-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     Sep 29 2018 12:24:41

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "main" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of main
entity main is
port (
    TVP_VIDEO : in std_logic_vector(9 downto 0);
    ADV_B : out std_logic_vector(7 downto 0);
    ADV_G : out std_logic_vector(7 downto 0);
    ADV_R : out std_logic_vector(7 downto 0);
    DEBUG : inout std_logic_vector(7 downto 0);
    TVP_CLK : in std_logic;
    ADV_CLK : out std_logic;
    TVP_HSYNC : in std_logic;
    ADV_HSYNC : out std_logic;
    TVP_VSYNC : in std_logic;
    ADV_VSYNC : out std_logic;
    ADV_BLANK_N : out std_logic;
    LED : out std_logic;
    ADV_SYNC_N : out std_logic);
end main;

-- Architecture of main
-- View name is \INTERFACE\
architecture \INTERFACE\ of main is

signal \N__24121\ : std_logic;
signal \N__24120\ : std_logic;
signal \N__24119\ : std_logic;
signal \N__24110\ : std_logic;
signal \N__24109\ : std_logic;
signal \N__24108\ : std_logic;
signal \N__24101\ : std_logic;
signal \N__24100\ : std_logic;
signal \N__24099\ : std_logic;
signal \N__24092\ : std_logic;
signal \N__24091\ : std_logic;
signal \N__24090\ : std_logic;
signal \N__24083\ : std_logic;
signal \N__24082\ : std_logic;
signal \N__24081\ : std_logic;
signal \N__24074\ : std_logic;
signal \N__24073\ : std_logic;
signal \N__24072\ : std_logic;
signal \N__24065\ : std_logic;
signal \N__24064\ : std_logic;
signal \N__24063\ : std_logic;
signal \N__24056\ : std_logic;
signal \N__24055\ : std_logic;
signal \N__24054\ : std_logic;
signal \N__24047\ : std_logic;
signal \N__24046\ : std_logic;
signal \N__24045\ : std_logic;
signal \N__24038\ : std_logic;
signal \N__24037\ : std_logic;
signal \N__24036\ : std_logic;
signal \N__24029\ : std_logic;
signal \N__24028\ : std_logic;
signal \N__24027\ : std_logic;
signal \N__24020\ : std_logic;
signal \N__24019\ : std_logic;
signal \N__24018\ : std_logic;
signal \N__24011\ : std_logic;
signal \N__24010\ : std_logic;
signal \N__24009\ : std_logic;
signal \N__24002\ : std_logic;
signal \N__24001\ : std_logic;
signal \N__24000\ : std_logic;
signal \N__23993\ : std_logic;
signal \N__23992\ : std_logic;
signal \N__23991\ : std_logic;
signal \N__23984\ : std_logic;
signal \N__23983\ : std_logic;
signal \N__23982\ : std_logic;
signal \N__23975\ : std_logic;
signal \N__23974\ : std_logic;
signal \N__23973\ : std_logic;
signal \N__23966\ : std_logic;
signal \N__23965\ : std_logic;
signal \N__23964\ : std_logic;
signal \N__23957\ : std_logic;
signal \N__23956\ : std_logic;
signal \N__23955\ : std_logic;
signal \N__23948\ : std_logic;
signal \N__23947\ : std_logic;
signal \N__23946\ : std_logic;
signal \N__23939\ : std_logic;
signal \N__23938\ : std_logic;
signal \N__23937\ : std_logic;
signal \N__23930\ : std_logic;
signal \N__23929\ : std_logic;
signal \N__23928\ : std_logic;
signal \N__23921\ : std_logic;
signal \N__23920\ : std_logic;
signal \N__23919\ : std_logic;
signal \N__23912\ : std_logic;
signal \N__23911\ : std_logic;
signal \N__23910\ : std_logic;
signal \N__23903\ : std_logic;
signal \N__23902\ : std_logic;
signal \N__23901\ : std_logic;
signal \N__23894\ : std_logic;
signal \N__23893\ : std_logic;
signal \N__23892\ : std_logic;
signal \N__23885\ : std_logic;
signal \N__23884\ : std_logic;
signal \N__23883\ : std_logic;
signal \N__23876\ : std_logic;
signal \N__23875\ : std_logic;
signal \N__23874\ : std_logic;
signal \N__23867\ : std_logic;
signal \N__23866\ : std_logic;
signal \N__23865\ : std_logic;
signal \N__23858\ : std_logic;
signal \N__23857\ : std_logic;
signal \N__23856\ : std_logic;
signal \N__23849\ : std_logic;
signal \N__23848\ : std_logic;
signal \N__23847\ : std_logic;
signal \N__23840\ : std_logic;
signal \N__23839\ : std_logic;
signal \N__23838\ : std_logic;
signal \N__23831\ : std_logic;
signal \N__23830\ : std_logic;
signal \N__23829\ : std_logic;
signal \N__23822\ : std_logic;
signal \N__23821\ : std_logic;
signal \N__23820\ : std_logic;
signal \N__23813\ : std_logic;
signal \N__23812\ : std_logic;
signal \N__23811\ : std_logic;
signal \N__23804\ : std_logic;
signal \N__23803\ : std_logic;
signal \N__23802\ : std_logic;
signal \N__23795\ : std_logic;
signal \N__23794\ : std_logic;
signal \N__23793\ : std_logic;
signal \N__23786\ : std_logic;
signal \N__23785\ : std_logic;
signal \N__23784\ : std_logic;
signal \N__23777\ : std_logic;
signal \N__23776\ : std_logic;
signal \N__23775\ : std_logic;
signal \N__23768\ : std_logic;
signal \N__23767\ : std_logic;
signal \N__23766\ : std_logic;
signal \N__23759\ : std_logic;
signal \N__23758\ : std_logic;
signal \N__23757\ : std_logic;
signal \N__23750\ : std_logic;
signal \N__23749\ : std_logic;
signal \N__23748\ : std_logic;
signal \N__23741\ : std_logic;
signal \N__23740\ : std_logic;
signal \N__23739\ : std_logic;
signal \N__23732\ : std_logic;
signal \N__23731\ : std_logic;
signal \N__23730\ : std_logic;
signal \N__23723\ : std_logic;
signal \N__23722\ : std_logic;
signal \N__23721\ : std_logic;
signal \N__23714\ : std_logic;
signal \N__23713\ : std_logic;
signal \N__23712\ : std_logic;
signal \N__23705\ : std_logic;
signal \N__23704\ : std_logic;
signal \N__23703\ : std_logic;
signal \N__23696\ : std_logic;
signal \N__23695\ : std_logic;
signal \N__23694\ : std_logic;
signal \N__23687\ : std_logic;
signal \N__23686\ : std_logic;
signal \N__23685\ : std_logic;
signal \N__23668\ : std_logic;
signal \N__23667\ : std_logic;
signal \N__23666\ : std_logic;
signal \N__23665\ : std_logic;
signal \N__23664\ : std_logic;
signal \N__23663\ : std_logic;
signal \N__23660\ : std_logic;
signal \N__23659\ : std_logic;
signal \N__23656\ : std_logic;
signal \N__23655\ : std_logic;
signal \N__23654\ : std_logic;
signal \N__23653\ : std_logic;
signal \N__23650\ : std_logic;
signal \N__23649\ : std_logic;
signal \N__23648\ : std_logic;
signal \N__23647\ : std_logic;
signal \N__23644\ : std_logic;
signal \N__23641\ : std_logic;
signal \N__23640\ : std_logic;
signal \N__23639\ : std_logic;
signal \N__23638\ : std_logic;
signal \N__23637\ : std_logic;
signal \N__23634\ : std_logic;
signal \N__23631\ : std_logic;
signal \N__23630\ : std_logic;
signal \N__23629\ : std_logic;
signal \N__23626\ : std_logic;
signal \N__23623\ : std_logic;
signal \N__23620\ : std_logic;
signal \N__23617\ : std_logic;
signal \N__23614\ : std_logic;
signal \N__23609\ : std_logic;
signal \N__23606\ : std_logic;
signal \N__23603\ : std_logic;
signal \N__23602\ : std_logic;
signal \N__23601\ : std_logic;
signal \N__23596\ : std_logic;
signal \N__23593\ : std_logic;
signal \N__23590\ : std_logic;
signal \N__23587\ : std_logic;
signal \N__23584\ : std_logic;
signal \N__23581\ : std_logic;
signal \N__23578\ : std_logic;
signal \N__23575\ : std_logic;
signal \N__23574\ : std_logic;
signal \N__23571\ : std_logic;
signal \N__23564\ : std_logic;
signal \N__23561\ : std_logic;
signal \N__23554\ : std_logic;
signal \N__23551\ : std_logic;
signal \N__23548\ : std_logic;
signal \N__23545\ : std_logic;
signal \N__23544\ : std_logic;
signal \N__23543\ : std_logic;
signal \N__23536\ : std_logic;
signal \N__23529\ : std_logic;
signal \N__23524\ : std_logic;
signal \N__23521\ : std_logic;
signal \N__23516\ : std_logic;
signal \N__23507\ : std_logic;
signal \N__23504\ : std_logic;
signal \N__23501\ : std_logic;
signal \N__23498\ : std_logic;
signal \N__23489\ : std_logic;
signal \N__23484\ : std_logic;
signal \N__23473\ : std_logic;
signal \N__23470\ : std_logic;
signal \N__23467\ : std_logic;
signal \N__23464\ : std_logic;
signal \N__23461\ : std_logic;
signal \N__23458\ : std_logic;
signal \N__23455\ : std_logic;
signal \N__23452\ : std_logic;
signal \N__23449\ : std_logic;
signal \N__23446\ : std_logic;
signal \N__23443\ : std_logic;
signal \N__23440\ : std_logic;
signal \N__23437\ : std_logic;
signal \N__23434\ : std_logic;
signal \N__23431\ : std_logic;
signal \N__23428\ : std_logic;
signal \N__23425\ : std_logic;
signal \N__23424\ : std_logic;
signal \N__23421\ : std_logic;
signal \N__23418\ : std_logic;
signal \N__23417\ : std_logic;
signal \N__23412\ : std_logic;
signal \N__23409\ : std_logic;
signal \N__23406\ : std_logic;
signal \N__23403\ : std_logic;
signal \N__23400\ : std_logic;
signal \N__23397\ : std_logic;
signal \N__23394\ : std_logic;
signal \N__23391\ : std_logic;
signal \N__23388\ : std_logic;
signal \N__23385\ : std_logic;
signal \N__23382\ : std_logic;
signal \N__23379\ : std_logic;
signal \N__23374\ : std_logic;
signal \N__23371\ : std_logic;
signal \N__23368\ : std_logic;
signal \N__23365\ : std_logic;
signal \N__23364\ : std_logic;
signal \N__23361\ : std_logic;
signal \N__23358\ : std_logic;
signal \N__23357\ : std_logic;
signal \N__23354\ : std_logic;
signal \N__23351\ : std_logic;
signal \N__23348\ : std_logic;
signal \N__23345\ : std_logic;
signal \N__23342\ : std_logic;
signal \N__23339\ : std_logic;
signal \N__23336\ : std_logic;
signal \N__23333\ : std_logic;
signal \N__23330\ : std_logic;
signal \N__23327\ : std_logic;
signal \N__23324\ : std_logic;
signal \N__23321\ : std_logic;
signal \N__23318\ : std_logic;
signal \N__23315\ : std_logic;
signal \N__23312\ : std_logic;
signal \N__23305\ : std_logic;
signal \N__23302\ : std_logic;
signal \N__23301\ : std_logic;
signal \N__23298\ : std_logic;
signal \N__23295\ : std_logic;
signal \N__23294\ : std_logic;
signal \N__23293\ : std_logic;
signal \N__23292\ : std_logic;
signal \N__23289\ : std_logic;
signal \N__23286\ : std_logic;
signal \N__23283\ : std_logic;
signal \N__23280\ : std_logic;
signal \N__23279\ : std_logic;
signal \N__23278\ : std_logic;
signal \N__23275\ : std_logic;
signal \N__23274\ : std_logic;
signal \N__23273\ : std_logic;
signal \N__23272\ : std_logic;
signal \N__23271\ : std_logic;
signal \N__23270\ : std_logic;
signal \N__23269\ : std_logic;
signal \N__23268\ : std_logic;
signal \N__23261\ : std_logic;
signal \N__23258\ : std_logic;
signal \N__23255\ : std_logic;
signal \N__23252\ : std_logic;
signal \N__23251\ : std_logic;
signal \N__23248\ : std_logic;
signal \N__23245\ : std_logic;
signal \N__23242\ : std_logic;
signal \N__23239\ : std_logic;
signal \N__23236\ : std_logic;
signal \N__23235\ : std_logic;
signal \N__23232\ : std_logic;
signal \N__23229\ : std_logic;
signal \N__23226\ : std_logic;
signal \N__23225\ : std_logic;
signal \N__23224\ : std_logic;
signal \N__23217\ : std_logic;
signal \N__23214\ : std_logic;
signal \N__23211\ : std_logic;
signal \N__23204\ : std_logic;
signal \N__23203\ : std_logic;
signal \N__23202\ : std_logic;
signal \N__23201\ : std_logic;
signal \N__23200\ : std_logic;
signal \N__23199\ : std_logic;
signal \N__23194\ : std_logic;
signal \N__23191\ : std_logic;
signal \N__23190\ : std_logic;
signal \N__23189\ : std_logic;
signal \N__23182\ : std_logic;
signal \N__23179\ : std_logic;
signal \N__23176\ : std_logic;
signal \N__23175\ : std_logic;
signal \N__23174\ : std_logic;
signal \N__23167\ : std_logic;
signal \N__23164\ : std_logic;
signal \N__23161\ : std_logic;
signal \N__23160\ : std_logic;
signal \N__23159\ : std_logic;
signal \N__23156\ : std_logic;
signal \N__23153\ : std_logic;
signal \N__23152\ : std_logic;
signal \N__23151\ : std_logic;
signal \N__23148\ : std_logic;
signal \N__23145\ : std_logic;
signal \N__23144\ : std_logic;
signal \N__23143\ : std_logic;
signal \N__23138\ : std_logic;
signal \N__23135\ : std_logic;
signal \N__23134\ : std_logic;
signal \N__23131\ : std_logic;
signal \N__23130\ : std_logic;
signal \N__23125\ : std_logic;
signal \N__23122\ : std_logic;
signal \N__23119\ : std_logic;
signal \N__23116\ : std_logic;
signal \N__23113\ : std_logic;
signal \N__23108\ : std_logic;
signal \N__23107\ : std_logic;
signal \N__23106\ : std_logic;
signal \N__23105\ : std_logic;
signal \N__23102\ : std_logic;
signal \N__23101\ : std_logic;
signal \N__23100\ : std_logic;
signal \N__23097\ : std_logic;
signal \N__23096\ : std_logic;
signal \N__23091\ : std_logic;
signal \N__23088\ : std_logic;
signal \N__23087\ : std_logic;
signal \N__23086\ : std_logic;
signal \N__23083\ : std_logic;
signal \N__23082\ : std_logic;
signal \N__23081\ : std_logic;
signal \N__23080\ : std_logic;
signal \N__23079\ : std_logic;
signal \N__23078\ : std_logic;
signal \N__23077\ : std_logic;
signal \N__23074\ : std_logic;
signal \N__23073\ : std_logic;
signal \N__23070\ : std_logic;
signal \N__23067\ : std_logic;
signal \N__23064\ : std_logic;
signal \N__23059\ : std_logic;
signal \N__23056\ : std_logic;
signal \N__23055\ : std_logic;
signal \N__23052\ : std_logic;
signal \N__23049\ : std_logic;
signal \N__23042\ : std_logic;
signal \N__23039\ : std_logic;
signal \N__23034\ : std_logic;
signal \N__23031\ : std_logic;
signal \N__23028\ : std_logic;
signal \N__23027\ : std_logic;
signal \N__23026\ : std_logic;
signal \N__23023\ : std_logic;
signal \N__23020\ : std_logic;
signal \N__23017\ : std_logic;
signal \N__23014\ : std_logic;
signal \N__23011\ : std_logic;
signal \N__23008\ : std_logic;
signal \N__23005\ : std_logic;
signal \N__23002\ : std_logic;
signal \N__22999\ : std_logic;
signal \N__22998\ : std_logic;
signal \N__22997\ : std_logic;
signal \N__22996\ : std_logic;
signal \N__22995\ : std_logic;
signal \N__22994\ : std_logic;
signal \N__22991\ : std_logic;
signal \N__22990\ : std_logic;
signal \N__22989\ : std_logic;
signal \N__22986\ : std_logic;
signal \N__22983\ : std_logic;
signal \N__22982\ : std_logic;
signal \N__22981\ : std_logic;
signal \N__22980\ : std_logic;
signal \N__22979\ : std_logic;
signal \N__22976\ : std_logic;
signal \N__22973\ : std_logic;
signal \N__22972\ : std_logic;
signal \N__22969\ : std_logic;
signal \N__22968\ : std_logic;
signal \N__22965\ : std_logic;
signal \N__22962\ : std_logic;
signal \N__22961\ : std_logic;
signal \N__22958\ : std_logic;
signal \N__22955\ : std_logic;
signal \N__22948\ : std_logic;
signal \N__22947\ : std_logic;
signal \N__22942\ : std_logic;
signal \N__22939\ : std_logic;
signal \N__22938\ : std_logic;
signal \N__22933\ : std_logic;
signal \N__22932\ : std_logic;
signal \N__22923\ : std_logic;
signal \N__22920\ : std_logic;
signal \N__22917\ : std_logic;
signal \N__22914\ : std_logic;
signal \N__22913\ : std_logic;
signal \N__22912\ : std_logic;
signal \N__22909\ : std_logic;
signal \N__22902\ : std_logic;
signal \N__22897\ : std_logic;
signal \N__22890\ : std_logic;
signal \N__22887\ : std_logic;
signal \N__22884\ : std_logic;
signal \N__22883\ : std_logic;
signal \N__22882\ : std_logic;
signal \N__22879\ : std_logic;
signal \N__22876\ : std_logic;
signal \N__22873\ : std_logic;
signal \N__22872\ : std_logic;
signal \N__22869\ : std_logic;
signal \N__22866\ : std_logic;
signal \N__22863\ : std_logic;
signal \N__22858\ : std_logic;
signal \N__22855\ : std_logic;
signal \N__22854\ : std_logic;
signal \N__22853\ : std_logic;
signal \N__22850\ : std_logic;
signal \N__22847\ : std_logic;
signal \N__22844\ : std_logic;
signal \N__22843\ : std_logic;
signal \N__22840\ : std_logic;
signal \N__22837\ : std_logic;
signal \N__22834\ : std_logic;
signal \N__22833\ : std_logic;
signal \N__22832\ : std_logic;
signal \N__22829\ : std_logic;
signal \N__22826\ : std_logic;
signal \N__22825\ : std_logic;
signal \N__22824\ : std_logic;
signal \N__22821\ : std_logic;
signal \N__22818\ : std_logic;
signal \N__22815\ : std_logic;
signal \N__22810\ : std_logic;
signal \N__22809\ : std_logic;
signal \N__22806\ : std_logic;
signal \N__22803\ : std_logic;
signal \N__22800\ : std_logic;
signal \N__22797\ : std_logic;
signal \N__22794\ : std_logic;
signal \N__22791\ : std_logic;
signal \N__22788\ : std_logic;
signal \N__22785\ : std_logic;
signal \N__22780\ : std_logic;
signal \N__22777\ : std_logic;
signal \N__22774\ : std_logic;
signal \N__22771\ : std_logic;
signal \N__22770\ : std_logic;
signal \N__22765\ : std_logic;
signal \N__22758\ : std_logic;
signal \N__22755\ : std_logic;
signal \N__22752\ : std_logic;
signal \N__22751\ : std_logic;
signal \N__22748\ : std_logic;
signal \N__22747\ : std_logic;
signal \N__22746\ : std_logic;
signal \N__22743\ : std_logic;
signal \N__22738\ : std_logic;
signal \N__22735\ : std_logic;
signal \N__22728\ : std_logic;
signal \N__22723\ : std_logic;
signal \N__22720\ : std_logic;
signal \N__22717\ : std_logic;
signal \N__22714\ : std_logic;
signal \N__22711\ : std_logic;
signal \N__22708\ : std_logic;
signal \N__22705\ : std_logic;
signal \N__22698\ : std_logic;
signal \N__22695\ : std_logic;
signal \N__22694\ : std_logic;
signal \N__22691\ : std_logic;
signal \N__22690\ : std_logic;
signal \N__22685\ : std_logic;
signal \N__22682\ : std_logic;
signal \N__22679\ : std_logic;
signal \N__22670\ : std_logic;
signal \N__22667\ : std_logic;
signal \N__22662\ : std_logic;
signal \N__22651\ : std_logic;
signal \N__22650\ : std_logic;
signal \N__22649\ : std_logic;
signal \N__22646\ : std_logic;
signal \N__22639\ : std_logic;
signal \N__22636\ : std_logic;
signal \N__22633\ : std_logic;
signal \N__22632\ : std_logic;
signal \N__22623\ : std_logic;
signal \N__22620\ : std_logic;
signal \N__22617\ : std_logic;
signal \N__22614\ : std_logic;
signal \N__22611\ : std_logic;
signal \N__22610\ : std_logic;
signal \N__22603\ : std_logic;
signal \N__22594\ : std_logic;
signal \N__22585\ : std_logic;
signal \N__22580\ : std_logic;
signal \N__22577\ : std_logic;
signal \N__22574\ : std_logic;
signal \N__22571\ : std_logic;
signal \N__22566\ : std_logic;
signal \N__22559\ : std_logic;
signal \N__22558\ : std_logic;
signal \N__22557\ : std_logic;
signal \N__22552\ : std_logic;
signal \N__22549\ : std_logic;
signal \N__22546\ : std_logic;
signal \N__22545\ : std_logic;
signal \N__22542\ : std_logic;
signal \N__22535\ : std_logic;
signal \N__22532\ : std_logic;
signal \N__22531\ : std_logic;
signal \N__22530\ : std_logic;
signal \N__22525\ : std_logic;
signal \N__22520\ : std_logic;
signal \N__22517\ : std_logic;
signal \N__22514\ : std_logic;
signal \N__22503\ : std_logic;
signal \N__22498\ : std_logic;
signal \N__22497\ : std_logic;
signal \N__22492\ : std_logic;
signal \N__22489\ : std_logic;
signal \N__22486\ : std_logic;
signal \N__22483\ : std_logic;
signal \N__22480\ : std_logic;
signal \N__22477\ : std_logic;
signal \N__22474\ : std_logic;
signal \N__22471\ : std_logic;
signal \N__22468\ : std_logic;
signal \N__22465\ : std_logic;
signal \N__22462\ : std_logic;
signal \N__22461\ : std_logic;
signal \N__22458\ : std_logic;
signal \N__22453\ : std_logic;
signal \N__22450\ : std_logic;
signal \N__22447\ : std_logic;
signal \N__22442\ : std_logic;
signal \N__22439\ : std_logic;
signal \N__22434\ : std_logic;
signal \N__22431\ : std_logic;
signal \N__22426\ : std_logic;
signal \N__22423\ : std_logic;
signal \N__22420\ : std_logic;
signal \N__22415\ : std_logic;
signal \N__22412\ : std_logic;
signal \N__22409\ : std_logic;
signal \N__22406\ : std_logic;
signal \N__22403\ : std_logic;
signal \N__22400\ : std_logic;
signal \N__22395\ : std_logic;
signal \N__22392\ : std_logic;
signal \N__22389\ : std_logic;
signal \N__22384\ : std_logic;
signal \N__22381\ : std_logic;
signal \N__22376\ : std_logic;
signal \N__22369\ : std_logic;
signal \N__22366\ : std_logic;
signal \N__22363\ : std_logic;
signal \N__22358\ : std_logic;
signal \N__22355\ : std_logic;
signal \N__22350\ : std_logic;
signal \N__22347\ : std_logic;
signal \N__22340\ : std_logic;
signal \N__22327\ : std_logic;
signal \N__22326\ : std_logic;
signal \N__22323\ : std_logic;
signal \N__22322\ : std_logic;
signal \N__22321\ : std_logic;
signal \N__22320\ : std_logic;
signal \N__22319\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22315\ : std_logic;
signal \N__22312\ : std_logic;
signal \N__22309\ : std_logic;
signal \N__22306\ : std_logic;
signal \N__22303\ : std_logic;
signal \N__22300\ : std_logic;
signal \N__22297\ : std_logic;
signal \N__22294\ : std_logic;
signal \N__22289\ : std_logic;
signal \N__22286\ : std_logic;
signal \N__22283\ : std_logic;
signal \N__22280\ : std_logic;
signal \N__22275\ : std_logic;
signal \N__22272\ : std_logic;
signal \N__22267\ : std_logic;
signal \N__22264\ : std_logic;
signal \N__22261\ : std_logic;
signal \N__22252\ : std_logic;
signal \N__22249\ : std_logic;
signal \N__22246\ : std_logic;
signal \N__22243\ : std_logic;
signal \N__22240\ : std_logic;
signal \N__22237\ : std_logic;
signal \N__22236\ : std_logic;
signal \N__22235\ : std_logic;
signal \N__22234\ : std_logic;
signal \N__22233\ : std_logic;
signal \N__22232\ : std_logic;
signal \N__22231\ : std_logic;
signal \N__22228\ : std_logic;
signal \N__22227\ : std_logic;
signal \N__22226\ : std_logic;
signal \N__22225\ : std_logic;
signal \N__22222\ : std_logic;
signal \N__22219\ : std_logic;
signal \N__22218\ : std_logic;
signal \N__22217\ : std_logic;
signal \N__22216\ : std_logic;
signal \N__22215\ : std_logic;
signal \N__22212\ : std_logic;
signal \N__22209\ : std_logic;
signal \N__22206\ : std_logic;
signal \N__22203\ : std_logic;
signal \N__22200\ : std_logic;
signal \N__22199\ : std_logic;
signal \N__22190\ : std_logic;
signal \N__22187\ : std_logic;
signal \N__22186\ : std_logic;
signal \N__22183\ : std_logic;
signal \N__22180\ : std_logic;
signal \N__22179\ : std_logic;
signal \N__22178\ : std_logic;
signal \N__22175\ : std_logic;
signal \N__22174\ : std_logic;
signal \N__22173\ : std_logic;
signal \N__22172\ : std_logic;
signal \N__22169\ : std_logic;
signal \N__22166\ : std_logic;
signal \N__22163\ : std_logic;
signal \N__22160\ : std_logic;
signal \N__22155\ : std_logic;
signal \N__22152\ : std_logic;
signal \N__22149\ : std_logic;
signal \N__22146\ : std_logic;
signal \N__22143\ : std_logic;
signal \N__22140\ : std_logic;
signal \N__22137\ : std_logic;
signal \N__22134\ : std_logic;
signal \N__22129\ : std_logic;
signal \N__22126\ : std_logic;
signal \N__22125\ : std_logic;
signal \N__22124\ : std_logic;
signal \N__22123\ : std_logic;
signal \N__22122\ : std_logic;
signal \N__22119\ : std_logic;
signal \N__22116\ : std_logic;
signal \N__22107\ : std_logic;
signal \N__22104\ : std_logic;
signal \N__22097\ : std_logic;
signal \N__22092\ : std_logic;
signal \N__22089\ : std_logic;
signal \N__22086\ : std_logic;
signal \N__22083\ : std_logic;
signal \N__22080\ : std_logic;
signal \N__22077\ : std_logic;
signal \N__22074\ : std_logic;
signal \N__22069\ : std_logic;
signal \N__22066\ : std_logic;
signal \N__22057\ : std_logic;
signal \N__22052\ : std_logic;
signal \N__22045\ : std_logic;
signal \N__22030\ : std_logic;
signal \N__22027\ : std_logic;
signal \N__22024\ : std_logic;
signal \N__22021\ : std_logic;
signal \N__22018\ : std_logic;
signal \N__22015\ : std_logic;
signal \N__22012\ : std_logic;
signal \N__22009\ : std_logic;
signal \N__22006\ : std_logic;
signal \N__22003\ : std_logic;
signal \N__22000\ : std_logic;
signal \N__21997\ : std_logic;
signal \N__21994\ : std_logic;
signal \N__21991\ : std_logic;
signal \N__21990\ : std_logic;
signal \N__21989\ : std_logic;
signal \N__21986\ : std_logic;
signal \N__21983\ : std_logic;
signal \N__21980\ : std_logic;
signal \N__21979\ : std_logic;
signal \N__21976\ : std_logic;
signal \N__21973\ : std_logic;
signal \N__21970\ : std_logic;
signal \N__21967\ : std_logic;
signal \N__21962\ : std_logic;
signal \N__21957\ : std_logic;
signal \N__21956\ : std_logic;
signal \N__21951\ : std_logic;
signal \N__21948\ : std_logic;
signal \N__21947\ : std_logic;
signal \N__21946\ : std_logic;
signal \N__21943\ : std_logic;
signal \N__21940\ : std_logic;
signal \N__21937\ : std_logic;
signal \N__21934\ : std_logic;
signal \N__21933\ : std_logic;
signal \N__21926\ : std_logic;
signal \N__21923\ : std_logic;
signal \N__21920\ : std_logic;
signal \N__21917\ : std_logic;
signal \N__21914\ : std_logic;
signal \N__21911\ : std_logic;
signal \N__21904\ : std_logic;
signal \N__21901\ : std_logic;
signal \N__21898\ : std_logic;
signal \N__21895\ : std_logic;
signal \N__21892\ : std_logic;
signal \N__21889\ : std_logic;
signal \N__21886\ : std_logic;
signal \N__21883\ : std_logic;
signal \N__21880\ : std_logic;
signal \N__21877\ : std_logic;
signal \N__21874\ : std_logic;
signal \N__21871\ : std_logic;
signal \N__21868\ : std_logic;
signal \N__21865\ : std_logic;
signal \N__21862\ : std_logic;
signal \N__21859\ : std_logic;
signal \N__21856\ : std_logic;
signal \N__21853\ : std_logic;
signal \N__21850\ : std_logic;
signal \N__21847\ : std_logic;
signal \N__21844\ : std_logic;
signal \N__21841\ : std_logic;
signal \N__21838\ : std_logic;
signal \N__21835\ : std_logic;
signal \N__21832\ : std_logic;
signal \N__21829\ : std_logic;
signal \N__21826\ : std_logic;
signal \N__21823\ : std_logic;
signal \N__21820\ : std_logic;
signal \N__21817\ : std_logic;
signal \N__21814\ : std_logic;
signal \N__21811\ : std_logic;
signal \N__21808\ : std_logic;
signal \N__21805\ : std_logic;
signal \N__21802\ : std_logic;
signal \N__21799\ : std_logic;
signal \N__21796\ : std_logic;
signal \N__21793\ : std_logic;
signal \N__21790\ : std_logic;
signal \N__21787\ : std_logic;
signal \N__21784\ : std_logic;
signal \N__21781\ : std_logic;
signal \N__21778\ : std_logic;
signal \N__21775\ : std_logic;
signal \N__21772\ : std_logic;
signal \N__21769\ : std_logic;
signal \N__21766\ : std_logic;
signal \N__21763\ : std_logic;
signal \N__21760\ : std_logic;
signal \N__21757\ : std_logic;
signal \N__21754\ : std_logic;
signal \N__21751\ : std_logic;
signal \N__21748\ : std_logic;
signal \N__21745\ : std_logic;
signal \N__21742\ : std_logic;
signal \N__21739\ : std_logic;
signal \N__21736\ : std_logic;
signal \N__21733\ : std_logic;
signal \N__21730\ : std_logic;
signal \N__21727\ : std_logic;
signal \N__21724\ : std_logic;
signal \N__21721\ : std_logic;
signal \N__21718\ : std_logic;
signal \N__21715\ : std_logic;
signal \N__21712\ : std_logic;
signal \N__21709\ : std_logic;
signal \N__21706\ : std_logic;
signal \N__21703\ : std_logic;
signal \N__21700\ : std_logic;
signal \N__21697\ : std_logic;
signal \N__21694\ : std_logic;
signal \N__21693\ : std_logic;
signal \N__21692\ : std_logic;
signal \N__21691\ : std_logic;
signal \N__21688\ : std_logic;
signal \N__21685\ : std_logic;
signal \N__21684\ : std_logic;
signal \N__21683\ : std_logic;
signal \N__21682\ : std_logic;
signal \N__21679\ : std_logic;
signal \N__21676\ : std_logic;
signal \N__21675\ : std_logic;
signal \N__21674\ : std_logic;
signal \N__21671\ : std_logic;
signal \N__21668\ : std_logic;
signal \N__21665\ : std_logic;
signal \N__21662\ : std_logic;
signal \N__21661\ : std_logic;
signal \N__21658\ : std_logic;
signal \N__21653\ : std_logic;
signal \N__21652\ : std_logic;
signal \N__21649\ : std_logic;
signal \N__21646\ : std_logic;
signal \N__21645\ : std_logic;
signal \N__21644\ : std_logic;
signal \N__21641\ : std_logic;
signal \N__21636\ : std_logic;
signal \N__21633\ : std_logic;
signal \N__21628\ : std_logic;
signal \N__21625\ : std_logic;
signal \N__21622\ : std_logic;
signal \N__21617\ : std_logic;
signal \N__21614\ : std_logic;
signal \N__21611\ : std_logic;
signal \N__21606\ : std_logic;
signal \N__21603\ : std_logic;
signal \N__21594\ : std_logic;
signal \N__21591\ : std_logic;
signal \N__21580\ : std_logic;
signal \N__21577\ : std_logic;
signal \N__21574\ : std_logic;
signal \N__21571\ : std_logic;
signal \N__21568\ : std_logic;
signal \N__21565\ : std_logic;
signal \N__21562\ : std_logic;
signal \N__21559\ : std_logic;
signal \N__21558\ : std_logic;
signal \N__21555\ : std_logic;
signal \N__21552\ : std_logic;
signal \N__21549\ : std_logic;
signal \N__21546\ : std_logic;
signal \N__21545\ : std_logic;
signal \N__21542\ : std_logic;
signal \N__21539\ : std_logic;
signal \N__21536\ : std_logic;
signal \N__21533\ : std_logic;
signal \N__21530\ : std_logic;
signal \N__21527\ : std_logic;
signal \N__21522\ : std_logic;
signal \N__21519\ : std_logic;
signal \N__21516\ : std_logic;
signal \N__21513\ : std_logic;
signal \N__21510\ : std_logic;
signal \N__21507\ : std_logic;
signal \N__21502\ : std_logic;
signal \N__21499\ : std_logic;
signal \N__21496\ : std_logic;
signal \N__21493\ : std_logic;
signal \N__21490\ : std_logic;
signal \N__21489\ : std_logic;
signal \N__21488\ : std_logic;
signal \N__21485\ : std_logic;
signal \N__21484\ : std_logic;
signal \N__21483\ : std_logic;
signal \N__21482\ : std_logic;
signal \N__21479\ : std_logic;
signal \N__21478\ : std_logic;
signal \N__21475\ : std_logic;
signal \N__21474\ : std_logic;
signal \N__21471\ : std_logic;
signal \N__21468\ : std_logic;
signal \N__21465\ : std_logic;
signal \N__21462\ : std_logic;
signal \N__21461\ : std_logic;
signal \N__21460\ : std_logic;
signal \N__21459\ : std_logic;
signal \N__21458\ : std_logic;
signal \N__21457\ : std_logic;
signal \N__21454\ : std_logic;
signal \N__21453\ : std_logic;
signal \N__21450\ : std_logic;
signal \N__21449\ : std_logic;
signal \N__21446\ : std_logic;
signal \N__21443\ : std_logic;
signal \N__21438\ : std_logic;
signal \N__21433\ : std_logic;
signal \N__21430\ : std_logic;
signal \N__21427\ : std_logic;
signal \N__21424\ : std_logic;
signal \N__21421\ : std_logic;
signal \N__21418\ : std_logic;
signal \N__21415\ : std_logic;
signal \N__21412\ : std_logic;
signal \N__21409\ : std_logic;
signal \N__21406\ : std_logic;
signal \N__21403\ : std_logic;
signal \N__21400\ : std_logic;
signal \N__21393\ : std_logic;
signal \N__21390\ : std_logic;
signal \N__21387\ : std_logic;
signal \N__21382\ : std_logic;
signal \N__21377\ : std_logic;
signal \N__21368\ : std_logic;
signal \N__21359\ : std_logic;
signal \N__21352\ : std_logic;
signal \N__21351\ : std_logic;
signal \N__21350\ : std_logic;
signal \N__21349\ : std_logic;
signal \N__21348\ : std_logic;
signal \N__21347\ : std_logic;
signal \N__21344\ : std_logic;
signal \N__21341\ : std_logic;
signal \N__21338\ : std_logic;
signal \N__21335\ : std_logic;
signal \N__21332\ : std_logic;
signal \N__21331\ : std_logic;
signal \N__21330\ : std_logic;
signal \N__21329\ : std_logic;
signal \N__21326\ : std_logic;
signal \N__21325\ : std_logic;
signal \N__21324\ : std_logic;
signal \N__21321\ : std_logic;
signal \N__21320\ : std_logic;
signal \N__21319\ : std_logic;
signal \N__21318\ : std_logic;
signal \N__21315\ : std_logic;
signal \N__21308\ : std_logic;
signal \N__21305\ : std_logic;
signal \N__21304\ : std_logic;
signal \N__21303\ : std_logic;
signal \N__21302\ : std_logic;
signal \N__21301\ : std_logic;
signal \N__21300\ : std_logic;
signal \N__21297\ : std_logic;
signal \N__21294\ : std_logic;
signal \N__21291\ : std_logic;
signal \N__21288\ : std_logic;
signal \N__21285\ : std_logic;
signal \N__21284\ : std_logic;
signal \N__21283\ : std_logic;
signal \N__21282\ : std_logic;
signal \N__21281\ : std_logic;
signal \N__21280\ : std_logic;
signal \N__21277\ : std_logic;
signal \N__21276\ : std_logic;
signal \N__21275\ : std_logic;
signal \N__21272\ : std_logic;
signal \N__21269\ : std_logic;
signal \N__21268\ : std_logic;
signal \N__21267\ : std_logic;
signal \N__21266\ : std_logic;
signal \N__21265\ : std_logic;
signal \N__21262\ : std_logic;
signal \N__21261\ : std_logic;
signal \N__21260\ : std_logic;
signal \N__21259\ : std_logic;
signal \N__21258\ : std_logic;
signal \N__21251\ : std_logic;
signal \N__21248\ : std_logic;
signal \N__21245\ : std_logic;
signal \N__21242\ : std_logic;
signal \N__21239\ : std_logic;
signal \N__21236\ : std_logic;
signal \N__21235\ : std_logic;
signal \N__21234\ : std_logic;
signal \N__21233\ : std_logic;
signal \N__21230\ : std_logic;
signal \N__21221\ : std_logic;
signal \N__21218\ : std_logic;
signal \N__21215\ : std_logic;
signal \N__21212\ : std_logic;
signal \N__21209\ : std_logic;
signal \N__21206\ : std_logic;
signal \N__21205\ : std_logic;
signal \N__21202\ : std_logic;
signal \N__21199\ : std_logic;
signal \N__21196\ : std_logic;
signal \N__21195\ : std_logic;
signal \N__21192\ : std_logic;
signal \N__21189\ : std_logic;
signal \N__21186\ : std_logic;
signal \N__21185\ : std_logic;
signal \N__21182\ : std_logic;
signal \N__21179\ : std_logic;
signal \N__21178\ : std_logic;
signal \N__21175\ : std_logic;
signal \N__21172\ : std_logic;
signal \N__21171\ : std_logic;
signal \N__21168\ : std_logic;
signal \N__21167\ : std_logic;
signal \N__21166\ : std_logic;
signal \N__21163\ : std_logic;
signal \N__21160\ : std_logic;
signal \N__21157\ : std_logic;
signal \N__21152\ : std_logic;
signal \N__21145\ : std_logic;
signal \N__21142\ : std_logic;
signal \N__21139\ : std_logic;
signal \N__21138\ : std_logic;
signal \N__21135\ : std_logic;
signal \N__21132\ : std_logic;
signal \N__21131\ : std_logic;
signal \N__21124\ : std_logic;
signal \N__21121\ : std_logic;
signal \N__21120\ : std_logic;
signal \N__21119\ : std_logic;
signal \N__21118\ : std_logic;
signal \N__21117\ : std_logic;
signal \N__21114\ : std_logic;
signal \N__21111\ : std_logic;
signal \N__21108\ : std_logic;
signal \N__21105\ : std_logic;
signal \N__21102\ : std_logic;
signal \N__21097\ : std_logic;
signal \N__21094\ : std_logic;
signal \N__21089\ : std_logic;
signal \N__21086\ : std_logic;
signal \N__21083\ : std_logic;
signal \N__21080\ : std_logic;
signal \N__21077\ : std_logic;
signal \N__21072\ : std_logic;
signal \N__21069\ : std_logic;
signal \N__21066\ : std_logic;
signal \N__21063\ : std_logic;
signal \N__21060\ : std_logic;
signal \N__21059\ : std_logic;
signal \N__21056\ : std_logic;
signal \N__21055\ : std_logic;
signal \N__21054\ : std_logic;
signal \N__21053\ : std_logic;
signal \N__21052\ : std_logic;
signal \N__21051\ : std_logic;
signal \N__21050\ : std_logic;
signal \N__21049\ : std_logic;
signal \N__21048\ : std_logic;
signal \N__21045\ : std_logic;
signal \N__21040\ : std_logic;
signal \N__21037\ : std_logic;
signal \N__21030\ : std_logic;
signal \N__21027\ : std_logic;
signal \N__21020\ : std_logic;
signal \N__21017\ : std_logic;
signal \N__21014\ : std_logic;
signal \N__21009\ : std_logic;
signal \N__21006\ : std_logic;
signal \N__21005\ : std_logic;
signal \N__21004\ : std_logic;
signal \N__21003\ : std_logic;
signal \N__21002\ : std_logic;
signal \N__20999\ : std_logic;
signal \N__20992\ : std_logic;
signal \N__20989\ : std_logic;
signal \N__20982\ : std_logic;
signal \N__20977\ : std_logic;
signal \N__20974\ : std_logic;
signal \N__20969\ : std_logic;
signal \N__20966\ : std_logic;
signal \N__20963\ : std_logic;
signal \N__20960\ : std_logic;
signal \N__20957\ : std_logic;
signal \N__20952\ : std_logic;
signal \N__20945\ : std_logic;
signal \N__20942\ : std_logic;
signal \N__20937\ : std_logic;
signal \N__20934\ : std_logic;
signal \N__20931\ : std_logic;
signal \N__20928\ : std_logic;
signal \N__20925\ : std_logic;
signal \N__20918\ : std_logic;
signal \N__20915\ : std_logic;
signal \N__20908\ : std_logic;
signal \N__20903\ : std_logic;
signal \N__20898\ : std_logic;
signal \N__20893\ : std_logic;
signal \N__20886\ : std_logic;
signal \N__20873\ : std_logic;
signal \N__20864\ : std_logic;
signal \N__20833\ : std_logic;
signal \N__20830\ : std_logic;
signal \N__20827\ : std_logic;
signal \N__20824\ : std_logic;
signal \N__20821\ : std_logic;
signal \N__20818\ : std_logic;
signal \N__20815\ : std_logic;
signal \N__20812\ : std_logic;
signal \N__20809\ : std_logic;
signal \N__20806\ : std_logic;
signal \N__20803\ : std_logic;
signal \N__20800\ : std_logic;
signal \N__20797\ : std_logic;
signal \N__20794\ : std_logic;
signal \N__20791\ : std_logic;
signal \N__20788\ : std_logic;
signal \N__20785\ : std_logic;
signal \N__20782\ : std_logic;
signal \N__20779\ : std_logic;
signal \N__20776\ : std_logic;
signal \N__20773\ : std_logic;
signal \N__20770\ : std_logic;
signal \N__20767\ : std_logic;
signal \N__20764\ : std_logic;
signal \N__20761\ : std_logic;
signal \N__20758\ : std_logic;
signal \N__20755\ : std_logic;
signal \N__20752\ : std_logic;
signal \N__20749\ : std_logic;
signal \N__20746\ : std_logic;
signal \N__20743\ : std_logic;
signal \N__20740\ : std_logic;
signal \N__20737\ : std_logic;
signal \N__20734\ : std_logic;
signal \N__20731\ : std_logic;
signal \N__20728\ : std_logic;
signal \N__20725\ : std_logic;
signal \N__20722\ : std_logic;
signal \N__20719\ : std_logic;
signal \N__20716\ : std_logic;
signal \N__20713\ : std_logic;
signal \N__20710\ : std_logic;
signal \N__20707\ : std_logic;
signal \N__20704\ : std_logic;
signal \N__20701\ : std_logic;
signal \N__20698\ : std_logic;
signal \N__20697\ : std_logic;
signal \N__20696\ : std_logic;
signal \N__20695\ : std_logic;
signal \N__20694\ : std_logic;
signal \N__20693\ : std_logic;
signal \N__20680\ : std_logic;
signal \N__20679\ : std_logic;
signal \N__20678\ : std_logic;
signal \N__20675\ : std_logic;
signal \N__20674\ : std_logic;
signal \N__20673\ : std_logic;
signal \N__20672\ : std_logic;
signal \N__20669\ : std_logic;
signal \N__20666\ : std_logic;
signal \N__20663\ : std_logic;
signal \N__20658\ : std_logic;
signal \N__20655\ : std_logic;
signal \N__20652\ : std_logic;
signal \N__20647\ : std_logic;
signal \N__20644\ : std_logic;
signal \N__20637\ : std_logic;
signal \N__20636\ : std_logic;
signal \N__20635\ : std_logic;
signal \N__20634\ : std_logic;
signal \N__20633\ : std_logic;
signal \N__20632\ : std_logic;
signal \N__20631\ : std_logic;
signal \N__20630\ : std_logic;
signal \N__20629\ : std_logic;
signal \N__20628\ : std_logic;
signal \N__20625\ : std_logic;
signal \N__20622\ : std_logic;
signal \N__20617\ : std_logic;
signal \N__20614\ : std_logic;
signal \N__20611\ : std_logic;
signal \N__20608\ : std_logic;
signal \N__20599\ : std_logic;
signal \N__20584\ : std_logic;
signal \N__20581\ : std_logic;
signal \N__20578\ : std_logic;
signal \N__20575\ : std_logic;
signal \N__20572\ : std_logic;
signal \N__20569\ : std_logic;
signal \N__20568\ : std_logic;
signal \N__20567\ : std_logic;
signal \N__20566\ : std_logic;
signal \N__20565\ : std_logic;
signal \N__20564\ : std_logic;
signal \N__20561\ : std_logic;
signal \N__20558\ : std_logic;
signal \N__20557\ : std_logic;
signal \N__20554\ : std_logic;
signal \N__20551\ : std_logic;
signal \N__20546\ : std_logic;
signal \N__20537\ : std_logic;
signal \N__20536\ : std_logic;
signal \N__20535\ : std_logic;
signal \N__20534\ : std_logic;
signal \N__20531\ : std_logic;
signal \N__20528\ : std_logic;
signal \N__20525\ : std_logic;
signal \N__20522\ : std_logic;
signal \N__20521\ : std_logic;
signal \N__20518\ : std_logic;
signal \N__20515\ : std_logic;
signal \N__20512\ : std_logic;
signal \N__20507\ : std_logic;
signal \N__20504\ : std_logic;
signal \N__20503\ : std_logic;
signal \N__20498\ : std_logic;
signal \N__20495\ : std_logic;
signal \N__20492\ : std_logic;
signal \N__20487\ : std_logic;
signal \N__20484\ : std_logic;
signal \N__20483\ : std_logic;
signal \N__20480\ : std_logic;
signal \N__20477\ : std_logic;
signal \N__20472\ : std_logic;
signal \N__20469\ : std_logic;
signal \N__20466\ : std_logic;
signal \N__20465\ : std_logic;
signal \N__20464\ : std_logic;
signal \N__20463\ : std_logic;
signal \N__20462\ : std_logic;
signal \N__20459\ : std_logic;
signal \N__20456\ : std_logic;
signal \N__20449\ : std_logic;
signal \N__20446\ : std_logic;
signal \N__20439\ : std_logic;
signal \N__20436\ : std_logic;
signal \N__20427\ : std_logic;
signal \N__20422\ : std_logic;
signal \N__20421\ : std_logic;
signal \N__20418\ : std_logic;
signal \N__20415\ : std_logic;
signal \N__20412\ : std_logic;
signal \N__20409\ : std_logic;
signal \N__20406\ : std_logic;
signal \N__20403\ : std_logic;
signal \N__20400\ : std_logic;
signal \N__20397\ : std_logic;
signal \N__20394\ : std_logic;
signal \N__20391\ : std_logic;
signal \N__20388\ : std_logic;
signal \N__20385\ : std_logic;
signal \N__20382\ : std_logic;
signal \N__20379\ : std_logic;
signal \N__20376\ : std_logic;
signal \N__20373\ : std_logic;
signal \N__20370\ : std_logic;
signal \N__20367\ : std_logic;
signal \N__20364\ : std_logic;
signal \N__20361\ : std_logic;
signal \N__20358\ : std_logic;
signal \N__20355\ : std_logic;
signal \N__20352\ : std_logic;
signal \N__20349\ : std_logic;
signal \N__20346\ : std_logic;
signal \N__20343\ : std_logic;
signal \N__20340\ : std_logic;
signal \N__20337\ : std_logic;
signal \N__20334\ : std_logic;
signal \N__20331\ : std_logic;
signal \N__20328\ : std_logic;
signal \N__20325\ : std_logic;
signal \N__20322\ : std_logic;
signal \N__20319\ : std_logic;
signal \N__20316\ : std_logic;
signal \N__20313\ : std_logic;
signal \N__20310\ : std_logic;
signal \N__20307\ : std_logic;
signal \N__20304\ : std_logic;
signal \N__20301\ : std_logic;
signal \N__20298\ : std_logic;
signal \N__20295\ : std_logic;
signal \N__20292\ : std_logic;
signal \N__20289\ : std_logic;
signal \N__20286\ : std_logic;
signal \N__20283\ : std_logic;
signal \N__20280\ : std_logic;
signal \N__20277\ : std_logic;
signal \N__20274\ : std_logic;
signal \N__20271\ : std_logic;
signal \N__20268\ : std_logic;
signal \N__20265\ : std_logic;
signal \N__20262\ : std_logic;
signal \N__20259\ : std_logic;
signal \N__20256\ : std_logic;
signal \N__20253\ : std_logic;
signal \N__20250\ : std_logic;
signal \N__20247\ : std_logic;
signal \N__20244\ : std_logic;
signal \N__20241\ : std_logic;
signal \N__20240\ : std_logic;
signal \N__20237\ : std_logic;
signal \N__20234\ : std_logic;
signal \N__20231\ : std_logic;
signal \N__20228\ : std_logic;
signal \N__20225\ : std_logic;
signal \N__20222\ : std_logic;
signal \N__20219\ : std_logic;
signal \N__20216\ : std_logic;
signal \N__20213\ : std_logic;
signal \N__20210\ : std_logic;
signal \N__20209\ : std_logic;
signal \N__20206\ : std_logic;
signal \N__20203\ : std_logic;
signal \N__20200\ : std_logic;
signal \N__20197\ : std_logic;
signal \N__20194\ : std_logic;
signal \N__20189\ : std_logic;
signal \N__20182\ : std_logic;
signal \N__20179\ : std_logic;
signal \N__20178\ : std_logic;
signal \N__20177\ : std_logic;
signal \N__20176\ : std_logic;
signal \N__20175\ : std_logic;
signal \N__20174\ : std_logic;
signal \N__20173\ : std_logic;
signal \N__20172\ : std_logic;
signal \N__20171\ : std_logic;
signal \N__20170\ : std_logic;
signal \N__20167\ : std_logic;
signal \N__20166\ : std_logic;
signal \N__20165\ : std_logic;
signal \N__20164\ : std_logic;
signal \N__20163\ : std_logic;
signal \N__20162\ : std_logic;
signal \N__20161\ : std_logic;
signal \N__20160\ : std_logic;
signal \N__20159\ : std_logic;
signal \N__20158\ : std_logic;
signal \N__20157\ : std_logic;
signal \N__20156\ : std_logic;
signal \N__20155\ : std_logic;
signal \N__20154\ : std_logic;
signal \N__20153\ : std_logic;
signal \N__20152\ : std_logic;
signal \N__20151\ : std_logic;
signal \N__20150\ : std_logic;
signal \N__20149\ : std_logic;
signal \N__20148\ : std_logic;
signal \N__20147\ : std_logic;
signal \N__20146\ : std_logic;
signal \N__20145\ : std_logic;
signal \N__20144\ : std_logic;
signal \N__20143\ : std_logic;
signal \N__20142\ : std_logic;
signal \N__20141\ : std_logic;
signal \N__20140\ : std_logic;
signal \N__20139\ : std_logic;
signal \N__20138\ : std_logic;
signal \N__20137\ : std_logic;
signal \N__20136\ : std_logic;
signal \N__20135\ : std_logic;
signal \N__20134\ : std_logic;
signal \N__20133\ : std_logic;
signal \N__20132\ : std_logic;
signal \N__20131\ : std_logic;
signal \N__20130\ : std_logic;
signal \N__20129\ : std_logic;
signal \N__20128\ : std_logic;
signal \N__20029\ : std_logic;
signal \N__20026\ : std_logic;
signal \N__20023\ : std_logic;
signal \N__20020\ : std_logic;
signal \N__20017\ : std_logic;
signal \N__20014\ : std_logic;
signal \N__20011\ : std_logic;
signal \N__20008\ : std_logic;
signal \N__20005\ : std_logic;
signal \N__20002\ : std_logic;
signal \N__19999\ : std_logic;
signal \N__19996\ : std_logic;
signal \N__19993\ : std_logic;
signal \N__19990\ : std_logic;
signal \N__19987\ : std_logic;
signal \N__19984\ : std_logic;
signal \N__19981\ : std_logic;
signal \N__19978\ : std_logic;
signal \N__19975\ : std_logic;
signal \N__19972\ : std_logic;
signal \N__19969\ : std_logic;
signal \N__19966\ : std_logic;
signal \N__19963\ : std_logic;
signal \N__19960\ : std_logic;
signal \N__19957\ : std_logic;
signal \N__19954\ : std_logic;
signal \N__19951\ : std_logic;
signal \N__19948\ : std_logic;
signal \N__19945\ : std_logic;
signal \N__19942\ : std_logic;
signal \N__19939\ : std_logic;
signal \N__19936\ : std_logic;
signal \N__19933\ : std_logic;
signal \N__19930\ : std_logic;
signal \N__19927\ : std_logic;
signal \N__19924\ : std_logic;
signal \N__19921\ : std_logic;
signal \N__19918\ : std_logic;
signal \N__19915\ : std_logic;
signal \N__19912\ : std_logic;
signal \N__19909\ : std_logic;
signal \N__19906\ : std_logic;
signal \N__19905\ : std_logic;
signal \N__19902\ : std_logic;
signal \N__19899\ : std_logic;
signal \N__19898\ : std_logic;
signal \N__19895\ : std_logic;
signal \N__19892\ : std_logic;
signal \N__19889\ : std_logic;
signal \N__19886\ : std_logic;
signal \N__19883\ : std_logic;
signal \N__19880\ : std_logic;
signal \N__19877\ : std_logic;
signal \N__19874\ : std_logic;
signal \N__19871\ : std_logic;
signal \N__19866\ : std_logic;
signal \N__19863\ : std_logic;
signal \N__19860\ : std_logic;
signal \N__19855\ : std_logic;
signal \N__19852\ : std_logic;
signal \N__19851\ : std_logic;
signal \N__19850\ : std_logic;
signal \N__19847\ : std_logic;
signal \N__19844\ : std_logic;
signal \N__19843\ : std_logic;
signal \N__19840\ : std_logic;
signal \N__19839\ : std_logic;
signal \N__19838\ : std_logic;
signal \N__19833\ : std_logic;
signal \N__19830\ : std_logic;
signal \N__19829\ : std_logic;
signal \N__19826\ : std_logic;
signal \N__19823\ : std_logic;
signal \N__19820\ : std_logic;
signal \N__19819\ : std_logic;
signal \N__19818\ : std_logic;
signal \N__19813\ : std_logic;
signal \N__19810\ : std_logic;
signal \N__19809\ : std_logic;
signal \N__19808\ : std_logic;
signal \N__19807\ : std_logic;
signal \N__19802\ : std_logic;
signal \N__19799\ : std_logic;
signal \N__19796\ : std_logic;
signal \N__19793\ : std_logic;
signal \N__19792\ : std_logic;
signal \N__19791\ : std_logic;
signal \N__19786\ : std_logic;
signal \N__19783\ : std_logic;
signal \N__19780\ : std_logic;
signal \N__19777\ : std_logic;
signal \N__19776\ : std_logic;
signal \N__19769\ : std_logic;
signal \N__19766\ : std_logic;
signal \N__19763\ : std_logic;
signal \N__19760\ : std_logic;
signal \N__19759\ : std_logic;
signal \N__19758\ : std_logic;
signal \N__19757\ : std_logic;
signal \N__19752\ : std_logic;
signal \N__19747\ : std_logic;
signal \N__19744\ : std_logic;
signal \N__19743\ : std_logic;
signal \N__19742\ : std_logic;
signal \N__19739\ : std_logic;
signal \N__19734\ : std_logic;
signal \N__19731\ : std_logic;
signal \N__19728\ : std_logic;
signal \N__19725\ : std_logic;
signal \N__19724\ : std_logic;
signal \N__19723\ : std_logic;
signal \N__19720\ : std_logic;
signal \N__19719\ : std_logic;
signal \N__19718\ : std_logic;
signal \N__19715\ : std_logic;
signal \N__19712\ : std_logic;
signal \N__19709\ : std_logic;
signal \N__19706\ : std_logic;
signal \N__19705\ : std_logic;
signal \N__19704\ : std_logic;
signal \N__19701\ : std_logic;
signal \N__19700\ : std_logic;
signal \N__19699\ : std_logic;
signal \N__19690\ : std_logic;
signal \N__19687\ : std_logic;
signal \N__19684\ : std_logic;
signal \N__19681\ : std_logic;
signal \N__19680\ : std_logic;
signal \N__19677\ : std_logic;
signal \N__19674\ : std_logic;
signal \N__19671\ : std_logic;
signal \N__19668\ : std_logic;
signal \N__19661\ : std_logic;
signal \N__19658\ : std_logic;
signal \N__19657\ : std_logic;
signal \N__19656\ : std_logic;
signal \N__19653\ : std_logic;
signal \N__19652\ : std_logic;
signal \N__19649\ : std_logic;
signal \N__19646\ : std_logic;
signal \N__19643\ : std_logic;
signal \N__19636\ : std_logic;
signal \N__19633\ : std_logic;
signal \N__19630\ : std_logic;
signal \N__19629\ : std_logic;
signal \N__19622\ : std_logic;
signal \N__19615\ : std_logic;
signal \N__19612\ : std_logic;
signal \N__19609\ : std_logic;
signal \N__19606\ : std_logic;
signal \N__19603\ : std_logic;
signal \N__19602\ : std_logic;
signal \N__19595\ : std_logic;
signal \N__19588\ : std_logic;
signal \N__19585\ : std_logic;
signal \N__19580\ : std_logic;
signal \N__19575\ : std_logic;
signal \N__19572\ : std_logic;
signal \N__19569\ : std_logic;
signal \N__19566\ : std_logic;
signal \N__19563\ : std_logic;
signal \N__19558\ : std_logic;
signal \N__19555\ : std_logic;
signal \N__19552\ : std_logic;
signal \N__19547\ : std_logic;
signal \N__19544\ : std_logic;
signal \N__19539\ : std_logic;
signal \N__19534\ : std_logic;
signal \N__19529\ : std_logic;
signal \N__19526\ : std_logic;
signal \N__19519\ : std_logic;
signal \N__19516\ : std_logic;
signal \N__19513\ : std_logic;
signal \N__19510\ : std_logic;
signal \N__19507\ : std_logic;
signal \N__19504\ : std_logic;
signal \N__19501\ : std_logic;
signal \N__19498\ : std_logic;
signal \N__19495\ : std_logic;
signal \N__19492\ : std_logic;
signal \N__19489\ : std_logic;
signal \N__19486\ : std_logic;
signal \N__19483\ : std_logic;
signal \N__19480\ : std_logic;
signal \N__19477\ : std_logic;
signal \N__19474\ : std_logic;
signal \N__19471\ : std_logic;
signal \N__19468\ : std_logic;
signal \N__19465\ : std_logic;
signal \N__19462\ : std_logic;
signal \N__19459\ : std_logic;
signal \N__19456\ : std_logic;
signal \N__19453\ : std_logic;
signal \N__19450\ : std_logic;
signal \N__19447\ : std_logic;
signal \N__19444\ : std_logic;
signal \N__19441\ : std_logic;
signal \N__19438\ : std_logic;
signal \N__19435\ : std_logic;
signal \N__19432\ : std_logic;
signal \N__19429\ : std_logic;
signal \N__19426\ : std_logic;
signal \N__19423\ : std_logic;
signal \N__19420\ : std_logic;
signal \N__19417\ : std_logic;
signal \N__19414\ : std_logic;
signal \N__19411\ : std_logic;
signal \N__19408\ : std_logic;
signal \N__19405\ : std_logic;
signal \N__19402\ : std_logic;
signal \N__19399\ : std_logic;
signal \N__19396\ : std_logic;
signal \N__19393\ : std_logic;
signal \N__19390\ : std_logic;
signal \N__19387\ : std_logic;
signal \N__19384\ : std_logic;
signal \N__19381\ : std_logic;
signal \N__19378\ : std_logic;
signal \N__19375\ : std_logic;
signal \N__19372\ : std_logic;
signal \N__19369\ : std_logic;
signal \N__19366\ : std_logic;
signal \N__19363\ : std_logic;
signal \N__19360\ : std_logic;
signal \N__19357\ : std_logic;
signal \N__19354\ : std_logic;
signal \N__19351\ : std_logic;
signal \N__19348\ : std_logic;
signal \N__19345\ : std_logic;
signal \N__19342\ : std_logic;
signal \N__19339\ : std_logic;
signal \N__19338\ : std_logic;
signal \N__19337\ : std_logic;
signal \N__19334\ : std_logic;
signal \N__19329\ : std_logic;
signal \N__19324\ : std_logic;
signal \N__19321\ : std_logic;
signal \N__19320\ : std_logic;
signal \N__19319\ : std_logic;
signal \N__19316\ : std_logic;
signal \N__19311\ : std_logic;
signal \N__19306\ : std_logic;
signal \N__19303\ : std_logic;
signal \N__19302\ : std_logic;
signal \N__19301\ : std_logic;
signal \N__19298\ : std_logic;
signal \N__19293\ : std_logic;
signal \N__19288\ : std_logic;
signal \N__19285\ : std_logic;
signal \N__19284\ : std_logic;
signal \N__19283\ : std_logic;
signal \N__19280\ : std_logic;
signal \N__19275\ : std_logic;
signal \N__19270\ : std_logic;
signal \N__19267\ : std_logic;
signal \N__19266\ : std_logic;
signal \N__19263\ : std_logic;
signal \N__19260\ : std_logic;
signal \N__19255\ : std_logic;
signal \N__19252\ : std_logic;
signal \N__19249\ : std_logic;
signal \N__19248\ : std_logic;
signal \N__19245\ : std_logic;
signal \N__19242\ : std_logic;
signal \N__19239\ : std_logic;
signal \N__19234\ : std_logic;
signal \N__19233\ : std_logic;
signal \N__19230\ : std_logic;
signal \N__19227\ : std_logic;
signal \N__19224\ : std_logic;
signal \N__19221\ : std_logic;
signal \N__19218\ : std_logic;
signal \N__19213\ : std_logic;
signal \N__19210\ : std_logic;
signal \N__19207\ : std_logic;
signal \N__19204\ : std_logic;
signal \N__19201\ : std_logic;
signal \N__19198\ : std_logic;
signal \N__19195\ : std_logic;
signal \N__19192\ : std_logic;
signal \N__19189\ : std_logic;
signal \N__19186\ : std_logic;
signal \N__19183\ : std_logic;
signal \N__19180\ : std_logic;
signal \N__19177\ : std_logic;
signal \N__19174\ : std_logic;
signal \N__19171\ : std_logic;
signal \N__19168\ : std_logic;
signal \N__19165\ : std_logic;
signal \N__19162\ : std_logic;
signal \N__19159\ : std_logic;
signal \N__19156\ : std_logic;
signal \N__19153\ : std_logic;
signal \N__19150\ : std_logic;
signal \N__19147\ : std_logic;
signal \N__19144\ : std_logic;
signal \N__19141\ : std_logic;
signal \N__19138\ : std_logic;
signal \N__19135\ : std_logic;
signal \N__19132\ : std_logic;
signal \N__19129\ : std_logic;
signal \N__19126\ : std_logic;
signal \N__19123\ : std_logic;
signal \N__19120\ : std_logic;
signal \N__19117\ : std_logic;
signal \N__19114\ : std_logic;
signal \N__19113\ : std_logic;
signal \N__19110\ : std_logic;
signal \N__19109\ : std_logic;
signal \N__19106\ : std_logic;
signal \N__19103\ : std_logic;
signal \N__19100\ : std_logic;
signal \N__19099\ : std_logic;
signal \N__19098\ : std_logic;
signal \N__19097\ : std_logic;
signal \N__19094\ : std_logic;
signal \N__19093\ : std_logic;
signal \N__19090\ : std_logic;
signal \N__19087\ : std_logic;
signal \N__19086\ : std_logic;
signal \N__19083\ : std_logic;
signal \N__19082\ : std_logic;
signal \N__19081\ : std_logic;
signal \N__19080\ : std_logic;
signal \N__19079\ : std_logic;
signal \N__19078\ : std_logic;
signal \N__19077\ : std_logic;
signal \N__19072\ : std_logic;
signal \N__19069\ : std_logic;
signal \N__19068\ : std_logic;
signal \N__19067\ : std_logic;
signal \N__19066\ : std_logic;
signal \N__19065\ : std_logic;
signal \N__19064\ : std_logic;
signal \N__19061\ : std_logic;
signal \N__19060\ : std_logic;
signal \N__19059\ : std_logic;
signal \N__19054\ : std_logic;
signal \N__19051\ : std_logic;
signal \N__19048\ : std_logic;
signal \N__19043\ : std_logic;
signal \N__19034\ : std_logic;
signal \N__19031\ : std_logic;
signal \N__19028\ : std_logic;
signal \N__19025\ : std_logic;
signal \N__19024\ : std_logic;
signal \N__19023\ : std_logic;
signal \N__19022\ : std_logic;
signal \N__19019\ : std_logic;
signal \N__19014\ : std_logic;
signal \N__19011\ : std_logic;
signal \N__19008\ : std_logic;
signal \N__19003\ : std_logic;
signal \N__18998\ : std_logic;
signal \N__18993\ : std_logic;
signal \N__18990\ : std_logic;
signal \N__18989\ : std_logic;
signal \N__18988\ : std_logic;
signal \N__18987\ : std_logic;
signal \N__18982\ : std_logic;
signal \N__18979\ : std_logic;
signal \N__18976\ : std_logic;
signal \N__18971\ : std_logic;
signal \N__18966\ : std_logic;
signal \N__18957\ : std_logic;
signal \N__18954\ : std_logic;
signal \N__18951\ : std_logic;
signal \N__18948\ : std_logic;
signal \N__18943\ : std_logic;
signal \N__18940\ : std_logic;
signal \N__18929\ : std_logic;
signal \N__18916\ : std_logic;
signal \N__18913\ : std_logic;
signal \N__18912\ : std_logic;
signal \N__18909\ : std_logic;
signal \N__18906\ : std_logic;
signal \N__18903\ : std_logic;
signal \N__18898\ : std_logic;
signal \N__18895\ : std_logic;
signal \N__18892\ : std_logic;
signal \N__18889\ : std_logic;
signal \N__18886\ : std_logic;
signal \N__18885\ : std_logic;
signal \N__18882\ : std_logic;
signal \N__18879\ : std_logic;
signal \N__18876\ : std_logic;
signal \N__18873\ : std_logic;
signal \N__18870\ : std_logic;
signal \N__18867\ : std_logic;
signal \N__18864\ : std_logic;
signal \N__18861\ : std_logic;
signal \N__18858\ : std_logic;
signal \N__18855\ : std_logic;
signal \N__18852\ : std_logic;
signal \N__18849\ : std_logic;
signal \N__18846\ : std_logic;
signal \N__18843\ : std_logic;
signal \N__18840\ : std_logic;
signal \N__18837\ : std_logic;
signal \N__18834\ : std_logic;
signal \N__18831\ : std_logic;
signal \N__18828\ : std_logic;
signal \N__18825\ : std_logic;
signal \N__18822\ : std_logic;
signal \N__18819\ : std_logic;
signal \N__18816\ : std_logic;
signal \N__18813\ : std_logic;
signal \N__18810\ : std_logic;
signal \N__18807\ : std_logic;
signal \N__18804\ : std_logic;
signal \N__18801\ : std_logic;
signal \N__18798\ : std_logic;
signal \N__18795\ : std_logic;
signal \N__18792\ : std_logic;
signal \N__18789\ : std_logic;
signal \N__18786\ : std_logic;
signal \N__18783\ : std_logic;
signal \N__18780\ : std_logic;
signal \N__18777\ : std_logic;
signal \N__18774\ : std_logic;
signal \N__18771\ : std_logic;
signal \N__18768\ : std_logic;
signal \N__18765\ : std_logic;
signal \N__18762\ : std_logic;
signal \N__18759\ : std_logic;
signal \N__18756\ : std_logic;
signal \N__18753\ : std_logic;
signal \N__18750\ : std_logic;
signal \N__18747\ : std_logic;
signal \N__18744\ : std_logic;
signal \N__18741\ : std_logic;
signal \N__18738\ : std_logic;
signal \N__18735\ : std_logic;
signal \N__18732\ : std_logic;
signal \N__18729\ : std_logic;
signal \N__18726\ : std_logic;
signal \N__18723\ : std_logic;
signal \N__18720\ : std_logic;
signal \N__18717\ : std_logic;
signal \N__18714\ : std_logic;
signal \N__18711\ : std_logic;
signal \N__18708\ : std_logic;
signal \N__18705\ : std_logic;
signal \N__18702\ : std_logic;
signal \N__18699\ : std_logic;
signal \N__18696\ : std_logic;
signal \N__18693\ : std_logic;
signal \N__18690\ : std_logic;
signal \N__18687\ : std_logic;
signal \N__18684\ : std_logic;
signal \N__18681\ : std_logic;
signal \N__18678\ : std_logic;
signal \N__18675\ : std_logic;
signal \N__18672\ : std_logic;
signal \N__18669\ : std_logic;
signal \N__18664\ : std_logic;
signal \N__18661\ : std_logic;
signal \N__18658\ : std_logic;
signal \N__18655\ : std_logic;
signal \N__18652\ : std_logic;
signal \N__18651\ : std_logic;
signal \N__18646\ : std_logic;
signal \N__18645\ : std_logic;
signal \N__18642\ : std_logic;
signal \N__18639\ : std_logic;
signal \N__18636\ : std_logic;
signal \N__18633\ : std_logic;
signal \N__18628\ : std_logic;
signal \N__18625\ : std_logic;
signal \N__18622\ : std_logic;
signal \N__18619\ : std_logic;
signal \N__18616\ : std_logic;
signal \N__18613\ : std_logic;
signal \N__18610\ : std_logic;
signal \N__18607\ : std_logic;
signal \N__18604\ : std_logic;
signal \N__18601\ : std_logic;
signal \N__18598\ : std_logic;
signal \N__18595\ : std_logic;
signal \N__18594\ : std_logic;
signal \N__18593\ : std_logic;
signal \N__18590\ : std_logic;
signal \N__18585\ : std_logic;
signal \N__18580\ : std_logic;
signal \N__18577\ : std_logic;
signal \N__18574\ : std_logic;
signal \N__18571\ : std_logic;
signal \N__18568\ : std_logic;
signal \N__18567\ : std_logic;
signal \N__18564\ : std_logic;
signal \N__18561\ : std_logic;
signal \N__18556\ : std_logic;
signal \N__18553\ : std_logic;
signal \N__18550\ : std_logic;
signal \N__18549\ : std_logic;
signal \N__18546\ : std_logic;
signal \N__18543\ : std_logic;
signal \N__18538\ : std_logic;
signal \N__18535\ : std_logic;
signal \N__18534\ : std_logic;
signal \N__18531\ : std_logic;
signal \N__18528\ : std_logic;
signal \N__18525\ : std_logic;
signal \N__18522\ : std_logic;
signal \N__18519\ : std_logic;
signal \N__18516\ : std_logic;
signal \N__18513\ : std_logic;
signal \N__18510\ : std_logic;
signal \N__18507\ : std_logic;
signal \N__18504\ : std_logic;
signal \N__18501\ : std_logic;
signal \N__18498\ : std_logic;
signal \N__18495\ : std_logic;
signal \N__18492\ : std_logic;
signal \N__18489\ : std_logic;
signal \N__18486\ : std_logic;
signal \N__18483\ : std_logic;
signal \N__18480\ : std_logic;
signal \N__18477\ : std_logic;
signal \N__18474\ : std_logic;
signal \N__18471\ : std_logic;
signal \N__18468\ : std_logic;
signal \N__18465\ : std_logic;
signal \N__18462\ : std_logic;
signal \N__18459\ : std_logic;
signal \N__18456\ : std_logic;
signal \N__18453\ : std_logic;
signal \N__18450\ : std_logic;
signal \N__18447\ : std_logic;
signal \N__18444\ : std_logic;
signal \N__18441\ : std_logic;
signal \N__18438\ : std_logic;
signal \N__18435\ : std_logic;
signal \N__18432\ : std_logic;
signal \N__18429\ : std_logic;
signal \N__18426\ : std_logic;
signal \N__18423\ : std_logic;
signal \N__18420\ : std_logic;
signal \N__18417\ : std_logic;
signal \N__18414\ : std_logic;
signal \N__18411\ : std_logic;
signal \N__18408\ : std_logic;
signal \N__18405\ : std_logic;
signal \N__18402\ : std_logic;
signal \N__18399\ : std_logic;
signal \N__18396\ : std_logic;
signal \N__18393\ : std_logic;
signal \N__18390\ : std_logic;
signal \N__18387\ : std_logic;
signal \N__18384\ : std_logic;
signal \N__18381\ : std_logic;
signal \N__18378\ : std_logic;
signal \N__18375\ : std_logic;
signal \N__18372\ : std_logic;
signal \N__18369\ : std_logic;
signal \N__18366\ : std_logic;
signal \N__18363\ : std_logic;
signal \N__18360\ : std_logic;
signal \N__18357\ : std_logic;
signal \N__18354\ : std_logic;
signal \N__18351\ : std_logic;
signal \N__18348\ : std_logic;
signal \N__18345\ : std_logic;
signal \N__18342\ : std_logic;
signal \N__18339\ : std_logic;
signal \N__18336\ : std_logic;
signal \N__18333\ : std_logic;
signal \N__18330\ : std_logic;
signal \N__18327\ : std_logic;
signal \N__18324\ : std_logic;
signal \N__18319\ : std_logic;
signal \N__18316\ : std_logic;
signal \N__18315\ : std_logic;
signal \N__18314\ : std_logic;
signal \N__18311\ : std_logic;
signal \N__18308\ : std_logic;
signal \N__18307\ : std_logic;
signal \N__18304\ : std_logic;
signal \N__18303\ : std_logic;
signal \N__18302\ : std_logic;
signal \N__18301\ : std_logic;
signal \N__18300\ : std_logic;
signal \N__18299\ : std_logic;
signal \N__18298\ : std_logic;
signal \N__18295\ : std_logic;
signal \N__18294\ : std_logic;
signal \N__18291\ : std_logic;
signal \N__18288\ : std_logic;
signal \N__18285\ : std_logic;
signal \N__18280\ : std_logic;
signal \N__18275\ : std_logic;
signal \N__18274\ : std_logic;
signal \N__18273\ : std_logic;
signal \N__18270\ : std_logic;
signal \N__18269\ : std_logic;
signal \N__18266\ : std_logic;
signal \N__18263\ : std_logic;
signal \N__18260\ : std_logic;
signal \N__18257\ : std_logic;
signal \N__18250\ : std_logic;
signal \N__18247\ : std_logic;
signal \N__18242\ : std_logic;
signal \N__18237\ : std_logic;
signal \N__18220\ : std_logic;
signal \N__18217\ : std_logic;
signal \N__18214\ : std_logic;
signal \N__18211\ : std_logic;
signal \N__18208\ : std_logic;
signal \N__18205\ : std_logic;
signal \N__18202\ : std_logic;
signal \N__18199\ : std_logic;
signal \N__18196\ : std_logic;
signal \N__18193\ : std_logic;
signal \N__18192\ : std_logic;
signal \N__18189\ : std_logic;
signal \N__18186\ : std_logic;
signal \N__18183\ : std_logic;
signal \N__18180\ : std_logic;
signal \N__18177\ : std_logic;
signal \N__18174\ : std_logic;
signal \N__18171\ : std_logic;
signal \N__18168\ : std_logic;
signal \N__18165\ : std_logic;
signal \N__18162\ : std_logic;
signal \N__18159\ : std_logic;
signal \N__18156\ : std_logic;
signal \N__18153\ : std_logic;
signal \N__18150\ : std_logic;
signal \N__18147\ : std_logic;
signal \N__18144\ : std_logic;
signal \N__18141\ : std_logic;
signal \N__18138\ : std_logic;
signal \N__18135\ : std_logic;
signal \N__18132\ : std_logic;
signal \N__18129\ : std_logic;
signal \N__18126\ : std_logic;
signal \N__18123\ : std_logic;
signal \N__18120\ : std_logic;
signal \N__18117\ : std_logic;
signal \N__18114\ : std_logic;
signal \N__18111\ : std_logic;
signal \N__18108\ : std_logic;
signal \N__18105\ : std_logic;
signal \N__18102\ : std_logic;
signal \N__18099\ : std_logic;
signal \N__18096\ : std_logic;
signal \N__18093\ : std_logic;
signal \N__18090\ : std_logic;
signal \N__18087\ : std_logic;
signal \N__18084\ : std_logic;
signal \N__18081\ : std_logic;
signal \N__18078\ : std_logic;
signal \N__18075\ : std_logic;
signal \N__18072\ : std_logic;
signal \N__18069\ : std_logic;
signal \N__18066\ : std_logic;
signal \N__18063\ : std_logic;
signal \N__18060\ : std_logic;
signal \N__18057\ : std_logic;
signal \N__18054\ : std_logic;
signal \N__18051\ : std_logic;
signal \N__18048\ : std_logic;
signal \N__18045\ : std_logic;
signal \N__18042\ : std_logic;
signal \N__18039\ : std_logic;
signal \N__18036\ : std_logic;
signal \N__18033\ : std_logic;
signal \N__18030\ : std_logic;
signal \N__18027\ : std_logic;
signal \N__18024\ : std_logic;
signal \N__18021\ : std_logic;
signal \N__18018\ : std_logic;
signal \N__18015\ : std_logic;
signal \N__18012\ : std_logic;
signal \N__18009\ : std_logic;
signal \N__18006\ : std_logic;
signal \N__18003\ : std_logic;
signal \N__18000\ : std_logic;
signal \N__17997\ : std_logic;
signal \N__17994\ : std_logic;
signal \N__17991\ : std_logic;
signal \N__17988\ : std_logic;
signal \N__17983\ : std_logic;
signal \N__17980\ : std_logic;
signal \N__17979\ : std_logic;
signal \N__17976\ : std_logic;
signal \N__17973\ : std_logic;
signal \N__17972\ : std_logic;
signal \N__17969\ : std_logic;
signal \N__17966\ : std_logic;
signal \N__17963\ : std_logic;
signal \N__17956\ : std_logic;
signal \N__17955\ : std_logic;
signal \N__17952\ : std_logic;
signal \N__17949\ : std_logic;
signal \N__17944\ : std_logic;
signal \N__17941\ : std_logic;
signal \N__17938\ : std_logic;
signal \N__17937\ : std_logic;
signal \N__17934\ : std_logic;
signal \N__17933\ : std_logic;
signal \N__17930\ : std_logic;
signal \N__17929\ : std_logic;
signal \N__17928\ : std_logic;
signal \N__17927\ : std_logic;
signal \N__17924\ : std_logic;
signal \N__17921\ : std_logic;
signal \N__17918\ : std_logic;
signal \N__17915\ : std_logic;
signal \N__17912\ : std_logic;
signal \N__17909\ : std_logic;
signal \N__17908\ : std_logic;
signal \N__17907\ : std_logic;
signal \N__17906\ : std_logic;
signal \N__17905\ : std_logic;
signal \N__17900\ : std_logic;
signal \N__17897\ : std_logic;
signal \N__17894\ : std_logic;
signal \N__17891\ : std_logic;
signal \N__17888\ : std_logic;
signal \N__17885\ : std_logic;
signal \N__17884\ : std_logic;
signal \N__17883\ : std_logic;
signal \N__17882\ : std_logic;
signal \N__17881\ : std_logic;
signal \N__17878\ : std_logic;
signal \N__17875\ : std_logic;
signal \N__17872\ : std_logic;
signal \N__17863\ : std_logic;
signal \N__17858\ : std_logic;
signal \N__17855\ : std_logic;
signal \N__17852\ : std_logic;
signal \N__17849\ : std_logic;
signal \N__17846\ : std_logic;
signal \N__17827\ : std_logic;
signal \N__17824\ : std_logic;
signal \N__17821\ : std_logic;
signal \N__17820\ : std_logic;
signal \N__17817\ : std_logic;
signal \N__17814\ : std_logic;
signal \N__17809\ : std_logic;
signal \N__17808\ : std_logic;
signal \N__17807\ : std_logic;
signal \N__17800\ : std_logic;
signal \N__17797\ : std_logic;
signal \N__17796\ : std_logic;
signal \N__17793\ : std_logic;
signal \N__17790\ : std_logic;
signal \N__17785\ : std_logic;
signal \N__17782\ : std_logic;
signal \N__17779\ : std_logic;
signal \N__17778\ : std_logic;
signal \N__17775\ : std_logic;
signal \N__17774\ : std_logic;
signal \N__17771\ : std_logic;
signal \N__17770\ : std_logic;
signal \N__17767\ : std_logic;
signal \N__17766\ : std_logic;
signal \N__17763\ : std_logic;
signal \N__17762\ : std_logic;
signal \N__17759\ : std_logic;
signal \N__17756\ : std_logic;
signal \N__17753\ : std_logic;
signal \N__17750\ : std_logic;
signal \N__17747\ : std_logic;
signal \N__17744\ : std_logic;
signal \N__17743\ : std_logic;
signal \N__17738\ : std_logic;
signal \N__17733\ : std_logic;
signal \N__17728\ : std_logic;
signal \N__17725\ : std_logic;
signal \N__17720\ : std_logic;
signal \N__17717\ : std_logic;
signal \N__17714\ : std_logic;
signal \N__17707\ : std_logic;
signal \N__17704\ : std_logic;
signal \N__17701\ : std_logic;
signal \N__17698\ : std_logic;
signal \N__17697\ : std_logic;
signal \N__17694\ : std_logic;
signal \N__17693\ : std_logic;
signal \N__17690\ : std_logic;
signal \N__17687\ : std_logic;
signal \N__17684\ : std_logic;
signal \N__17681\ : std_logic;
signal \N__17678\ : std_logic;
signal \N__17675\ : std_logic;
signal \N__17672\ : std_logic;
signal \N__17669\ : std_logic;
signal \N__17666\ : std_logic;
signal \N__17663\ : std_logic;
signal \N__17660\ : std_logic;
signal \N__17657\ : std_logic;
signal \N__17654\ : std_logic;
signal \N__17651\ : std_logic;
signal \N__17646\ : std_logic;
signal \N__17643\ : std_logic;
signal \N__17638\ : std_logic;
signal \N__17635\ : std_logic;
signal \N__17632\ : std_logic;
signal \N__17629\ : std_logic;
signal \N__17628\ : std_logic;
signal \N__17625\ : std_logic;
signal \N__17624\ : std_logic;
signal \N__17621\ : std_logic;
signal \N__17618\ : std_logic;
signal \N__17615\ : std_logic;
signal \N__17612\ : std_logic;
signal \N__17609\ : std_logic;
signal \N__17606\ : std_logic;
signal \N__17601\ : std_logic;
signal \N__17598\ : std_logic;
signal \N__17595\ : std_logic;
signal \N__17592\ : std_logic;
signal \N__17589\ : std_logic;
signal \N__17586\ : std_logic;
signal \N__17581\ : std_logic;
signal \N__17578\ : std_logic;
signal \N__17575\ : std_logic;
signal \N__17572\ : std_logic;
signal \N__17569\ : std_logic;
signal \N__17566\ : std_logic;
signal \N__17563\ : std_logic;
signal \N__17560\ : std_logic;
signal \N__17557\ : std_logic;
signal \N__17554\ : std_logic;
signal \N__17551\ : std_logic;
signal \N__17548\ : std_logic;
signal \N__17545\ : std_logic;
signal \N__17542\ : std_logic;
signal \N__17539\ : std_logic;
signal \N__17536\ : std_logic;
signal \N__17533\ : std_logic;
signal \N__17530\ : std_logic;
signal \N__17527\ : std_logic;
signal \N__17524\ : std_logic;
signal \N__17521\ : std_logic;
signal \N__17518\ : std_logic;
signal \N__17515\ : std_logic;
signal \N__17512\ : std_logic;
signal \N__17509\ : std_logic;
signal \N__17506\ : std_logic;
signal \N__17503\ : std_logic;
signal \N__17500\ : std_logic;
signal \N__17497\ : std_logic;
signal \N__17494\ : std_logic;
signal \N__17491\ : std_logic;
signal \N__17488\ : std_logic;
signal \N__17485\ : std_logic;
signal \N__17482\ : std_logic;
signal \N__17479\ : std_logic;
signal \N__17476\ : std_logic;
signal \N__17473\ : std_logic;
signal \N__17470\ : std_logic;
signal \N__17467\ : std_logic;
signal \N__17464\ : std_logic;
signal \N__17461\ : std_logic;
signal \N__17458\ : std_logic;
signal \N__17455\ : std_logic;
signal \N__17452\ : std_logic;
signal \N__17449\ : std_logic;
signal \N__17446\ : std_logic;
signal \N__17443\ : std_logic;
signal \N__17440\ : std_logic;
signal \N__17437\ : std_logic;
signal \N__17434\ : std_logic;
signal \N__17431\ : std_logic;
signal \N__17428\ : std_logic;
signal \N__17425\ : std_logic;
signal \N__17422\ : std_logic;
signal \N__17419\ : std_logic;
signal \N__17416\ : std_logic;
signal \N__17413\ : std_logic;
signal \N__17410\ : std_logic;
signal \N__17407\ : std_logic;
signal \N__17404\ : std_logic;
signal \N__17401\ : std_logic;
signal \N__17398\ : std_logic;
signal \N__17395\ : std_logic;
signal \N__17392\ : std_logic;
signal \N__17389\ : std_logic;
signal \N__17386\ : std_logic;
signal \N__17383\ : std_logic;
signal \N__17380\ : std_logic;
signal \N__17377\ : std_logic;
signal \N__17374\ : std_logic;
signal \N__17371\ : std_logic;
signal \N__17368\ : std_logic;
signal \N__17365\ : std_logic;
signal \N__17362\ : std_logic;
signal \N__17359\ : std_logic;
signal \N__17356\ : std_logic;
signal \N__17353\ : std_logic;
signal \N__17352\ : std_logic;
signal \N__17351\ : std_logic;
signal \N__17350\ : std_logic;
signal \N__17347\ : std_logic;
signal \N__17342\ : std_logic;
signal \N__17337\ : std_logic;
signal \N__17332\ : std_logic;
signal \N__17331\ : std_logic;
signal \N__17330\ : std_logic;
signal \N__17329\ : std_logic;
signal \N__17326\ : std_logic;
signal \N__17323\ : std_logic;
signal \N__17320\ : std_logic;
signal \N__17315\ : std_logic;
signal \N__17308\ : std_logic;
signal \N__17305\ : std_logic;
signal \N__17302\ : std_logic;
signal \N__17299\ : std_logic;
signal \N__17296\ : std_logic;
signal \N__17293\ : std_logic;
signal \N__17292\ : std_logic;
signal \N__17287\ : std_logic;
signal \N__17284\ : std_logic;
signal \N__17283\ : std_logic;
signal \N__17280\ : std_logic;
signal \N__17277\ : std_logic;
signal \N__17274\ : std_logic;
signal \N__17271\ : std_logic;
signal \N__17268\ : std_logic;
signal \N__17265\ : std_logic;
signal \N__17262\ : std_logic;
signal \N__17259\ : std_logic;
signal \N__17256\ : std_logic;
signal \N__17253\ : std_logic;
signal \N__17250\ : std_logic;
signal \N__17247\ : std_logic;
signal \N__17244\ : std_logic;
signal \N__17241\ : std_logic;
signal \N__17238\ : std_logic;
signal \N__17235\ : std_logic;
signal \N__17232\ : std_logic;
signal \N__17229\ : std_logic;
signal \N__17226\ : std_logic;
signal \N__17223\ : std_logic;
signal \N__17220\ : std_logic;
signal \N__17217\ : std_logic;
signal \N__17214\ : std_logic;
signal \N__17211\ : std_logic;
signal \N__17208\ : std_logic;
signal \N__17205\ : std_logic;
signal \N__17202\ : std_logic;
signal \N__17199\ : std_logic;
signal \N__17196\ : std_logic;
signal \N__17193\ : std_logic;
signal \N__17190\ : std_logic;
signal \N__17187\ : std_logic;
signal \N__17184\ : std_logic;
signal \N__17181\ : std_logic;
signal \N__17178\ : std_logic;
signal \N__17175\ : std_logic;
signal \N__17172\ : std_logic;
signal \N__17169\ : std_logic;
signal \N__17166\ : std_logic;
signal \N__17163\ : std_logic;
signal \N__17160\ : std_logic;
signal \N__17157\ : std_logic;
signal \N__17154\ : std_logic;
signal \N__17151\ : std_logic;
signal \N__17148\ : std_logic;
signal \N__17145\ : std_logic;
signal \N__17142\ : std_logic;
signal \N__17139\ : std_logic;
signal \N__17136\ : std_logic;
signal \N__17133\ : std_logic;
signal \N__17130\ : std_logic;
signal \N__17127\ : std_logic;
signal \N__17124\ : std_logic;
signal \N__17121\ : std_logic;
signal \N__17118\ : std_logic;
signal \N__17115\ : std_logic;
signal \N__17112\ : std_logic;
signal \N__17109\ : std_logic;
signal \N__17106\ : std_logic;
signal \N__17103\ : std_logic;
signal \N__17100\ : std_logic;
signal \N__17097\ : std_logic;
signal \N__17094\ : std_logic;
signal \N__17091\ : std_logic;
signal \N__17088\ : std_logic;
signal \N__17085\ : std_logic;
signal \N__17082\ : std_logic;
signal \N__17079\ : std_logic;
signal \N__17076\ : std_logic;
signal \N__17073\ : std_logic;
signal \N__17070\ : std_logic;
signal \N__17067\ : std_logic;
signal \N__17064\ : std_logic;
signal \N__17061\ : std_logic;
signal \N__17058\ : std_logic;
signal \N__17053\ : std_logic;
signal \N__17050\ : std_logic;
signal \N__17047\ : std_logic;
signal \N__17044\ : std_logic;
signal \N__17041\ : std_logic;
signal \N__17040\ : std_logic;
signal \N__17037\ : std_logic;
signal \N__17034\ : std_logic;
signal \N__17033\ : std_logic;
signal \N__17028\ : std_logic;
signal \N__17025\ : std_logic;
signal \N__17024\ : std_logic;
signal \N__17019\ : std_logic;
signal \N__17016\ : std_logic;
signal \N__17013\ : std_logic;
signal \N__17010\ : std_logic;
signal \N__17007\ : std_logic;
signal \N__17004\ : std_logic;
signal \N__17001\ : std_logic;
signal \N__16998\ : std_logic;
signal \N__16995\ : std_logic;
signal \N__16992\ : std_logic;
signal \N__16987\ : std_logic;
signal \N__16986\ : std_logic;
signal \N__16983\ : std_logic;
signal \N__16980\ : std_logic;
signal \N__16977\ : std_logic;
signal \N__16976\ : std_logic;
signal \N__16973\ : std_logic;
signal \N__16972\ : std_logic;
signal \N__16969\ : std_logic;
signal \N__16966\ : std_logic;
signal \N__16963\ : std_logic;
signal \N__16960\ : std_logic;
signal \N__16957\ : std_logic;
signal \N__16954\ : std_logic;
signal \N__16949\ : std_logic;
signal \N__16942\ : std_logic;
signal \N__16939\ : std_logic;
signal \N__16936\ : std_logic;
signal \N__16935\ : std_logic;
signal \N__16932\ : std_logic;
signal \N__16929\ : std_logic;
signal \N__16928\ : std_logic;
signal \N__16925\ : std_logic;
signal \N__16922\ : std_logic;
signal \N__16919\ : std_logic;
signal \N__16912\ : std_logic;
signal \N__16909\ : std_logic;
signal \N__16908\ : std_logic;
signal \N__16905\ : std_logic;
signal \N__16902\ : std_logic;
signal \N__16897\ : std_logic;
signal \N__16894\ : std_logic;
signal \N__16891\ : std_logic;
signal \N__16888\ : std_logic;
signal \N__16885\ : std_logic;
signal \N__16882\ : std_logic;
signal \N__16879\ : std_logic;
signal \N__16876\ : std_logic;
signal \N__16873\ : std_logic;
signal \N__16870\ : std_logic;
signal \N__16867\ : std_logic;
signal \N__16864\ : std_logic;
signal \N__16863\ : std_logic;
signal \N__16862\ : std_logic;
signal \N__16859\ : std_logic;
signal \N__16858\ : std_logic;
signal \N__16855\ : std_logic;
signal \N__16852\ : std_logic;
signal \N__16849\ : std_logic;
signal \N__16846\ : std_logic;
signal \N__16843\ : std_logic;
signal \N__16834\ : std_logic;
signal \N__16831\ : std_logic;
signal \N__16828\ : std_logic;
signal \N__16825\ : std_logic;
signal \N__16824\ : std_logic;
signal \N__16821\ : std_logic;
signal \N__16818\ : std_logic;
signal \N__16817\ : std_logic;
signal \N__16812\ : std_logic;
signal \N__16809\ : std_logic;
signal \N__16808\ : std_logic;
signal \N__16803\ : std_logic;
signal \N__16800\ : std_logic;
signal \N__16795\ : std_logic;
signal \N__16792\ : std_logic;
signal \N__16789\ : std_logic;
signal \N__16786\ : std_logic;
signal \N__16785\ : std_logic;
signal \N__16784\ : std_logic;
signal \N__16783\ : std_logic;
signal \N__16782\ : std_logic;
signal \N__16781\ : std_logic;
signal \N__16780\ : std_logic;
signal \N__16779\ : std_logic;
signal \N__16776\ : std_logic;
signal \N__16773\ : std_logic;
signal \N__16772\ : std_logic;
signal \N__16769\ : std_logic;
signal \N__16762\ : std_logic;
signal \N__16757\ : std_logic;
signal \N__16750\ : std_logic;
signal \N__16741\ : std_logic;
signal \N__16740\ : std_logic;
signal \N__16739\ : std_logic;
signal \N__16738\ : std_logic;
signal \N__16737\ : std_logic;
signal \N__16736\ : std_logic;
signal \N__16735\ : std_logic;
signal \N__16732\ : std_logic;
signal \N__16729\ : std_logic;
signal \N__16726\ : std_logic;
signal \N__16725\ : std_logic;
signal \N__16724\ : std_logic;
signal \N__16721\ : std_logic;
signal \N__16718\ : std_logic;
signal \N__16711\ : std_logic;
signal \N__16708\ : std_logic;
signal \N__16705\ : std_logic;
signal \N__16698\ : std_logic;
signal \N__16687\ : std_logic;
signal \N__16686\ : std_logic;
signal \N__16685\ : std_logic;
signal \N__16682\ : std_logic;
signal \N__16679\ : std_logic;
signal \N__16678\ : std_logic;
signal \N__16677\ : std_logic;
signal \N__16676\ : std_logic;
signal \N__16675\ : std_logic;
signal \N__16674\ : std_logic;
signal \N__16673\ : std_logic;
signal \N__16670\ : std_logic;
signal \N__16665\ : std_logic;
signal \N__16662\ : std_logic;
signal \N__16657\ : std_logic;
signal \N__16650\ : std_logic;
signal \N__16639\ : std_logic;
signal \N__16638\ : std_logic;
signal \N__16635\ : std_logic;
signal \N__16634\ : std_logic;
signal \N__16631\ : std_logic;
signal \N__16628\ : std_logic;
signal \N__16625\ : std_logic;
signal \N__16624\ : std_logic;
signal \N__16621\ : std_logic;
signal \N__16618\ : std_logic;
signal \N__16615\ : std_logic;
signal \N__16612\ : std_logic;
signal \N__16609\ : std_logic;
signal \N__16604\ : std_logic;
signal \N__16601\ : std_logic;
signal \N__16598\ : std_logic;
signal \N__16595\ : std_logic;
signal \N__16592\ : std_logic;
signal \N__16587\ : std_logic;
signal \N__16584\ : std_logic;
signal \N__16581\ : std_logic;
signal \N__16578\ : std_logic;
signal \N__16573\ : std_logic;
signal \N__16570\ : std_logic;
signal \N__16567\ : std_logic;
signal \N__16564\ : std_logic;
signal \N__16561\ : std_logic;
signal \N__16558\ : std_logic;
signal \N__16555\ : std_logic;
signal \N__16552\ : std_logic;
signal \N__16549\ : std_logic;
signal \N__16546\ : std_logic;
signal \N__16543\ : std_logic;
signal \N__16540\ : std_logic;
signal \N__16537\ : std_logic;
signal \N__16534\ : std_logic;
signal \N__16531\ : std_logic;
signal \N__16528\ : std_logic;
signal \N__16525\ : std_logic;
signal \N__16522\ : std_logic;
signal \N__16519\ : std_logic;
signal \N__16516\ : std_logic;
signal \N__16513\ : std_logic;
signal \N__16510\ : std_logic;
signal \N__16507\ : std_logic;
signal \N__16504\ : std_logic;
signal \N__16501\ : std_logic;
signal \N__16498\ : std_logic;
signal \N__16495\ : std_logic;
signal \N__16492\ : std_logic;
signal \N__16491\ : std_logic;
signal \N__16490\ : std_logic;
signal \N__16487\ : std_logic;
signal \N__16484\ : std_logic;
signal \N__16483\ : std_logic;
signal \N__16480\ : std_logic;
signal \N__16475\ : std_logic;
signal \N__16472\ : std_logic;
signal \N__16469\ : std_logic;
signal \N__16464\ : std_logic;
signal \N__16461\ : std_logic;
signal \N__16458\ : std_logic;
signal \N__16455\ : std_logic;
signal \N__16452\ : std_logic;
signal \N__16447\ : std_logic;
signal \N__16446\ : std_logic;
signal \N__16443\ : std_logic;
signal \N__16440\ : std_logic;
signal \N__16439\ : std_logic;
signal \N__16438\ : std_logic;
signal \N__16433\ : std_logic;
signal \N__16430\ : std_logic;
signal \N__16427\ : std_logic;
signal \N__16420\ : std_logic;
signal \N__16417\ : std_logic;
signal \N__16414\ : std_logic;
signal \N__16411\ : std_logic;
signal \N__16408\ : std_logic;
signal \N__16405\ : std_logic;
signal \N__16404\ : std_logic;
signal \N__16401\ : std_logic;
signal \N__16398\ : std_logic;
signal \N__16397\ : std_logic;
signal \N__16396\ : std_logic;
signal \N__16391\ : std_logic;
signal \N__16388\ : std_logic;
signal \N__16385\ : std_logic;
signal \N__16380\ : std_logic;
signal \N__16377\ : std_logic;
signal \N__16374\ : std_logic;
signal \N__16371\ : std_logic;
signal \N__16368\ : std_logic;
signal \N__16365\ : std_logic;
signal \N__16362\ : std_logic;
signal \N__16357\ : std_logic;
signal \N__16356\ : std_logic;
signal \N__16353\ : std_logic;
signal \N__16350\ : std_logic;
signal \N__16345\ : std_logic;
signal \N__16342\ : std_logic;
signal \N__16341\ : std_logic;
signal \N__16338\ : std_logic;
signal \N__16335\ : std_logic;
signal \N__16330\ : std_logic;
signal \N__16327\ : std_logic;
signal \N__16326\ : std_logic;
signal \N__16323\ : std_logic;
signal \N__16320\ : std_logic;
signal \N__16315\ : std_logic;
signal \N__16312\ : std_logic;
signal \N__16311\ : std_logic;
signal \N__16308\ : std_logic;
signal \N__16305\ : std_logic;
signal \N__16300\ : std_logic;
signal \N__16297\ : std_logic;
signal \N__16296\ : std_logic;
signal \N__16293\ : std_logic;
signal \N__16290\ : std_logic;
signal \N__16285\ : std_logic;
signal \N__16282\ : std_logic;
signal \N__16279\ : std_logic;
signal \N__16278\ : std_logic;
signal \N__16275\ : std_logic;
signal \N__16272\ : std_logic;
signal \N__16267\ : std_logic;
signal \N__16266\ : std_logic;
signal \N__16263\ : std_logic;
signal \N__16260\ : std_logic;
signal \N__16257\ : std_logic;
signal \N__16254\ : std_logic;
signal \N__16251\ : std_logic;
signal \N__16248\ : std_logic;
signal \N__16243\ : std_logic;
signal \N__16240\ : std_logic;
signal \N__16237\ : std_logic;
signal \N__16234\ : std_logic;
signal \N__16231\ : std_logic;
signal \N__16228\ : std_logic;
signal \N__16225\ : std_logic;
signal \N__16222\ : std_logic;
signal \N__16219\ : std_logic;
signal \N__16216\ : std_logic;
signal \N__16215\ : std_logic;
signal \N__16212\ : std_logic;
signal \N__16209\ : std_logic;
signal \N__16206\ : std_logic;
signal \N__16203\ : std_logic;
signal \N__16200\ : std_logic;
signal \N__16197\ : std_logic;
signal \N__16194\ : std_logic;
signal \N__16191\ : std_logic;
signal \N__16188\ : std_logic;
signal \N__16185\ : std_logic;
signal \N__16182\ : std_logic;
signal \N__16179\ : std_logic;
signal \N__16176\ : std_logic;
signal \N__16173\ : std_logic;
signal \N__16170\ : std_logic;
signal \N__16167\ : std_logic;
signal \N__16164\ : std_logic;
signal \N__16161\ : std_logic;
signal \N__16158\ : std_logic;
signal \N__16155\ : std_logic;
signal \N__16152\ : std_logic;
signal \N__16149\ : std_logic;
signal \N__16146\ : std_logic;
signal \N__16143\ : std_logic;
signal \N__16140\ : std_logic;
signal \N__16137\ : std_logic;
signal \N__16134\ : std_logic;
signal \N__16131\ : std_logic;
signal \N__16128\ : std_logic;
signal \N__16125\ : std_logic;
signal \N__16122\ : std_logic;
signal \N__16119\ : std_logic;
signal \N__16116\ : std_logic;
signal \N__16113\ : std_logic;
signal \N__16110\ : std_logic;
signal \N__16107\ : std_logic;
signal \N__16104\ : std_logic;
signal \N__16101\ : std_logic;
signal \N__16098\ : std_logic;
signal \N__16095\ : std_logic;
signal \N__16092\ : std_logic;
signal \N__16089\ : std_logic;
signal \N__16086\ : std_logic;
signal \N__16083\ : std_logic;
signal \N__16080\ : std_logic;
signal \N__16077\ : std_logic;
signal \N__16074\ : std_logic;
signal \N__16071\ : std_logic;
signal \N__16068\ : std_logic;
signal \N__16065\ : std_logic;
signal \N__16062\ : std_logic;
signal \N__16059\ : std_logic;
signal \N__16056\ : std_logic;
signal \N__16053\ : std_logic;
signal \N__16050\ : std_logic;
signal \N__16047\ : std_logic;
signal \N__16044\ : std_logic;
signal \N__16041\ : std_logic;
signal \N__16038\ : std_logic;
signal \N__16035\ : std_logic;
signal \N__16032\ : std_logic;
signal \N__16029\ : std_logic;
signal \N__16026\ : std_logic;
signal \N__16023\ : std_logic;
signal \N__16020\ : std_logic;
signal \N__16017\ : std_logic;
signal \N__16014\ : std_logic;
signal \N__16011\ : std_logic;
signal \N__16010\ : std_logic;
signal \N__16007\ : std_logic;
signal \N__16004\ : std_logic;
signal \N__16001\ : std_logic;
signal \N__15998\ : std_logic;
signal \N__15995\ : std_logic;
signal \N__15994\ : std_logic;
signal \N__15991\ : std_logic;
signal \N__15986\ : std_logic;
signal \N__15983\ : std_logic;
signal \N__15978\ : std_logic;
signal \N__15973\ : std_logic;
signal \N__15970\ : std_logic;
signal \N__15967\ : std_logic;
signal \N__15964\ : std_logic;
signal \N__15961\ : std_logic;
signal \N__15958\ : std_logic;
signal \N__15957\ : std_logic;
signal \N__15954\ : std_logic;
signal \N__15951\ : std_logic;
signal \N__15948\ : std_logic;
signal \N__15945\ : std_logic;
signal \N__15942\ : std_logic;
signal \N__15939\ : std_logic;
signal \N__15936\ : std_logic;
signal \N__15933\ : std_logic;
signal \N__15930\ : std_logic;
signal \N__15927\ : std_logic;
signal \N__15924\ : std_logic;
signal \N__15921\ : std_logic;
signal \N__15918\ : std_logic;
signal \N__15915\ : std_logic;
signal \N__15912\ : std_logic;
signal \N__15909\ : std_logic;
signal \N__15906\ : std_logic;
signal \N__15903\ : std_logic;
signal \N__15900\ : std_logic;
signal \N__15897\ : std_logic;
signal \N__15894\ : std_logic;
signal \N__15891\ : std_logic;
signal \N__15888\ : std_logic;
signal \N__15885\ : std_logic;
signal \N__15882\ : std_logic;
signal \N__15879\ : std_logic;
signal \N__15876\ : std_logic;
signal \N__15873\ : std_logic;
signal \N__15870\ : std_logic;
signal \N__15867\ : std_logic;
signal \N__15864\ : std_logic;
signal \N__15861\ : std_logic;
signal \N__15858\ : std_logic;
signal \N__15855\ : std_logic;
signal \N__15852\ : std_logic;
signal \N__15849\ : std_logic;
signal \N__15846\ : std_logic;
signal \N__15843\ : std_logic;
signal \N__15840\ : std_logic;
signal \N__15837\ : std_logic;
signal \N__15834\ : std_logic;
signal \N__15831\ : std_logic;
signal \N__15828\ : std_logic;
signal \N__15825\ : std_logic;
signal \N__15822\ : std_logic;
signal \N__15819\ : std_logic;
signal \N__15816\ : std_logic;
signal \N__15813\ : std_logic;
signal \N__15810\ : std_logic;
signal \N__15807\ : std_logic;
signal \N__15804\ : std_logic;
signal \N__15801\ : std_logic;
signal \N__15798\ : std_logic;
signal \N__15795\ : std_logic;
signal \N__15792\ : std_logic;
signal \N__15789\ : std_logic;
signal \N__15786\ : std_logic;
signal \N__15783\ : std_logic;
signal \N__15780\ : std_logic;
signal \N__15777\ : std_logic;
signal \N__15774\ : std_logic;
signal \N__15771\ : std_logic;
signal \N__15768\ : std_logic;
signal \N__15765\ : std_logic;
signal \N__15762\ : std_logic;
signal \N__15759\ : std_logic;
signal \N__15758\ : std_logic;
signal \N__15755\ : std_logic;
signal \N__15752\ : std_logic;
signal \N__15751\ : std_logic;
signal \N__15748\ : std_logic;
signal \N__15745\ : std_logic;
signal \N__15742\ : std_logic;
signal \N__15739\ : std_logic;
signal \N__15736\ : std_logic;
signal \N__15733\ : std_logic;
signal \N__15730\ : std_logic;
signal \N__15725\ : std_logic;
signal \N__15720\ : std_logic;
signal \N__15715\ : std_logic;
signal \N__15712\ : std_logic;
signal \N__15709\ : std_logic;
signal \N__15706\ : std_logic;
signal \N__15703\ : std_logic;
signal \N__15700\ : std_logic;
signal \N__15697\ : std_logic;
signal \N__15694\ : std_logic;
signal \N__15691\ : std_logic;
signal \N__15688\ : std_logic;
signal \N__15685\ : std_logic;
signal \N__15682\ : std_logic;
signal \N__15679\ : std_logic;
signal \N__15676\ : std_logic;
signal \N__15673\ : std_logic;
signal \N__15670\ : std_logic;
signal \N__15667\ : std_logic;
signal \N__15664\ : std_logic;
signal \N__15661\ : std_logic;
signal \N__15658\ : std_logic;
signal \N__15657\ : std_logic;
signal \N__15654\ : std_logic;
signal \N__15651\ : std_logic;
signal \N__15648\ : std_logic;
signal \N__15645\ : std_logic;
signal \N__15642\ : std_logic;
signal \N__15639\ : std_logic;
signal \N__15636\ : std_logic;
signal \N__15633\ : std_logic;
signal \N__15630\ : std_logic;
signal \N__15627\ : std_logic;
signal \N__15624\ : std_logic;
signal \N__15621\ : std_logic;
signal \N__15618\ : std_logic;
signal \N__15615\ : std_logic;
signal \N__15612\ : std_logic;
signal \N__15609\ : std_logic;
signal \N__15606\ : std_logic;
signal \N__15603\ : std_logic;
signal \N__15600\ : std_logic;
signal \N__15597\ : std_logic;
signal \N__15594\ : std_logic;
signal \N__15591\ : std_logic;
signal \N__15588\ : std_logic;
signal \N__15585\ : std_logic;
signal \N__15582\ : std_logic;
signal \N__15579\ : std_logic;
signal \N__15576\ : std_logic;
signal \N__15573\ : std_logic;
signal \N__15570\ : std_logic;
signal \N__15567\ : std_logic;
signal \N__15564\ : std_logic;
signal \N__15561\ : std_logic;
signal \N__15558\ : std_logic;
signal \N__15555\ : std_logic;
signal \N__15552\ : std_logic;
signal \N__15549\ : std_logic;
signal \N__15546\ : std_logic;
signal \N__15543\ : std_logic;
signal \N__15540\ : std_logic;
signal \N__15537\ : std_logic;
signal \N__15534\ : std_logic;
signal \N__15531\ : std_logic;
signal \N__15528\ : std_logic;
signal \N__15525\ : std_logic;
signal \N__15522\ : std_logic;
signal \N__15519\ : std_logic;
signal \N__15516\ : std_logic;
signal \N__15513\ : std_logic;
signal \N__15510\ : std_logic;
signal \N__15507\ : std_logic;
signal \N__15504\ : std_logic;
signal \N__15501\ : std_logic;
signal \N__15498\ : std_logic;
signal \N__15495\ : std_logic;
signal \N__15492\ : std_logic;
signal \N__15489\ : std_logic;
signal \N__15486\ : std_logic;
signal \N__15483\ : std_logic;
signal \N__15480\ : std_logic;
signal \N__15479\ : std_logic;
signal \N__15476\ : std_logic;
signal \N__15473\ : std_logic;
signal \N__15470\ : std_logic;
signal \N__15467\ : std_logic;
signal \N__15464\ : std_logic;
signal \N__15461\ : std_logic;
signal \N__15458\ : std_logic;
signal \N__15455\ : std_logic;
signal \N__15452\ : std_logic;
signal \N__15449\ : std_logic;
signal \N__15446\ : std_logic;
signal \N__15443\ : std_logic;
signal \N__15442\ : std_logic;
signal \N__15439\ : std_logic;
signal \N__15436\ : std_logic;
signal \N__15433\ : std_logic;
signal \N__15430\ : std_logic;
signal \N__15427\ : std_logic;
signal \N__15424\ : std_logic;
signal \N__15415\ : std_logic;
signal \N__15412\ : std_logic;
signal \N__15409\ : std_logic;
signal \N__15406\ : std_logic;
signal \N__15403\ : std_logic;
signal \N__15400\ : std_logic;
signal \N__15399\ : std_logic;
signal \N__15396\ : std_logic;
signal \N__15393\ : std_logic;
signal \N__15390\ : std_logic;
signal \N__15387\ : std_logic;
signal \N__15384\ : std_logic;
signal \N__15381\ : std_logic;
signal \N__15378\ : std_logic;
signal \N__15375\ : std_logic;
signal \N__15372\ : std_logic;
signal \N__15369\ : std_logic;
signal \N__15366\ : std_logic;
signal \N__15363\ : std_logic;
signal \N__15360\ : std_logic;
signal \N__15357\ : std_logic;
signal \N__15354\ : std_logic;
signal \N__15351\ : std_logic;
signal \N__15348\ : std_logic;
signal \N__15345\ : std_logic;
signal \N__15342\ : std_logic;
signal \N__15339\ : std_logic;
signal \N__15336\ : std_logic;
signal \N__15333\ : std_logic;
signal \N__15330\ : std_logic;
signal \N__15327\ : std_logic;
signal \N__15324\ : std_logic;
signal \N__15321\ : std_logic;
signal \N__15318\ : std_logic;
signal \N__15315\ : std_logic;
signal \N__15312\ : std_logic;
signal \N__15309\ : std_logic;
signal \N__15306\ : std_logic;
signal \N__15303\ : std_logic;
signal \N__15300\ : std_logic;
signal \N__15297\ : std_logic;
signal \N__15294\ : std_logic;
signal \N__15291\ : std_logic;
signal \N__15288\ : std_logic;
signal \N__15285\ : std_logic;
signal \N__15282\ : std_logic;
signal \N__15279\ : std_logic;
signal \N__15276\ : std_logic;
signal \N__15273\ : std_logic;
signal \N__15270\ : std_logic;
signal \N__15267\ : std_logic;
signal \N__15264\ : std_logic;
signal \N__15261\ : std_logic;
signal \N__15258\ : std_logic;
signal \N__15255\ : std_logic;
signal \N__15252\ : std_logic;
signal \N__15249\ : std_logic;
signal \N__15246\ : std_logic;
signal \N__15243\ : std_logic;
signal \N__15240\ : std_logic;
signal \N__15237\ : std_logic;
signal \N__15234\ : std_logic;
signal \N__15231\ : std_logic;
signal \N__15228\ : std_logic;
signal \N__15225\ : std_logic;
signal \N__15222\ : std_logic;
signal \N__15219\ : std_logic;
signal \N__15218\ : std_logic;
signal \N__15215\ : std_logic;
signal \N__15212\ : std_logic;
signal \N__15209\ : std_logic;
signal \N__15206\ : std_logic;
signal \N__15203\ : std_logic;
signal \N__15202\ : std_logic;
signal \N__15199\ : std_logic;
signal \N__15196\ : std_logic;
signal \N__15193\ : std_logic;
signal \N__15190\ : std_logic;
signal \N__15183\ : std_logic;
signal \N__15178\ : std_logic;
signal \N__15175\ : std_logic;
signal \N__15172\ : std_logic;
signal \N__15169\ : std_logic;
signal \N__15166\ : std_logic;
signal \N__15163\ : std_logic;
signal \N__15162\ : std_logic;
signal \N__15159\ : std_logic;
signal \N__15156\ : std_logic;
signal \N__15153\ : std_logic;
signal \N__15150\ : std_logic;
signal \N__15147\ : std_logic;
signal \N__15144\ : std_logic;
signal \N__15141\ : std_logic;
signal \N__15138\ : std_logic;
signal \N__15135\ : std_logic;
signal \N__15132\ : std_logic;
signal \N__15129\ : std_logic;
signal \N__15126\ : std_logic;
signal \N__15123\ : std_logic;
signal \N__15120\ : std_logic;
signal \N__15117\ : std_logic;
signal \N__15114\ : std_logic;
signal \N__15111\ : std_logic;
signal \N__15108\ : std_logic;
signal \N__15105\ : std_logic;
signal \N__15102\ : std_logic;
signal \N__15099\ : std_logic;
signal \N__15096\ : std_logic;
signal \N__15093\ : std_logic;
signal \N__15090\ : std_logic;
signal \N__15087\ : std_logic;
signal \N__15084\ : std_logic;
signal \N__15081\ : std_logic;
signal \N__15078\ : std_logic;
signal \N__15075\ : std_logic;
signal \N__15072\ : std_logic;
signal \N__15069\ : std_logic;
signal \N__15066\ : std_logic;
signal \N__15063\ : std_logic;
signal \N__15060\ : std_logic;
signal \N__15057\ : std_logic;
signal \N__15054\ : std_logic;
signal \N__15051\ : std_logic;
signal \N__15048\ : std_logic;
signal \N__15045\ : std_logic;
signal \N__15042\ : std_logic;
signal \N__15039\ : std_logic;
signal \N__15036\ : std_logic;
signal \N__15033\ : std_logic;
signal \N__15030\ : std_logic;
signal \N__15027\ : std_logic;
signal \N__15024\ : std_logic;
signal \N__15021\ : std_logic;
signal \N__15018\ : std_logic;
signal \N__15015\ : std_logic;
signal \N__15012\ : std_logic;
signal \N__15009\ : std_logic;
signal \N__15006\ : std_logic;
signal \N__15003\ : std_logic;
signal \N__15000\ : std_logic;
signal \N__14997\ : std_logic;
signal \N__14994\ : std_logic;
signal \N__14991\ : std_logic;
signal \N__14990\ : std_logic;
signal \N__14987\ : std_logic;
signal \N__14984\ : std_logic;
signal \N__14981\ : std_logic;
signal \N__14978\ : std_logic;
signal \N__14975\ : std_logic;
signal \N__14972\ : std_logic;
signal \N__14969\ : std_logic;
signal \N__14966\ : std_logic;
signal \N__14963\ : std_logic;
signal \N__14960\ : std_logic;
signal \N__14957\ : std_logic;
signal \N__14956\ : std_logic;
signal \N__14953\ : std_logic;
signal \N__14950\ : std_logic;
signal \N__14947\ : std_logic;
signal \N__14944\ : std_logic;
signal \N__14941\ : std_logic;
signal \N__14938\ : std_logic;
signal \N__14935\ : std_logic;
signal \N__14932\ : std_logic;
signal \N__14929\ : std_logic;
signal \N__14926\ : std_logic;
signal \N__14923\ : std_logic;
signal \N__14914\ : std_logic;
signal \N__14911\ : std_logic;
signal \N__14908\ : std_logic;
signal \N__14905\ : std_logic;
signal \N__14902\ : std_logic;
signal \N__14899\ : std_logic;
signal \N__14896\ : std_logic;
signal \N__14895\ : std_logic;
signal \N__14892\ : std_logic;
signal \N__14889\ : std_logic;
signal \N__14886\ : std_logic;
signal \N__14883\ : std_logic;
signal \N__14880\ : std_logic;
signal \N__14877\ : std_logic;
signal \N__14874\ : std_logic;
signal \N__14871\ : std_logic;
signal \N__14868\ : std_logic;
signal \N__14865\ : std_logic;
signal \N__14862\ : std_logic;
signal \N__14859\ : std_logic;
signal \N__14856\ : std_logic;
signal \N__14853\ : std_logic;
signal \N__14850\ : std_logic;
signal \N__14847\ : std_logic;
signal \N__14844\ : std_logic;
signal \N__14841\ : std_logic;
signal \N__14838\ : std_logic;
signal \N__14835\ : std_logic;
signal \N__14832\ : std_logic;
signal \N__14829\ : std_logic;
signal \N__14826\ : std_logic;
signal \N__14823\ : std_logic;
signal \N__14820\ : std_logic;
signal \N__14817\ : std_logic;
signal \N__14814\ : std_logic;
signal \N__14811\ : std_logic;
signal \N__14808\ : std_logic;
signal \N__14805\ : std_logic;
signal \N__14802\ : std_logic;
signal \N__14799\ : std_logic;
signal \N__14796\ : std_logic;
signal \N__14793\ : std_logic;
signal \N__14790\ : std_logic;
signal \N__14787\ : std_logic;
signal \N__14784\ : std_logic;
signal \N__14781\ : std_logic;
signal \N__14778\ : std_logic;
signal \N__14775\ : std_logic;
signal \N__14772\ : std_logic;
signal \N__14769\ : std_logic;
signal \N__14766\ : std_logic;
signal \N__14763\ : std_logic;
signal \N__14760\ : std_logic;
signal \N__14757\ : std_logic;
signal \N__14754\ : std_logic;
signal \N__14751\ : std_logic;
signal \N__14748\ : std_logic;
signal \N__14745\ : std_logic;
signal \N__14742\ : std_logic;
signal \N__14739\ : std_logic;
signal \N__14736\ : std_logic;
signal \N__14733\ : std_logic;
signal \N__14730\ : std_logic;
signal \N__14727\ : std_logic;
signal \N__14724\ : std_logic;
signal \N__14721\ : std_logic;
signal \N__14718\ : std_logic;
signal \N__14715\ : std_logic;
signal \N__14714\ : std_logic;
signal \N__14711\ : std_logic;
signal \N__14708\ : std_logic;
signal \N__14705\ : std_logic;
signal \N__14702\ : std_logic;
signal \N__14699\ : std_logic;
signal \N__14696\ : std_logic;
signal \N__14693\ : std_logic;
signal \N__14690\ : std_logic;
signal \N__14687\ : std_logic;
signal \N__14686\ : std_logic;
signal \N__14683\ : std_logic;
signal \N__14680\ : std_logic;
signal \N__14677\ : std_logic;
signal \N__14674\ : std_logic;
signal \N__14669\ : std_logic;
signal \N__14662\ : std_logic;
signal \N__14659\ : std_logic;
signal \N__14656\ : std_logic;
signal \N__14653\ : std_logic;
signal \N__14650\ : std_logic;
signal \N__14647\ : std_logic;
signal \N__14646\ : std_logic;
signal \N__14643\ : std_logic;
signal \N__14640\ : std_logic;
signal \N__14637\ : std_logic;
signal \N__14634\ : std_logic;
signal \N__14631\ : std_logic;
signal \N__14628\ : std_logic;
signal \N__14625\ : std_logic;
signal \N__14622\ : std_logic;
signal \N__14619\ : std_logic;
signal \N__14616\ : std_logic;
signal \N__14613\ : std_logic;
signal \N__14610\ : std_logic;
signal \N__14607\ : std_logic;
signal \N__14604\ : std_logic;
signal \N__14601\ : std_logic;
signal \N__14598\ : std_logic;
signal \N__14595\ : std_logic;
signal \N__14592\ : std_logic;
signal \N__14589\ : std_logic;
signal \N__14586\ : std_logic;
signal \N__14583\ : std_logic;
signal \N__14580\ : std_logic;
signal \N__14577\ : std_logic;
signal \N__14574\ : std_logic;
signal \N__14571\ : std_logic;
signal \N__14568\ : std_logic;
signal \N__14565\ : std_logic;
signal \N__14562\ : std_logic;
signal \N__14559\ : std_logic;
signal \N__14556\ : std_logic;
signal \N__14553\ : std_logic;
signal \N__14550\ : std_logic;
signal \N__14547\ : std_logic;
signal \N__14544\ : std_logic;
signal \N__14541\ : std_logic;
signal \N__14538\ : std_logic;
signal \N__14535\ : std_logic;
signal \N__14532\ : std_logic;
signal \N__14529\ : std_logic;
signal \N__14526\ : std_logic;
signal \N__14523\ : std_logic;
signal \N__14520\ : std_logic;
signal \N__14517\ : std_logic;
signal \N__14514\ : std_logic;
signal \N__14511\ : std_logic;
signal \N__14508\ : std_logic;
signal \N__14505\ : std_logic;
signal \N__14502\ : std_logic;
signal \N__14499\ : std_logic;
signal \N__14496\ : std_logic;
signal \N__14493\ : std_logic;
signal \N__14490\ : std_logic;
signal \N__14487\ : std_logic;
signal \N__14484\ : std_logic;
signal \N__14481\ : std_logic;
signal \N__14478\ : std_logic;
signal \N__14475\ : std_logic;
signal \N__14472\ : std_logic;
signal \N__14469\ : std_logic;
signal \N__14466\ : std_logic;
signal \N__14463\ : std_logic;
signal \N__14462\ : std_logic;
signal \N__14459\ : std_logic;
signal \N__14456\ : std_logic;
signal \N__14453\ : std_logic;
signal \N__14450\ : std_logic;
signal \N__14447\ : std_logic;
signal \N__14446\ : std_logic;
signal \N__14443\ : std_logic;
signal \N__14440\ : std_logic;
signal \N__14437\ : std_logic;
signal \N__14434\ : std_logic;
signal \N__14431\ : std_logic;
signal \N__14428\ : std_logic;
signal \N__14425\ : std_logic;
signal \N__14422\ : std_logic;
signal \N__14419\ : std_logic;
signal \N__14414\ : std_logic;
signal \N__14407\ : std_logic;
signal \N__14404\ : std_logic;
signal \N__14401\ : std_logic;
signal \N__14398\ : std_logic;
signal \N__14395\ : std_logic;
signal \N__14392\ : std_logic;
signal \N__14391\ : std_logic;
signal \N__14388\ : std_logic;
signal \N__14385\ : std_logic;
signal \N__14382\ : std_logic;
signal \N__14379\ : std_logic;
signal \N__14376\ : std_logic;
signal \N__14373\ : std_logic;
signal \N__14370\ : std_logic;
signal \N__14367\ : std_logic;
signal \N__14364\ : std_logic;
signal \N__14361\ : std_logic;
signal \N__14358\ : std_logic;
signal \N__14355\ : std_logic;
signal \N__14352\ : std_logic;
signal \N__14349\ : std_logic;
signal \N__14346\ : std_logic;
signal \N__14343\ : std_logic;
signal \N__14340\ : std_logic;
signal \N__14337\ : std_logic;
signal \N__14334\ : std_logic;
signal \N__14331\ : std_logic;
signal \N__14328\ : std_logic;
signal \N__14325\ : std_logic;
signal \N__14322\ : std_logic;
signal \N__14319\ : std_logic;
signal \N__14316\ : std_logic;
signal \N__14313\ : std_logic;
signal \N__14310\ : std_logic;
signal \N__14307\ : std_logic;
signal \N__14304\ : std_logic;
signal \N__14301\ : std_logic;
signal \N__14298\ : std_logic;
signal \N__14295\ : std_logic;
signal \N__14292\ : std_logic;
signal \N__14289\ : std_logic;
signal \N__14286\ : std_logic;
signal \N__14283\ : std_logic;
signal \N__14280\ : std_logic;
signal \N__14277\ : std_logic;
signal \N__14274\ : std_logic;
signal \N__14271\ : std_logic;
signal \N__14268\ : std_logic;
signal \N__14265\ : std_logic;
signal \N__14262\ : std_logic;
signal \N__14259\ : std_logic;
signal \N__14256\ : std_logic;
signal \N__14253\ : std_logic;
signal \N__14250\ : std_logic;
signal \N__14247\ : std_logic;
signal \N__14244\ : std_logic;
signal \N__14241\ : std_logic;
signal \N__14238\ : std_logic;
signal \N__14235\ : std_logic;
signal \N__14232\ : std_logic;
signal \N__14229\ : std_logic;
signal \N__14226\ : std_logic;
signal \N__14223\ : std_logic;
signal \N__14220\ : std_logic;
signal \N__14217\ : std_logic;
signal \N__14214\ : std_logic;
signal \N__14211\ : std_logic;
signal \N__14210\ : std_logic;
signal \N__14207\ : std_logic;
signal \N__14204\ : std_logic;
signal \N__14201\ : std_logic;
signal \N__14198\ : std_logic;
signal \N__14195\ : std_logic;
signal \N__14192\ : std_logic;
signal \N__14189\ : std_logic;
signal \N__14186\ : std_logic;
signal \N__14183\ : std_logic;
signal \N__14182\ : std_logic;
signal \N__14179\ : std_logic;
signal \N__14176\ : std_logic;
signal \N__14173\ : std_logic;
signal \N__14170\ : std_logic;
signal \N__14165\ : std_logic;
signal \N__14158\ : std_logic;
signal \N__14155\ : std_logic;
signal \N__14152\ : std_logic;
signal \N__14149\ : std_logic;
signal \N__14146\ : std_logic;
signal \N__14143\ : std_logic;
signal \N__14140\ : std_logic;
signal \N__14139\ : std_logic;
signal \N__14136\ : std_logic;
signal \N__14133\ : std_logic;
signal \N__14130\ : std_logic;
signal \N__14127\ : std_logic;
signal \N__14124\ : std_logic;
signal \N__14121\ : std_logic;
signal \N__14118\ : std_logic;
signal \N__14115\ : std_logic;
signal \N__14112\ : std_logic;
signal \N__14109\ : std_logic;
signal \N__14106\ : std_logic;
signal \N__14103\ : std_logic;
signal \N__14100\ : std_logic;
signal \N__14097\ : std_logic;
signal \N__14094\ : std_logic;
signal \N__14091\ : std_logic;
signal \N__14088\ : std_logic;
signal \N__14085\ : std_logic;
signal \N__14082\ : std_logic;
signal \N__14079\ : std_logic;
signal \N__14076\ : std_logic;
signal \N__14073\ : std_logic;
signal \N__14070\ : std_logic;
signal \N__14067\ : std_logic;
signal \N__14064\ : std_logic;
signal \N__14061\ : std_logic;
signal \N__14058\ : std_logic;
signal \N__14055\ : std_logic;
signal \N__14052\ : std_logic;
signal \N__14049\ : std_logic;
signal \N__14046\ : std_logic;
signal \N__14043\ : std_logic;
signal \N__14040\ : std_logic;
signal \N__14037\ : std_logic;
signal \N__14034\ : std_logic;
signal \N__14031\ : std_logic;
signal \N__14028\ : std_logic;
signal \N__14025\ : std_logic;
signal \N__14022\ : std_logic;
signal \N__14019\ : std_logic;
signal \N__14016\ : std_logic;
signal \N__14013\ : std_logic;
signal \N__14010\ : std_logic;
signal \N__14007\ : std_logic;
signal \N__14004\ : std_logic;
signal \N__14001\ : std_logic;
signal \N__13998\ : std_logic;
signal \N__13995\ : std_logic;
signal \N__13992\ : std_logic;
signal \N__13989\ : std_logic;
signal \N__13986\ : std_logic;
signal \N__13983\ : std_logic;
signal \N__13980\ : std_logic;
signal \N__13977\ : std_logic;
signal \N__13976\ : std_logic;
signal \N__13973\ : std_logic;
signal \N__13970\ : std_logic;
signal \N__13967\ : std_logic;
signal \N__13964\ : std_logic;
signal \N__13961\ : std_logic;
signal \N__13958\ : std_logic;
signal \N__13955\ : std_logic;
signal \N__13952\ : std_logic;
signal \N__13949\ : std_logic;
signal \N__13946\ : std_logic;
signal \N__13943\ : std_logic;
signal \N__13942\ : std_logic;
signal \N__13939\ : std_logic;
signal \N__13936\ : std_logic;
signal \N__13933\ : std_logic;
signal \N__13930\ : std_logic;
signal \N__13927\ : std_logic;
signal \N__13924\ : std_logic;
signal \N__13921\ : std_logic;
signal \N__13918\ : std_logic;
signal \N__13915\ : std_logic;
signal \N__13912\ : std_logic;
signal \N__13909\ : std_logic;
signal \N__13900\ : std_logic;
signal \N__13897\ : std_logic;
signal \N__13894\ : std_logic;
signal \N__13891\ : std_logic;
signal \N__13888\ : std_logic;
signal \N__13885\ : std_logic;
signal \N__13882\ : std_logic;
signal \N__13879\ : std_logic;
signal \N__13876\ : std_logic;
signal \N__13873\ : std_logic;
signal \N__13870\ : std_logic;
signal \N__13867\ : std_logic;
signal \N__13864\ : std_logic;
signal \N__13861\ : std_logic;
signal \N__13858\ : std_logic;
signal \N__13855\ : std_logic;
signal \N__13852\ : std_logic;
signal \N__13849\ : std_logic;
signal \N__13846\ : std_logic;
signal \N__13843\ : std_logic;
signal \N__13842\ : std_logic;
signal \N__13839\ : std_logic;
signal \N__13836\ : std_logic;
signal \N__13833\ : std_logic;
signal \N__13830\ : std_logic;
signal \N__13827\ : std_logic;
signal \N__13822\ : std_logic;
signal \N__13819\ : std_logic;
signal \N__13816\ : std_logic;
signal \N__13813\ : std_logic;
signal \N__13810\ : std_logic;
signal \N__13807\ : std_logic;
signal \N__13804\ : std_logic;
signal \N__13801\ : std_logic;
signal \N__13798\ : std_logic;
signal \N__13795\ : std_logic;
signal \N__13792\ : std_logic;
signal \N__13789\ : std_logic;
signal \N__13786\ : std_logic;
signal \N__13783\ : std_logic;
signal \N__13782\ : std_logic;
signal \N__13779\ : std_logic;
signal \N__13776\ : std_logic;
signal \N__13773\ : std_logic;
signal \N__13770\ : std_logic;
signal \N__13767\ : std_logic;
signal \N__13764\ : std_logic;
signal \N__13761\ : std_logic;
signal \N__13758\ : std_logic;
signal \N__13755\ : std_logic;
signal \N__13752\ : std_logic;
signal \N__13749\ : std_logic;
signal \N__13746\ : std_logic;
signal \N__13743\ : std_logic;
signal \N__13740\ : std_logic;
signal \N__13737\ : std_logic;
signal \N__13734\ : std_logic;
signal \N__13731\ : std_logic;
signal \N__13728\ : std_logic;
signal \N__13725\ : std_logic;
signal \N__13722\ : std_logic;
signal \N__13719\ : std_logic;
signal \N__13716\ : std_logic;
signal \N__13713\ : std_logic;
signal \N__13710\ : std_logic;
signal \N__13707\ : std_logic;
signal \N__13704\ : std_logic;
signal \N__13701\ : std_logic;
signal \N__13698\ : std_logic;
signal \N__13695\ : std_logic;
signal \N__13692\ : std_logic;
signal \N__13689\ : std_logic;
signal \N__13686\ : std_logic;
signal \N__13683\ : std_logic;
signal \N__13680\ : std_logic;
signal \N__13677\ : std_logic;
signal \N__13674\ : std_logic;
signal \N__13671\ : std_logic;
signal \N__13668\ : std_logic;
signal \N__13665\ : std_logic;
signal \N__13662\ : std_logic;
signal \N__13659\ : std_logic;
signal \N__13656\ : std_logic;
signal \N__13653\ : std_logic;
signal \N__13650\ : std_logic;
signal \N__13647\ : std_logic;
signal \N__13644\ : std_logic;
signal \N__13641\ : std_logic;
signal \N__13638\ : std_logic;
signal \N__13635\ : std_logic;
signal \N__13632\ : std_logic;
signal \N__13629\ : std_logic;
signal \N__13626\ : std_logic;
signal \N__13623\ : std_logic;
signal \N__13620\ : std_logic;
signal \N__13617\ : std_logic;
signal \N__13614\ : std_logic;
signal \N__13611\ : std_logic;
signal \N__13608\ : std_logic;
signal \N__13605\ : std_logic;
signal \N__13602\ : std_logic;
signal \N__13599\ : std_logic;
signal \N__13596\ : std_logic;
signal \N__13593\ : std_logic;
signal \N__13590\ : std_logic;
signal \N__13589\ : std_logic;
signal \N__13586\ : std_logic;
signal \N__13583\ : std_logic;
signal \N__13580\ : std_logic;
signal \N__13577\ : std_logic;
signal \N__13574\ : std_logic;
signal \N__13571\ : std_logic;
signal \N__13570\ : std_logic;
signal \N__13567\ : std_logic;
signal \N__13564\ : std_logic;
signal \N__13561\ : std_logic;
signal \N__13558\ : std_logic;
signal \N__13553\ : std_logic;
signal \N__13546\ : std_logic;
signal \N__13545\ : std_logic;
signal \N__13544\ : std_logic;
signal \N__13543\ : std_logic;
signal \N__13540\ : std_logic;
signal \N__13537\ : std_logic;
signal \N__13534\ : std_logic;
signal \N__13531\ : std_logic;
signal \N__13528\ : std_logic;
signal \N__13525\ : std_logic;
signal \N__13522\ : std_logic;
signal \N__13513\ : std_logic;
signal \N__13510\ : std_logic;
signal \N__13507\ : std_logic;
signal \N__13504\ : std_logic;
signal \N__13501\ : std_logic;
signal \N__13498\ : std_logic;
signal \N__13497\ : std_logic;
signal \N__13496\ : std_logic;
signal \N__13495\ : std_logic;
signal \N__13492\ : std_logic;
signal \N__13487\ : std_logic;
signal \N__13484\ : std_logic;
signal \N__13477\ : std_logic;
signal \N__13474\ : std_logic;
signal \N__13471\ : std_logic;
signal \N__13468\ : std_logic;
signal \N__13465\ : std_logic;
signal \N__13462\ : std_logic;
signal \N__13459\ : std_logic;
signal \N__13456\ : std_logic;
signal \N__13455\ : std_logic;
signal \N__13454\ : std_logic;
signal \N__13451\ : std_logic;
signal \N__13448\ : std_logic;
signal \N__13445\ : std_logic;
signal \N__13440\ : std_logic;
signal \N__13439\ : std_logic;
signal \N__13434\ : std_logic;
signal \N__13431\ : std_logic;
signal \N__13426\ : std_logic;
signal \N__13423\ : std_logic;
signal \N__13422\ : std_logic;
signal \N__13419\ : std_logic;
signal \N__13416\ : std_logic;
signal \N__13413\ : std_logic;
signal \N__13410\ : std_logic;
signal \N__13407\ : std_logic;
signal \N__13404\ : std_logic;
signal \N__13399\ : std_logic;
signal \N__13396\ : std_logic;
signal \N__13393\ : std_logic;
signal \N__13390\ : std_logic;
signal \N__13389\ : std_logic;
signal \N__13386\ : std_logic;
signal \N__13385\ : std_logic;
signal \N__13384\ : std_logic;
signal \N__13381\ : std_logic;
signal \N__13378\ : std_logic;
signal \N__13373\ : std_logic;
signal \N__13370\ : std_logic;
signal \N__13363\ : std_logic;
signal \N__13360\ : std_logic;
signal \N__13357\ : std_logic;
signal \N__13354\ : std_logic;
signal \N__13351\ : std_logic;
signal \N__13348\ : std_logic;
signal \N__13345\ : std_logic;
signal \N__13342\ : std_logic;
signal \N__13339\ : std_logic;
signal \N__13338\ : std_logic;
signal \N__13337\ : std_logic;
signal \N__13336\ : std_logic;
signal \N__13333\ : std_logic;
signal \N__13330\ : std_logic;
signal \N__13327\ : std_logic;
signal \N__13324\ : std_logic;
signal \N__13315\ : std_logic;
signal \N__13312\ : std_logic;
signal \N__13309\ : std_logic;
signal \N__13306\ : std_logic;
signal \N__13305\ : std_logic;
signal \N__13304\ : std_logic;
signal \N__13301\ : std_logic;
signal \N__13298\ : std_logic;
signal \N__13297\ : std_logic;
signal \N__13294\ : std_logic;
signal \N__13289\ : std_logic;
signal \N__13286\ : std_logic;
signal \N__13283\ : std_logic;
signal \N__13276\ : std_logic;
signal \N__13273\ : std_logic;
signal \N__13270\ : std_logic;
signal \N__13267\ : std_logic;
signal \N__13266\ : std_logic;
signal \N__13265\ : std_logic;
signal \N__13262\ : std_logic;
signal \N__13259\ : std_logic;
signal \N__13258\ : std_logic;
signal \N__13255\ : std_logic;
signal \N__13252\ : std_logic;
signal \N__13249\ : std_logic;
signal \N__13246\ : std_logic;
signal \N__13243\ : std_logic;
signal \N__13234\ : std_logic;
signal \N__13231\ : std_logic;
signal \N__13228\ : std_logic;
signal \N__13225\ : std_logic;
signal \N__13222\ : std_logic;
signal \N__13219\ : std_logic;
signal \N__13216\ : std_logic;
signal \N__13213\ : std_logic;
signal \N__13210\ : std_logic;
signal \N__13207\ : std_logic;
signal \N__13204\ : std_logic;
signal \N__13201\ : std_logic;
signal \N__13198\ : std_logic;
signal \N__13195\ : std_logic;
signal \N__13192\ : std_logic;
signal \N__13189\ : std_logic;
signal \N__13186\ : std_logic;
signal \N__13183\ : std_logic;
signal \N__13180\ : std_logic;
signal \N__13177\ : std_logic;
signal \N__13174\ : std_logic;
signal \N__13171\ : std_logic;
signal \N__13168\ : std_logic;
signal \N__13165\ : std_logic;
signal \N__13164\ : std_logic;
signal \N__13161\ : std_logic;
signal \N__13160\ : std_logic;
signal \N__13159\ : std_logic;
signal \N__13156\ : std_logic;
signal \N__13153\ : std_logic;
signal \N__13148\ : std_logic;
signal \N__13141\ : std_logic;
signal \N__13140\ : std_logic;
signal \N__13137\ : std_logic;
signal \N__13134\ : std_logic;
signal \N__13129\ : std_logic;
signal \N__13126\ : std_logic;
signal \N__13123\ : std_logic;
signal \N__13122\ : std_logic;
signal \N__13121\ : std_logic;
signal \N__13120\ : std_logic;
signal \N__13117\ : std_logic;
signal \N__13114\ : std_logic;
signal \N__13109\ : std_logic;
signal \N__13102\ : std_logic;
signal \N__13099\ : std_logic;
signal \N__13096\ : std_logic;
signal \N__13093\ : std_logic;
signal \N__13092\ : std_logic;
signal \N__13089\ : std_logic;
signal \N__13086\ : std_logic;
signal \N__13083\ : std_logic;
signal \N__13080\ : std_logic;
signal \N__13075\ : std_logic;
signal \N__13072\ : std_logic;
signal \N__13069\ : std_logic;
signal \N__13066\ : std_logic;
signal \N__13063\ : std_logic;
signal \N__13060\ : std_logic;
signal \N__13057\ : std_logic;
signal \N__13054\ : std_logic;
signal \N__13053\ : std_logic;
signal \N__13050\ : std_logic;
signal \N__13047\ : std_logic;
signal \N__13044\ : std_logic;
signal \N__13041\ : std_logic;
signal \N__13038\ : std_logic;
signal \N__13033\ : std_logic;
signal \N__13030\ : std_logic;
signal \N__13027\ : std_logic;
signal \N__13024\ : std_logic;
signal \N__13021\ : std_logic;
signal \N__13018\ : std_logic;
signal \N__13015\ : std_logic;
signal \N__13014\ : std_logic;
signal \N__13011\ : std_logic;
signal \N__13008\ : std_logic;
signal \N__13005\ : std_logic;
signal \N__13002\ : std_logic;
signal \N__12999\ : std_logic;
signal \N__12996\ : std_logic;
signal \N__12993\ : std_logic;
signal \N__12990\ : std_logic;
signal \N__12987\ : std_logic;
signal \N__12984\ : std_logic;
signal \N__12981\ : std_logic;
signal \N__12978\ : std_logic;
signal \N__12975\ : std_logic;
signal \N__12972\ : std_logic;
signal \N__12969\ : std_logic;
signal \N__12966\ : std_logic;
signal \N__12963\ : std_logic;
signal \N__12960\ : std_logic;
signal \N__12957\ : std_logic;
signal \N__12954\ : std_logic;
signal \N__12951\ : std_logic;
signal \N__12948\ : std_logic;
signal \N__12945\ : std_logic;
signal \N__12942\ : std_logic;
signal \N__12939\ : std_logic;
signal \N__12936\ : std_logic;
signal \N__12933\ : std_logic;
signal \N__12930\ : std_logic;
signal \N__12927\ : std_logic;
signal \N__12924\ : std_logic;
signal \N__12921\ : std_logic;
signal \N__12918\ : std_logic;
signal \N__12915\ : std_logic;
signal \N__12912\ : std_logic;
signal \N__12909\ : std_logic;
signal \N__12906\ : std_logic;
signal \N__12903\ : std_logic;
signal \N__12900\ : std_logic;
signal \N__12897\ : std_logic;
signal \N__12894\ : std_logic;
signal \N__12891\ : std_logic;
signal \N__12888\ : std_logic;
signal \N__12885\ : std_logic;
signal \N__12882\ : std_logic;
signal \N__12879\ : std_logic;
signal \N__12876\ : std_logic;
signal \N__12873\ : std_logic;
signal \N__12870\ : std_logic;
signal \N__12867\ : std_logic;
signal \N__12864\ : std_logic;
signal \N__12861\ : std_logic;
signal \N__12858\ : std_logic;
signal \N__12855\ : std_logic;
signal \N__12852\ : std_logic;
signal \N__12849\ : std_logic;
signal \N__12846\ : std_logic;
signal \N__12843\ : std_logic;
signal \N__12840\ : std_logic;
signal \N__12837\ : std_logic;
signal \N__12834\ : std_logic;
signal \N__12831\ : std_logic;
signal \N__12828\ : std_logic;
signal \N__12825\ : std_logic;
signal \N__12822\ : std_logic;
signal \N__12819\ : std_logic;
signal \N__12816\ : std_logic;
signal \N__12813\ : std_logic;
signal \N__12810\ : std_logic;
signal \N__12805\ : std_logic;
signal \N__12802\ : std_logic;
signal \N__12801\ : std_logic;
signal \N__12798\ : std_logic;
signal \N__12795\ : std_logic;
signal \N__12792\ : std_logic;
signal \N__12789\ : std_logic;
signal \N__12786\ : std_logic;
signal \N__12781\ : std_logic;
signal \N__12778\ : std_logic;
signal \N__12777\ : std_logic;
signal \N__12774\ : std_logic;
signal \N__12771\ : std_logic;
signal \N__12768\ : std_logic;
signal \N__12763\ : std_logic;
signal \N__12762\ : std_logic;
signal \N__12759\ : std_logic;
signal \N__12756\ : std_logic;
signal \N__12753\ : std_logic;
signal \N__12750\ : std_logic;
signal \N__12747\ : std_logic;
signal \N__12744\ : std_logic;
signal \N__12741\ : std_logic;
signal \N__12738\ : std_logic;
signal \N__12735\ : std_logic;
signal \N__12732\ : std_logic;
signal \N__12729\ : std_logic;
signal \N__12726\ : std_logic;
signal \N__12723\ : std_logic;
signal \N__12720\ : std_logic;
signal \N__12717\ : std_logic;
signal \N__12714\ : std_logic;
signal \N__12711\ : std_logic;
signal \N__12708\ : std_logic;
signal \N__12705\ : std_logic;
signal \N__12702\ : std_logic;
signal \N__12699\ : std_logic;
signal \N__12696\ : std_logic;
signal \N__12693\ : std_logic;
signal \N__12690\ : std_logic;
signal \N__12687\ : std_logic;
signal \N__12684\ : std_logic;
signal \N__12681\ : std_logic;
signal \N__12678\ : std_logic;
signal \N__12675\ : std_logic;
signal \N__12672\ : std_logic;
signal \N__12669\ : std_logic;
signal \N__12666\ : std_logic;
signal \N__12663\ : std_logic;
signal \N__12660\ : std_logic;
signal \N__12657\ : std_logic;
signal \N__12654\ : std_logic;
signal \N__12651\ : std_logic;
signal \N__12648\ : std_logic;
signal \N__12645\ : std_logic;
signal \N__12642\ : std_logic;
signal \N__12639\ : std_logic;
signal \N__12636\ : std_logic;
signal \N__12633\ : std_logic;
signal \N__12630\ : std_logic;
signal \N__12627\ : std_logic;
signal \N__12624\ : std_logic;
signal \N__12621\ : std_logic;
signal \N__12618\ : std_logic;
signal \N__12615\ : std_logic;
signal \N__12612\ : std_logic;
signal \N__12609\ : std_logic;
signal \N__12606\ : std_logic;
signal \N__12603\ : std_logic;
signal \N__12600\ : std_logic;
signal \N__12597\ : std_logic;
signal \N__12594\ : std_logic;
signal \N__12591\ : std_logic;
signal \N__12588\ : std_logic;
signal \N__12585\ : std_logic;
signal \N__12582\ : std_logic;
signal \N__12579\ : std_logic;
signal \N__12576\ : std_logic;
signal \N__12573\ : std_logic;
signal \N__12570\ : std_logic;
signal \N__12567\ : std_logic;
signal \N__12564\ : std_logic;
signal \N__12561\ : std_logic;
signal \N__12558\ : std_logic;
signal \N__12553\ : std_logic;
signal \N__12550\ : std_logic;
signal \N__12547\ : std_logic;
signal \N__12544\ : std_logic;
signal \N__12543\ : std_logic;
signal \N__12540\ : std_logic;
signal \N__12537\ : std_logic;
signal \N__12532\ : std_logic;
signal \N__12529\ : std_logic;
signal \N__12526\ : std_logic;
signal \N__12523\ : std_logic;
signal \N__12520\ : std_logic;
signal \N__12517\ : std_logic;
signal \N__12514\ : std_logic;
signal \N__12513\ : std_logic;
signal \N__12508\ : std_logic;
signal \N__12505\ : std_logic;
signal \N__12502\ : std_logic;
signal \N__12499\ : std_logic;
signal \N__12496\ : std_logic;
signal \N__12495\ : std_logic;
signal \N__12492\ : std_logic;
signal \N__12489\ : std_logic;
signal \N__12486\ : std_logic;
signal \N__12481\ : std_logic;
signal \N__12478\ : std_logic;
signal \N__12475\ : std_logic;
signal \N__12472\ : std_logic;
signal \N__12469\ : std_logic;
signal \N__12468\ : std_logic;
signal \N__12465\ : std_logic;
signal \N__12462\ : std_logic;
signal \N__12459\ : std_logic;
signal \N__12456\ : std_logic;
signal \N__12453\ : std_logic;
signal \N__12450\ : std_logic;
signal \N__12447\ : std_logic;
signal \N__12444\ : std_logic;
signal \N__12441\ : std_logic;
signal \N__12438\ : std_logic;
signal \N__12435\ : std_logic;
signal \N__12432\ : std_logic;
signal \N__12429\ : std_logic;
signal \N__12426\ : std_logic;
signal \N__12423\ : std_logic;
signal \N__12420\ : std_logic;
signal \N__12417\ : std_logic;
signal \N__12414\ : std_logic;
signal \N__12411\ : std_logic;
signal \N__12408\ : std_logic;
signal \N__12405\ : std_logic;
signal \N__12402\ : std_logic;
signal \N__12399\ : std_logic;
signal \N__12396\ : std_logic;
signal \N__12393\ : std_logic;
signal \N__12390\ : std_logic;
signal \N__12387\ : std_logic;
signal \N__12384\ : std_logic;
signal \N__12381\ : std_logic;
signal \N__12378\ : std_logic;
signal \N__12375\ : std_logic;
signal \N__12372\ : std_logic;
signal \N__12369\ : std_logic;
signal \N__12366\ : std_logic;
signal \N__12363\ : std_logic;
signal \N__12360\ : std_logic;
signal \N__12357\ : std_logic;
signal \N__12354\ : std_logic;
signal \N__12351\ : std_logic;
signal \N__12348\ : std_logic;
signal \N__12345\ : std_logic;
signal \N__12342\ : std_logic;
signal \N__12339\ : std_logic;
signal \N__12336\ : std_logic;
signal \N__12333\ : std_logic;
signal \N__12330\ : std_logic;
signal \N__12327\ : std_logic;
signal \N__12324\ : std_logic;
signal \N__12321\ : std_logic;
signal \N__12318\ : std_logic;
signal \N__12315\ : std_logic;
signal \N__12312\ : std_logic;
signal \N__12309\ : std_logic;
signal \N__12306\ : std_logic;
signal \N__12303\ : std_logic;
signal \N__12300\ : std_logic;
signal \N__12297\ : std_logic;
signal \N__12294\ : std_logic;
signal \N__12291\ : std_logic;
signal \N__12288\ : std_logic;
signal \N__12285\ : std_logic;
signal \N__12282\ : std_logic;
signal \N__12279\ : std_logic;
signal \N__12276\ : std_logic;
signal \N__12273\ : std_logic;
signal \N__12270\ : std_logic;
signal \N__12267\ : std_logic;
signal \N__12264\ : std_logic;
signal \N__12261\ : std_logic;
signal \N__12258\ : std_logic;
signal \N__12255\ : std_logic;
signal \N__12252\ : std_logic;
signal \N__12247\ : std_logic;
signal \N__12244\ : std_logic;
signal \N__12241\ : std_logic;
signal \N__12238\ : std_logic;
signal \N__12235\ : std_logic;
signal \N__12232\ : std_logic;
signal \N__12229\ : std_logic;
signal \N__12226\ : std_logic;
signal \N__12223\ : std_logic;
signal \N__12220\ : std_logic;
signal \N__12219\ : std_logic;
signal \N__12216\ : std_logic;
signal \N__12215\ : std_logic;
signal \N__12212\ : std_logic;
signal \N__12209\ : std_logic;
signal \N__12206\ : std_logic;
signal \N__12203\ : std_logic;
signal \N__12200\ : std_logic;
signal \N__12197\ : std_logic;
signal \N__12194\ : std_logic;
signal \N__12191\ : std_logic;
signal \N__12188\ : std_logic;
signal \N__12185\ : std_logic;
signal \N__12180\ : std_logic;
signal \N__12177\ : std_logic;
signal \N__12172\ : std_logic;
signal \N__12169\ : std_logic;
signal \N__12168\ : std_logic;
signal \N__12167\ : std_logic;
signal \N__12164\ : std_logic;
signal \N__12161\ : std_logic;
signal \N__12158\ : std_logic;
signal \N__12155\ : std_logic;
signal \N__12152\ : std_logic;
signal \N__12149\ : std_logic;
signal \N__12146\ : std_logic;
signal \N__12143\ : std_logic;
signal \N__12140\ : std_logic;
signal \N__12137\ : std_logic;
signal \N__12134\ : std_logic;
signal \N__12131\ : std_logic;
signal \N__12126\ : std_logic;
signal \N__12121\ : std_logic;
signal \N__12118\ : std_logic;
signal \N__12115\ : std_logic;
signal \N__12112\ : std_logic;
signal \N__12109\ : std_logic;
signal \N__12106\ : std_logic;
signal \N__12103\ : std_logic;
signal \N__12100\ : std_logic;
signal \N__12097\ : std_logic;
signal \N__12094\ : std_logic;
signal \N__12091\ : std_logic;
signal \N__12088\ : std_logic;
signal \N__12085\ : std_logic;
signal \N__12082\ : std_logic;
signal \N__12079\ : std_logic;
signal \N__12078\ : std_logic;
signal \N__12075\ : std_logic;
signal \N__12072\ : std_logic;
signal \N__12069\ : std_logic;
signal \N__12066\ : std_logic;
signal \N__12063\ : std_logic;
signal \N__12060\ : std_logic;
signal \N__12057\ : std_logic;
signal \N__12052\ : std_logic;
signal \N__12051\ : std_logic;
signal \N__12048\ : std_logic;
signal \N__12045\ : std_logic;
signal \N__12042\ : std_logic;
signal \N__12039\ : std_logic;
signal \N__12036\ : std_logic;
signal \N__12031\ : std_logic;
signal \N__12028\ : std_logic;
signal \N__12027\ : std_logic;
signal \N__12024\ : std_logic;
signal \N__12021\ : std_logic;
signal \N__12018\ : std_logic;
signal \N__12015\ : std_logic;
signal \N__12012\ : std_logic;
signal \N__12009\ : std_logic;
signal \N__12006\ : std_logic;
signal \N__12003\ : std_logic;
signal \N__12000\ : std_logic;
signal \N__11997\ : std_logic;
signal \N__11994\ : std_logic;
signal \N__11991\ : std_logic;
signal \N__11988\ : std_logic;
signal \N__11985\ : std_logic;
signal \N__11982\ : std_logic;
signal \N__11979\ : std_logic;
signal \N__11976\ : std_logic;
signal \N__11973\ : std_logic;
signal \N__11970\ : std_logic;
signal \N__11967\ : std_logic;
signal \N__11964\ : std_logic;
signal \N__11961\ : std_logic;
signal \N__11958\ : std_logic;
signal \N__11955\ : std_logic;
signal \N__11952\ : std_logic;
signal \N__11949\ : std_logic;
signal \N__11946\ : std_logic;
signal \N__11943\ : std_logic;
signal \N__11940\ : std_logic;
signal \N__11937\ : std_logic;
signal \N__11934\ : std_logic;
signal \N__11931\ : std_logic;
signal \N__11928\ : std_logic;
signal \N__11925\ : std_logic;
signal \N__11922\ : std_logic;
signal \N__11919\ : std_logic;
signal \N__11916\ : std_logic;
signal \N__11913\ : std_logic;
signal \N__11910\ : std_logic;
signal \N__11907\ : std_logic;
signal \N__11904\ : std_logic;
signal \N__11901\ : std_logic;
signal \N__11898\ : std_logic;
signal \N__11895\ : std_logic;
signal \N__11892\ : std_logic;
signal \N__11889\ : std_logic;
signal \N__11886\ : std_logic;
signal \N__11883\ : std_logic;
signal \N__11880\ : std_logic;
signal \N__11877\ : std_logic;
signal \N__11874\ : std_logic;
signal \N__11871\ : std_logic;
signal \N__11868\ : std_logic;
signal \N__11865\ : std_logic;
signal \N__11862\ : std_logic;
signal \N__11859\ : std_logic;
signal \N__11856\ : std_logic;
signal \N__11853\ : std_logic;
signal \N__11850\ : std_logic;
signal \N__11847\ : std_logic;
signal \N__11844\ : std_logic;
signal \N__11841\ : std_logic;
signal \N__11838\ : std_logic;
signal \N__11835\ : std_logic;
signal \N__11832\ : std_logic;
signal \N__11829\ : std_logic;
signal \N__11826\ : std_logic;
signal \N__11823\ : std_logic;
signal \N__11820\ : std_logic;
signal \N__11817\ : std_logic;
signal \N__11812\ : std_logic;
signal \N__11809\ : std_logic;
signal \N__11806\ : std_logic;
signal \N__11803\ : std_logic;
signal \N__11802\ : std_logic;
signal \N__11799\ : std_logic;
signal \N__11796\ : std_logic;
signal \N__11793\ : std_logic;
signal \N__11788\ : std_logic;
signal \N__11785\ : std_logic;
signal \N__11784\ : std_logic;
signal \N__11781\ : std_logic;
signal \N__11778\ : std_logic;
signal \N__11775\ : std_logic;
signal \N__11772\ : std_logic;
signal \N__11769\ : std_logic;
signal \N__11766\ : std_logic;
signal \N__11763\ : std_logic;
signal \N__11760\ : std_logic;
signal \N__11757\ : std_logic;
signal \N__11754\ : std_logic;
signal \N__11751\ : std_logic;
signal \N__11748\ : std_logic;
signal \N__11745\ : std_logic;
signal \N__11742\ : std_logic;
signal \N__11739\ : std_logic;
signal \N__11736\ : std_logic;
signal \N__11733\ : std_logic;
signal \N__11730\ : std_logic;
signal \N__11727\ : std_logic;
signal \N__11724\ : std_logic;
signal \N__11721\ : std_logic;
signal \N__11718\ : std_logic;
signal \N__11715\ : std_logic;
signal \N__11712\ : std_logic;
signal \N__11709\ : std_logic;
signal \N__11706\ : std_logic;
signal \N__11703\ : std_logic;
signal \N__11700\ : std_logic;
signal \N__11697\ : std_logic;
signal \N__11694\ : std_logic;
signal \N__11691\ : std_logic;
signal \N__11688\ : std_logic;
signal \N__11685\ : std_logic;
signal \N__11682\ : std_logic;
signal \N__11679\ : std_logic;
signal \N__11676\ : std_logic;
signal \N__11673\ : std_logic;
signal \N__11670\ : std_logic;
signal \N__11667\ : std_logic;
signal \N__11664\ : std_logic;
signal \N__11661\ : std_logic;
signal \N__11658\ : std_logic;
signal \N__11655\ : std_logic;
signal \N__11652\ : std_logic;
signal \N__11649\ : std_logic;
signal \N__11646\ : std_logic;
signal \N__11643\ : std_logic;
signal \N__11640\ : std_logic;
signal \N__11637\ : std_logic;
signal \N__11634\ : std_logic;
signal \N__11631\ : std_logic;
signal \N__11628\ : std_logic;
signal \N__11625\ : std_logic;
signal \N__11622\ : std_logic;
signal \N__11619\ : std_logic;
signal \N__11616\ : std_logic;
signal \N__11613\ : std_logic;
signal \N__11610\ : std_logic;
signal \N__11607\ : std_logic;
signal \N__11604\ : std_logic;
signal \N__11601\ : std_logic;
signal \N__11598\ : std_logic;
signal \N__11595\ : std_logic;
signal \N__11592\ : std_logic;
signal \N__11589\ : std_logic;
signal \N__11586\ : std_logic;
signal \N__11583\ : std_logic;
signal \N__11580\ : std_logic;
signal \N__11577\ : std_logic;
signal \N__11574\ : std_logic;
signal \N__11571\ : std_logic;
signal \N__11568\ : std_logic;
signal \N__11565\ : std_logic;
signal \N__11562\ : std_logic;
signal \N__11557\ : std_logic;
signal \N__11554\ : std_logic;
signal \N__11551\ : std_logic;
signal \N__11548\ : std_logic;
signal \N__11545\ : std_logic;
signal \N__11542\ : std_logic;
signal \N__11539\ : std_logic;
signal \N__11536\ : std_logic;
signal \N__11533\ : std_logic;
signal \N__11530\ : std_logic;
signal \N__11527\ : std_logic;
signal \N__11524\ : std_logic;
signal \N__11521\ : std_logic;
signal \N__11518\ : std_logic;
signal \N__11515\ : std_logic;
signal \N__11512\ : std_logic;
signal \N__11509\ : std_logic;
signal \N__11506\ : std_logic;
signal \N__11503\ : std_logic;
signal \N__11500\ : std_logic;
signal \N__11497\ : std_logic;
signal \N__11494\ : std_logic;
signal \N__11491\ : std_logic;
signal \N__11488\ : std_logic;
signal \N__11485\ : std_logic;
signal \N__11482\ : std_logic;
signal \N__11479\ : std_logic;
signal \N__11476\ : std_logic;
signal \N__11473\ : std_logic;
signal \N__11470\ : std_logic;
signal \N__11467\ : std_logic;
signal \N__11464\ : std_logic;
signal \N__11461\ : std_logic;
signal \N__11458\ : std_logic;
signal \N__11455\ : std_logic;
signal \N__11452\ : std_logic;
signal \N__11449\ : std_logic;
signal \N__11446\ : std_logic;
signal \N__11443\ : std_logic;
signal \N__11440\ : std_logic;
signal \N__11437\ : std_logic;
signal \N__11434\ : std_logic;
signal \N__11431\ : std_logic;
signal \N__11428\ : std_logic;
signal \N__11425\ : std_logic;
signal \N__11422\ : std_logic;
signal \N__11419\ : std_logic;
signal \N__11416\ : std_logic;
signal \N__11415\ : std_logic;
signal \N__11414\ : std_logic;
signal \N__11411\ : std_logic;
signal \N__11408\ : std_logic;
signal \N__11405\ : std_logic;
signal \N__11398\ : std_logic;
signal \N__11395\ : std_logic;
signal \N__11392\ : std_logic;
signal \N__11391\ : std_logic;
signal \N__11388\ : std_logic;
signal \N__11385\ : std_logic;
signal \N__11380\ : std_logic;
signal \N__11379\ : std_logic;
signal \N__11378\ : std_logic;
signal \N__11377\ : std_logic;
signal \N__11374\ : std_logic;
signal \N__11369\ : std_logic;
signal \N__11366\ : std_logic;
signal \N__11361\ : std_logic;
signal \N__11356\ : std_logic;
signal \N__11353\ : std_logic;
signal \N__11352\ : std_logic;
signal \N__11349\ : std_logic;
signal \N__11348\ : std_logic;
signal \N__11345\ : std_logic;
signal \N__11344\ : std_logic;
signal \N__11341\ : std_logic;
signal \N__11338\ : std_logic;
signal \N__11333\ : std_logic;
signal \N__11326\ : std_logic;
signal \N__11323\ : std_logic;
signal \N__11320\ : std_logic;
signal \N__11317\ : std_logic;
signal \N__11314\ : std_logic;
signal \N__11311\ : std_logic;
signal \N__11308\ : std_logic;
signal \N__11305\ : std_logic;
signal \N__11302\ : std_logic;
signal \N__11299\ : std_logic;
signal \N__11296\ : std_logic;
signal \N__11295\ : std_logic;
signal \N__11292\ : std_logic;
signal \N__11289\ : std_logic;
signal \N__11284\ : std_logic;
signal \N__11283\ : std_logic;
signal \N__11282\ : std_logic;
signal \N__11281\ : std_logic;
signal \N__11278\ : std_logic;
signal \N__11271\ : std_logic;
signal \N__11266\ : std_logic;
signal \N__11265\ : std_logic;
signal \N__11264\ : std_logic;
signal \N__11263\ : std_logic;
signal \N__11260\ : std_logic;
signal \N__11253\ : std_logic;
signal \N__11248\ : std_logic;
signal \N__11247\ : std_logic;
signal \N__11246\ : std_logic;
signal \N__11245\ : std_logic;
signal \N__11242\ : std_logic;
signal \N__11239\ : std_logic;
signal \N__11232\ : std_logic;
signal \N__11227\ : std_logic;
signal \N__11226\ : std_logic;
signal \N__11225\ : std_logic;
signal \N__11222\ : std_logic;
signal \N__11217\ : std_logic;
signal \N__11212\ : std_logic;
signal \N__11211\ : std_logic;
signal \N__11210\ : std_logic;
signal \N__11207\ : std_logic;
signal \N__11204\ : std_logic;
signal \N__11201\ : std_logic;
signal \N__11194\ : std_logic;
signal \N__11191\ : std_logic;
signal \N__11188\ : std_logic;
signal \N__11185\ : std_logic;
signal \N__11182\ : std_logic;
signal \N__11179\ : std_logic;
signal \N__11178\ : std_logic;
signal \N__11177\ : std_logic;
signal \N__11176\ : std_logic;
signal \N__11173\ : std_logic;
signal \N__11170\ : std_logic;
signal \N__11165\ : std_logic;
signal \N__11158\ : std_logic;
signal \N__11155\ : std_logic;
signal \N__11152\ : std_logic;
signal \N__11149\ : std_logic;
signal \N__11146\ : std_logic;
signal \N__11143\ : std_logic;
signal \N__11140\ : std_logic;
signal \N__11137\ : std_logic;
signal \N__11134\ : std_logic;
signal \N__11131\ : std_logic;
signal \N__11128\ : std_logic;
signal \N__11127\ : std_logic;
signal \N__11124\ : std_logic;
signal \N__11123\ : std_logic;
signal \N__11122\ : std_logic;
signal \N__11119\ : std_logic;
signal \N__11116\ : std_logic;
signal \N__11113\ : std_logic;
signal \N__11110\ : std_logic;
signal \N__11107\ : std_logic;
signal \N__11106\ : std_logic;
signal \N__11103\ : std_logic;
signal \N__11100\ : std_logic;
signal \N__11097\ : std_logic;
signal \N__11094\ : std_logic;
signal \N__11091\ : std_logic;
signal \N__11086\ : std_logic;
signal \N__11079\ : std_logic;
signal \N__11074\ : std_logic;
signal \N__11073\ : std_logic;
signal \N__11070\ : std_logic;
signal \N__11069\ : std_logic;
signal \N__11066\ : std_logic;
signal \N__11065\ : std_logic;
signal \N__11064\ : std_logic;
signal \N__11061\ : std_logic;
signal \N__11058\ : std_logic;
signal \N__11055\ : std_logic;
signal \N__11052\ : std_logic;
signal \N__11049\ : std_logic;
signal \N__11044\ : std_logic;
signal \N__11041\ : std_logic;
signal \N__11038\ : std_logic;
signal \N__11035\ : std_logic;
signal \N__11032\ : std_logic;
signal \N__11027\ : std_logic;
signal \N__11024\ : std_logic;
signal \N__11017\ : std_logic;
signal \N__11016\ : std_logic;
signal \N__11013\ : std_logic;
signal \N__11012\ : std_logic;
signal \N__11011\ : std_logic;
signal \N__11008\ : std_logic;
signal \N__11005\ : std_logic;
signal \N__11000\ : std_logic;
signal \N__10993\ : std_logic;
signal \N__10992\ : std_logic;
signal \N__10989\ : std_logic;
signal \N__10988\ : std_logic;
signal \N__10985\ : std_logic;
signal \N__10982\ : std_logic;
signal \N__10981\ : std_logic;
signal \N__10978\ : std_logic;
signal \N__10973\ : std_logic;
signal \N__10970\ : std_logic;
signal \N__10963\ : std_logic;
signal \N__10960\ : std_logic;
signal \N__10957\ : std_logic;
signal \N__10954\ : std_logic;
signal \N__10951\ : std_logic;
signal \N__10948\ : std_logic;
signal \N__10945\ : std_logic;
signal \N__10942\ : std_logic;
signal \N__10939\ : std_logic;
signal \N__10936\ : std_logic;
signal \N__10933\ : std_logic;
signal \N__10930\ : std_logic;
signal \N__10927\ : std_logic;
signal \N__10924\ : std_logic;
signal \N__10921\ : std_logic;
signal \N__10918\ : std_logic;
signal \N__10915\ : std_logic;
signal \N__10912\ : std_logic;
signal \N__10909\ : std_logic;
signal \N__10906\ : std_logic;
signal \N__10903\ : std_logic;
signal \N__10900\ : std_logic;
signal \N__10897\ : std_logic;
signal \N__10894\ : std_logic;
signal \N__10891\ : std_logic;
signal \N__10888\ : std_logic;
signal \N__10885\ : std_logic;
signal \N__10882\ : std_logic;
signal \N__10879\ : std_logic;
signal \N__10876\ : std_logic;
signal \N__10873\ : std_logic;
signal \N__10870\ : std_logic;
signal \N__10867\ : std_logic;
signal \N__10864\ : std_logic;
signal \N__10861\ : std_logic;
signal \N__10858\ : std_logic;
signal \N__10855\ : std_logic;
signal \N__10852\ : std_logic;
signal \N__10849\ : std_logic;
signal \N__10846\ : std_logic;
signal \N__10843\ : std_logic;
signal \N__10840\ : std_logic;
signal \N__10837\ : std_logic;
signal \N__10834\ : std_logic;
signal \N__10831\ : std_logic;
signal \N__10828\ : std_logic;
signal \N__10827\ : std_logic;
signal \N__10824\ : std_logic;
signal \N__10821\ : std_logic;
signal \N__10818\ : std_logic;
signal \N__10815\ : std_logic;
signal \N__10812\ : std_logic;
signal \N__10809\ : std_logic;
signal \N__10806\ : std_logic;
signal \N__10803\ : std_logic;
signal \N__10800\ : std_logic;
signal \N__10797\ : std_logic;
signal \N__10794\ : std_logic;
signal \N__10791\ : std_logic;
signal \N__10788\ : std_logic;
signal \N__10785\ : std_logic;
signal \N__10782\ : std_logic;
signal \N__10779\ : std_logic;
signal \N__10776\ : std_logic;
signal \N__10773\ : std_logic;
signal \N__10770\ : std_logic;
signal \N__10767\ : std_logic;
signal \N__10764\ : std_logic;
signal \N__10761\ : std_logic;
signal \N__10758\ : std_logic;
signal \N__10755\ : std_logic;
signal \N__10752\ : std_logic;
signal \N__10749\ : std_logic;
signal \N__10746\ : std_logic;
signal \N__10743\ : std_logic;
signal \N__10740\ : std_logic;
signal \N__10737\ : std_logic;
signal \N__10734\ : std_logic;
signal \N__10731\ : std_logic;
signal \N__10728\ : std_logic;
signal \N__10725\ : std_logic;
signal \N__10722\ : std_logic;
signal \N__10719\ : std_logic;
signal \N__10716\ : std_logic;
signal \N__10713\ : std_logic;
signal \N__10710\ : std_logic;
signal \N__10707\ : std_logic;
signal \N__10704\ : std_logic;
signal \N__10701\ : std_logic;
signal \N__10698\ : std_logic;
signal \N__10695\ : std_logic;
signal \N__10692\ : std_logic;
signal \N__10689\ : std_logic;
signal \N__10686\ : std_logic;
signal \N__10683\ : std_logic;
signal \N__10680\ : std_logic;
signal \N__10677\ : std_logic;
signal \N__10674\ : std_logic;
signal \N__10671\ : std_logic;
signal \N__10668\ : std_logic;
signal \N__10665\ : std_logic;
signal \N__10662\ : std_logic;
signal \N__10659\ : std_logic;
signal \N__10656\ : std_logic;
signal \N__10653\ : std_logic;
signal \N__10650\ : std_logic;
signal \N__10647\ : std_logic;
signal \N__10644\ : std_logic;
signal \N__10641\ : std_logic;
signal \N__10638\ : std_logic;
signal \N__10635\ : std_logic;
signal \N__10632\ : std_logic;
signal \N__10629\ : std_logic;
signal \N__10626\ : std_logic;
signal \N__10623\ : std_logic;
signal \N__10618\ : std_logic;
signal \N__10615\ : std_logic;
signal \N__10614\ : std_logic;
signal \N__10613\ : std_logic;
signal \N__10610\ : std_logic;
signal \N__10609\ : std_logic;
signal \N__10604\ : std_logic;
signal \N__10599\ : std_logic;
signal \N__10594\ : std_logic;
signal \N__10591\ : std_logic;
signal \N__10590\ : std_logic;
signal \N__10585\ : std_logic;
signal \N__10584\ : std_logic;
signal \N__10583\ : std_logic;
signal \N__10580\ : std_logic;
signal \N__10575\ : std_logic;
signal \N__10570\ : std_logic;
signal \N__10567\ : std_logic;
signal \N__10564\ : std_logic;
signal \N__10561\ : std_logic;
signal \N__10558\ : std_logic;
signal \N__10557\ : std_logic;
signal \N__10556\ : std_logic;
signal \N__10553\ : std_logic;
signal \N__10548\ : std_logic;
signal \N__10547\ : std_logic;
signal \N__10546\ : std_logic;
signal \N__10545\ : std_logic;
signal \N__10542\ : std_logic;
signal \N__10539\ : std_logic;
signal \N__10532\ : std_logic;
signal \N__10525\ : std_logic;
signal \N__10522\ : std_logic;
signal \N__10521\ : std_logic;
signal \N__10518\ : std_logic;
signal \N__10515\ : std_logic;
signal \N__10510\ : std_logic;
signal \N__10507\ : std_logic;
signal \N__10504\ : std_logic;
signal \N__10501\ : std_logic;
signal \N__10498\ : std_logic;
signal \N__10495\ : std_logic;
signal \N__10492\ : std_logic;
signal \N__10491\ : std_logic;
signal \N__10490\ : std_logic;
signal \N__10489\ : std_logic;
signal \N__10486\ : std_logic;
signal \N__10485\ : std_logic;
signal \N__10480\ : std_logic;
signal \N__10477\ : std_logic;
signal \N__10474\ : std_logic;
signal \N__10471\ : std_logic;
signal \N__10468\ : std_logic;
signal \N__10459\ : std_logic;
signal \N__10456\ : std_logic;
signal \N__10455\ : std_logic;
signal \N__10452\ : std_logic;
signal \N__10449\ : std_logic;
signal \N__10444\ : std_logic;
signal \N__10441\ : std_logic;
signal \N__10438\ : std_logic;
signal \N__10435\ : std_logic;
signal \N__10432\ : std_logic;
signal \N__10431\ : std_logic;
signal \N__10428\ : std_logic;
signal \N__10425\ : std_logic;
signal \N__10422\ : std_logic;
signal \N__10419\ : std_logic;
signal \N__10416\ : std_logic;
signal \N__10413\ : std_logic;
signal \N__10410\ : std_logic;
signal \N__10407\ : std_logic;
signal \N__10404\ : std_logic;
signal \N__10401\ : std_logic;
signal \N__10398\ : std_logic;
signal \N__10395\ : std_logic;
signal \N__10392\ : std_logic;
signal \N__10389\ : std_logic;
signal \N__10386\ : std_logic;
signal \N__10383\ : std_logic;
signal \N__10380\ : std_logic;
signal \N__10377\ : std_logic;
signal \N__10374\ : std_logic;
signal \N__10371\ : std_logic;
signal \N__10368\ : std_logic;
signal \N__10365\ : std_logic;
signal \N__10362\ : std_logic;
signal \N__10359\ : std_logic;
signal \N__10356\ : std_logic;
signal \N__10353\ : std_logic;
signal \N__10350\ : std_logic;
signal \N__10347\ : std_logic;
signal \N__10344\ : std_logic;
signal \N__10341\ : std_logic;
signal \N__10338\ : std_logic;
signal \N__10335\ : std_logic;
signal \N__10332\ : std_logic;
signal \N__10329\ : std_logic;
signal \N__10326\ : std_logic;
signal \N__10323\ : std_logic;
signal \N__10320\ : std_logic;
signal \N__10317\ : std_logic;
signal \N__10314\ : std_logic;
signal \N__10311\ : std_logic;
signal \N__10308\ : std_logic;
signal \N__10305\ : std_logic;
signal \N__10302\ : std_logic;
signal \N__10299\ : std_logic;
signal \N__10296\ : std_logic;
signal \N__10293\ : std_logic;
signal \N__10290\ : std_logic;
signal \N__10287\ : std_logic;
signal \N__10284\ : std_logic;
signal \N__10281\ : std_logic;
signal \N__10278\ : std_logic;
signal \N__10275\ : std_logic;
signal \N__10272\ : std_logic;
signal \N__10269\ : std_logic;
signal \N__10266\ : std_logic;
signal \N__10263\ : std_logic;
signal \N__10260\ : std_logic;
signal \N__10257\ : std_logic;
signal \N__10254\ : std_logic;
signal \N__10251\ : std_logic;
signal \N__10248\ : std_logic;
signal \N__10245\ : std_logic;
signal \N__10242\ : std_logic;
signal \N__10239\ : std_logic;
signal \N__10236\ : std_logic;
signal \N__10233\ : std_logic;
signal \N__10230\ : std_logic;
signal \N__10227\ : std_logic;
signal \N__10224\ : std_logic;
signal \N__10221\ : std_logic;
signal \N__10216\ : std_logic;
signal \N__10213\ : std_logic;
signal \N__10210\ : std_logic;
signal \N__10207\ : std_logic;
signal \N__10204\ : std_logic;
signal \N__10201\ : std_logic;
signal \N__10198\ : std_logic;
signal \N__10195\ : std_logic;
signal \N__10192\ : std_logic;
signal \N__10189\ : std_logic;
signal \N__10188\ : std_logic;
signal \N__10183\ : std_logic;
signal \N__10180\ : std_logic;
signal \N__10179\ : std_logic;
signal \N__10178\ : std_logic;
signal \N__10177\ : std_logic;
signal \N__10172\ : std_logic;
signal \N__10169\ : std_logic;
signal \N__10166\ : std_logic;
signal \N__10163\ : std_logic;
signal \N__10156\ : std_logic;
signal \N__10155\ : std_logic;
signal \N__10154\ : std_logic;
signal \N__10153\ : std_logic;
signal \N__10150\ : std_logic;
signal \N__10147\ : std_logic;
signal \N__10142\ : std_logic;
signal \N__10135\ : std_logic;
signal \N__10134\ : std_logic;
signal \N__10133\ : std_logic;
signal \N__10130\ : std_logic;
signal \N__10125\ : std_logic;
signal \N__10120\ : std_logic;
signal \N__10119\ : std_logic;
signal \N__10118\ : std_logic;
signal \N__10117\ : std_logic;
signal \N__10114\ : std_logic;
signal \N__10111\ : std_logic;
signal \N__10106\ : std_logic;
signal \N__10099\ : std_logic;
signal \N__10096\ : std_logic;
signal \N__10095\ : std_logic;
signal \N__10094\ : std_logic;
signal \N__10093\ : std_logic;
signal \N__10090\ : std_logic;
signal \N__10087\ : std_logic;
signal \N__10082\ : std_logic;
signal \N__10075\ : std_logic;
signal \N__10074\ : std_logic;
signal \N__10073\ : std_logic;
signal \N__10072\ : std_logic;
signal \N__10069\ : std_logic;
signal \N__10066\ : std_logic;
signal \N__10061\ : std_logic;
signal \N__10054\ : std_logic;
signal \N__10053\ : std_logic;
signal \N__10052\ : std_logic;
signal \N__10051\ : std_logic;
signal \N__10050\ : std_logic;
signal \N__10049\ : std_logic;
signal \N__10046\ : std_logic;
signal \N__10043\ : std_logic;
signal \N__10040\ : std_logic;
signal \N__10039\ : std_logic;
signal \N__10036\ : std_logic;
signal \N__10035\ : std_logic;
signal \N__10032\ : std_logic;
signal \N__10029\ : std_logic;
signal \N__10028\ : std_logic;
signal \N__10025\ : std_logic;
signal \N__10024\ : std_logic;
signal \N__10021\ : std_logic;
signal \N__10018\ : std_logic;
signal \N__10015\ : std_logic;
signal \N__10012\ : std_logic;
signal \N__10009\ : std_logic;
signal \N__10006\ : std_logic;
signal \N__10003\ : std_logic;
signal \N__10000\ : std_logic;
signal \N__9997\ : std_logic;
signal \N__9994\ : std_logic;
signal \N__9989\ : std_logic;
signal \N__9986\ : std_logic;
signal \N__9981\ : std_logic;
signal \N__9976\ : std_logic;
signal \N__9973\ : std_logic;
signal \N__9968\ : std_logic;
signal \N__9965\ : std_logic;
signal \N__9962\ : std_logic;
signal \N__9959\ : std_logic;
signal \N__9954\ : std_logic;
signal \N__9951\ : std_logic;
signal \N__9940\ : std_logic;
signal \N__9937\ : std_logic;
signal \N__9934\ : std_logic;
signal \N__9931\ : std_logic;
signal \N__9928\ : std_logic;
signal \N__9925\ : std_logic;
signal \N__9922\ : std_logic;
signal \N__9919\ : std_logic;
signal \N__9916\ : std_logic;
signal \N__9913\ : std_logic;
signal \N__9910\ : std_logic;
signal \N__9907\ : std_logic;
signal \N__9904\ : std_logic;
signal \N__9901\ : std_logic;
signal \N__9898\ : std_logic;
signal \N__9895\ : std_logic;
signal \N__9892\ : std_logic;
signal \N__9889\ : std_logic;
signal \N__9886\ : std_logic;
signal \N__9883\ : std_logic;
signal \N__9880\ : std_logic;
signal \N__9877\ : std_logic;
signal \N__9874\ : std_logic;
signal \N__9871\ : std_logic;
signal \N__9868\ : std_logic;
signal \N__9865\ : std_logic;
signal \N__9862\ : std_logic;
signal \N__9859\ : std_logic;
signal \N__9856\ : std_logic;
signal \N__9853\ : std_logic;
signal \N__9850\ : std_logic;
signal \N__9849\ : std_logic;
signal \N__9846\ : std_logic;
signal \N__9843\ : std_logic;
signal \N__9838\ : std_logic;
signal \N__9835\ : std_logic;
signal \N__9832\ : std_logic;
signal \N__9829\ : std_logic;
signal \N__9826\ : std_logic;
signal \N__9823\ : std_logic;
signal \N__9820\ : std_logic;
signal \N__9817\ : std_logic;
signal \N__9814\ : std_logic;
signal \N__9811\ : std_logic;
signal \N__9808\ : std_logic;
signal \N__9805\ : std_logic;
signal \N__9802\ : std_logic;
signal \N__9799\ : std_logic;
signal \N__9796\ : std_logic;
signal \N__9793\ : std_logic;
signal \N__9790\ : std_logic;
signal \N__9787\ : std_logic;
signal \N__9786\ : std_logic;
signal \N__9783\ : std_logic;
signal \N__9782\ : std_logic;
signal \N__9779\ : std_logic;
signal \N__9778\ : std_logic;
signal \N__9775\ : std_logic;
signal \N__9772\ : std_logic;
signal \N__9769\ : std_logic;
signal \N__9766\ : std_logic;
signal \N__9759\ : std_logic;
signal \N__9754\ : std_logic;
signal \N__9751\ : std_logic;
signal \N__9748\ : std_logic;
signal \N__9745\ : std_logic;
signal \N__9742\ : std_logic;
signal \N__9739\ : std_logic;
signal \N__9736\ : std_logic;
signal \N__9733\ : std_logic;
signal \N__9730\ : std_logic;
signal \N__9727\ : std_logic;
signal \N__9724\ : std_logic;
signal \N__9721\ : std_logic;
signal \N__9718\ : std_logic;
signal \N__9715\ : std_logic;
signal \N__9712\ : std_logic;
signal \N__9709\ : std_logic;
signal \N__9706\ : std_logic;
signal \N__9703\ : std_logic;
signal \N__9700\ : std_logic;
signal \N__9697\ : std_logic;
signal \N__9694\ : std_logic;
signal \N__9691\ : std_logic;
signal \N__9690\ : std_logic;
signal \N__9689\ : std_logic;
signal \N__9688\ : std_logic;
signal \N__9683\ : std_logic;
signal \N__9680\ : std_logic;
signal \N__9677\ : std_logic;
signal \N__9674\ : std_logic;
signal \N__9667\ : std_logic;
signal \N__9664\ : std_logic;
signal \N__9663\ : std_logic;
signal \N__9662\ : std_logic;
signal \N__9661\ : std_logic;
signal \N__9658\ : std_logic;
signal \N__9655\ : std_logic;
signal \N__9652\ : std_logic;
signal \N__9649\ : std_logic;
signal \N__9640\ : std_logic;
signal \N__9639\ : std_logic;
signal \N__9636\ : std_logic;
signal \N__9635\ : std_logic;
signal \N__9630\ : std_logic;
signal \N__9629\ : std_logic;
signal \N__9626\ : std_logic;
signal \N__9623\ : std_logic;
signal \N__9620\ : std_logic;
signal \N__9613\ : std_logic;
signal \N__9612\ : std_logic;
signal \N__9607\ : std_logic;
signal \N__9606\ : std_logic;
signal \N__9603\ : std_logic;
signal \N__9602\ : std_logic;
signal \N__9599\ : std_logic;
signal \N__9596\ : std_logic;
signal \N__9593\ : std_logic;
signal \N__9586\ : std_logic;
signal \N__9583\ : std_logic;
signal \N__9580\ : std_logic;
signal \N__9577\ : std_logic;
signal \N__9576\ : std_logic;
signal \N__9575\ : std_logic;
signal \N__9574\ : std_logic;
signal \N__9569\ : std_logic;
signal \N__9566\ : std_logic;
signal \N__9563\ : std_logic;
signal \N__9556\ : std_logic;
signal \N__9553\ : std_logic;
signal \N__9552\ : std_logic;
signal \N__9551\ : std_logic;
signal \N__9550\ : std_logic;
signal \N__9545\ : std_logic;
signal \N__9542\ : std_logic;
signal \N__9539\ : std_logic;
signal \N__9532\ : std_logic;
signal \N__9529\ : std_logic;
signal \N__9526\ : std_logic;
signal \N__9523\ : std_logic;
signal \N__9520\ : std_logic;
signal \N__9517\ : std_logic;
signal \N__9514\ : std_logic;
signal \N__9511\ : std_logic;
signal \N__9508\ : std_logic;
signal \N__9505\ : std_logic;
signal \N__9502\ : std_logic;
signal \N__9499\ : std_logic;
signal \N__9496\ : std_logic;
signal \N__9493\ : std_logic;
signal \N__9490\ : std_logic;
signal \N__9487\ : std_logic;
signal \N__9484\ : std_logic;
signal \N__9481\ : std_logic;
signal \N__9478\ : std_logic;
signal \N__9475\ : std_logic;
signal \N__9472\ : std_logic;
signal \N__9469\ : std_logic;
signal \N__9466\ : std_logic;
signal \N__9463\ : std_logic;
signal \N__9460\ : std_logic;
signal \N__9457\ : std_logic;
signal \N__9454\ : std_logic;
signal \N__9451\ : std_logic;
signal \N__9448\ : std_logic;
signal \N__9445\ : std_logic;
signal \N__9442\ : std_logic;
signal \N__9439\ : std_logic;
signal \N__9436\ : std_logic;
signal \N__9433\ : std_logic;
signal \N__9432\ : std_logic;
signal \N__9427\ : std_logic;
signal \N__9424\ : std_logic;
signal \N__9421\ : std_logic;
signal \N__9420\ : std_logic;
signal \N__9419\ : std_logic;
signal \N__9416\ : std_logic;
signal \N__9415\ : std_logic;
signal \N__9412\ : std_logic;
signal \N__9409\ : std_logic;
signal \N__9406\ : std_logic;
signal \N__9403\ : std_logic;
signal \N__9394\ : std_logic;
signal \N__9393\ : std_logic;
signal \N__9392\ : std_logic;
signal \N__9391\ : std_logic;
signal \N__9388\ : std_logic;
signal \N__9385\ : std_logic;
signal \N__9382\ : std_logic;
signal \N__9379\ : std_logic;
signal \N__9370\ : std_logic;
signal \N__9367\ : std_logic;
signal \N__9364\ : std_logic;
signal \N__9361\ : std_logic;
signal \N__9358\ : std_logic;
signal \N__9355\ : std_logic;
signal \N__9352\ : std_logic;
signal \N__9349\ : std_logic;
signal \N__9346\ : std_logic;
signal \N__9343\ : std_logic;
signal \N__9340\ : std_logic;
signal \N__9337\ : std_logic;
signal \N__9334\ : std_logic;
signal \N__9331\ : std_logic;
signal \N__9328\ : std_logic;
signal \N__9325\ : std_logic;
signal \N__9322\ : std_logic;
signal \N__9319\ : std_logic;
signal \N__9316\ : std_logic;
signal \N__9313\ : std_logic;
signal \N__9310\ : std_logic;
signal \N__9307\ : std_logic;
signal \N__9304\ : std_logic;
signal \N__9301\ : std_logic;
signal \N__9298\ : std_logic;
signal \N__9295\ : std_logic;
signal \N__9292\ : std_logic;
signal \N__9289\ : std_logic;
signal \N__9286\ : std_logic;
signal \N__9283\ : std_logic;
signal \N__9280\ : std_logic;
signal \N__9277\ : std_logic;
signal \N__9274\ : std_logic;
signal \N__9271\ : std_logic;
signal \N__9268\ : std_logic;
signal \N__9265\ : std_logic;
signal \N__9262\ : std_logic;
signal \N__9259\ : std_logic;
signal \N__9256\ : std_logic;
signal \N__9253\ : std_logic;
signal \N__9250\ : std_logic;
signal \N__9247\ : std_logic;
signal \N__9244\ : std_logic;
signal \N__9241\ : std_logic;
signal \N__9238\ : std_logic;
signal \N__9235\ : std_logic;
signal \N__9232\ : std_logic;
signal \N__9229\ : std_logic;
signal \N__9226\ : std_logic;
signal \N__9223\ : std_logic;
signal \N__9220\ : std_logic;
signal \N__9217\ : std_logic;
signal \N__9214\ : std_logic;
signal \N__9211\ : std_logic;
signal \N__9208\ : std_logic;
signal \N__9207\ : std_logic;
signal \N__9206\ : std_logic;
signal \N__9203\ : std_logic;
signal \N__9198\ : std_logic;
signal \N__9193\ : std_logic;
signal \N__9190\ : std_logic;
signal \N__9189\ : std_logic;
signal \N__9188\ : std_logic;
signal \N__9187\ : std_logic;
signal \N__9184\ : std_logic;
signal \N__9181\ : std_logic;
signal \N__9174\ : std_logic;
signal \N__9169\ : std_logic;
signal \N__9166\ : std_logic;
signal \N__9165\ : std_logic;
signal \N__9164\ : std_logic;
signal \N__9163\ : std_logic;
signal \N__9160\ : std_logic;
signal \N__9153\ : std_logic;
signal \N__9148\ : std_logic;
signal \N__9145\ : std_logic;
signal \N__9142\ : std_logic;
signal \N__9139\ : std_logic;
signal \N__9136\ : std_logic;
signal \N__9133\ : std_logic;
signal \N__9130\ : std_logic;
signal \N__9127\ : std_logic;
signal \N__9124\ : std_logic;
signal \N__9121\ : std_logic;
signal \N__9118\ : std_logic;
signal \N__9115\ : std_logic;
signal \N__9112\ : std_logic;
signal \N__9109\ : std_logic;
signal \N__9106\ : std_logic;
signal \N__9103\ : std_logic;
signal \N__9100\ : std_logic;
signal \N__9097\ : std_logic;
signal \N__9094\ : std_logic;
signal \N__9091\ : std_logic;
signal \N__9088\ : std_logic;
signal \N__9085\ : std_logic;
signal \N__9082\ : std_logic;
signal \N__9079\ : std_logic;
signal \N__9076\ : std_logic;
signal \N__9073\ : std_logic;
signal \N__9070\ : std_logic;
signal \N__9067\ : std_logic;
signal \N__9064\ : std_logic;
signal \N__9061\ : std_logic;
signal \N__9058\ : std_logic;
signal \N__9055\ : std_logic;
signal \N__9052\ : std_logic;
signal \N__9049\ : std_logic;
signal \N__9046\ : std_logic;
signal \N__9043\ : std_logic;
signal \N__9040\ : std_logic;
signal \N__9037\ : std_logic;
signal \N__9034\ : std_logic;
signal \N__9031\ : std_logic;
signal \N__9028\ : std_logic;
signal \N__9025\ : std_logic;
signal \N__9022\ : std_logic;
signal \N__9019\ : std_logic;
signal \N__9016\ : std_logic;
signal \N__9013\ : std_logic;
signal \N__9010\ : std_logic;
signal \N__9007\ : std_logic;
signal \N__9004\ : std_logic;
signal \N__9001\ : std_logic;
signal \N__8998\ : std_logic;
signal \N__8995\ : std_logic;
signal \N__8992\ : std_logic;
signal \N__8989\ : std_logic;
signal \N__8986\ : std_logic;
signal \N__8983\ : std_logic;
signal \N__8980\ : std_logic;
signal \N__8977\ : std_logic;
signal \N__8974\ : std_logic;
signal \N__8971\ : std_logic;
signal \N__8968\ : std_logic;
signal \N__8965\ : std_logic;
signal \N__8962\ : std_logic;
signal \N__8959\ : std_logic;
signal \N__8956\ : std_logic;
signal \N__8953\ : std_logic;
signal \N__8950\ : std_logic;
signal \N__8947\ : std_logic;
signal \N__8944\ : std_logic;
signal \N__8941\ : std_logic;
signal \N__8938\ : std_logic;
signal \N__8935\ : std_logic;
signal \N__8932\ : std_logic;
signal \N__8929\ : std_logic;
signal \N__8926\ : std_logic;
signal \N__8923\ : std_logic;
signal \N__8920\ : std_logic;
signal \N__8917\ : std_logic;
signal \N__8914\ : std_logic;
signal \N__8911\ : std_logic;
signal \N__8908\ : std_logic;
signal \N__8905\ : std_logic;
signal \N__8902\ : std_logic;
signal \N__8899\ : std_logic;
signal \N__8896\ : std_logic;
signal \N__8893\ : std_logic;
signal \N__8890\ : std_logic;
signal \N__8887\ : std_logic;
signal \N__8884\ : std_logic;
signal \N__8881\ : std_logic;
signal \N__8878\ : std_logic;
signal \N__8875\ : std_logic;
signal \N__8874\ : std_logic;
signal \N__8871\ : std_logic;
signal \N__8868\ : std_logic;
signal \N__8863\ : std_logic;
signal \N__8862\ : std_logic;
signal \N__8859\ : std_logic;
signal \N__8856\ : std_logic;
signal \N__8855\ : std_logic;
signal \N__8850\ : std_logic;
signal \N__8847\ : std_logic;
signal \N__8842\ : std_logic;
signal \N__8841\ : std_logic;
signal \N__8840\ : std_logic;
signal \N__8837\ : std_logic;
signal \N__8834\ : std_logic;
signal \N__8831\ : std_logic;
signal \N__8826\ : std_logic;
signal \N__8823\ : std_logic;
signal \N__8822\ : std_logic;
signal \N__8819\ : std_logic;
signal \N__8816\ : std_logic;
signal \N__8813\ : std_logic;
signal \N__8810\ : std_logic;
signal \N__8809\ : std_logic;
signal \N__8806\ : std_logic;
signal \N__8803\ : std_logic;
signal \N__8800\ : std_logic;
signal \N__8797\ : std_logic;
signal \N__8792\ : std_logic;
signal \N__8787\ : std_logic;
signal \N__8784\ : std_logic;
signal \N__8781\ : std_logic;
signal \N__8778\ : std_logic;
signal \N__8775\ : std_logic;
signal \N__8770\ : std_logic;
signal \N__8767\ : std_logic;
signal \N__8764\ : std_logic;
signal \N__8761\ : std_logic;
signal \N__8758\ : std_logic;
signal \N__8755\ : std_logic;
signal \N__8754\ : std_logic;
signal \N__8753\ : std_logic;
signal \N__8750\ : std_logic;
signal \N__8747\ : std_logic;
signal \N__8744\ : std_logic;
signal \N__8741\ : std_logic;
signal \N__8740\ : std_logic;
signal \N__8739\ : std_logic;
signal \N__8734\ : std_logic;
signal \N__8731\ : std_logic;
signal \N__8728\ : std_logic;
signal \N__8727\ : std_logic;
signal \N__8724\ : std_logic;
signal \N__8721\ : std_logic;
signal \N__8716\ : std_logic;
signal \N__8713\ : std_logic;
signal \N__8712\ : std_logic;
signal \N__8711\ : std_logic;
signal \N__8708\ : std_logic;
signal \N__8701\ : std_logic;
signal \N__8698\ : std_logic;
signal \N__8695\ : std_logic;
signal \N__8692\ : std_logic;
signal \N__8689\ : std_logic;
signal \N__8686\ : std_logic;
signal \N__8683\ : std_logic;
signal \N__8680\ : std_logic;
signal \N__8677\ : std_logic;
signal \N__8674\ : std_logic;
signal \N__8671\ : std_logic;
signal \N__8668\ : std_logic;
signal \N__8665\ : std_logic;
signal \N__8662\ : std_logic;
signal \N__8659\ : std_logic;
signal \N__8654\ : std_logic;
signal \N__8649\ : std_logic;
signal \N__8644\ : std_logic;
signal \N__8641\ : std_logic;
signal \N__8640\ : std_logic;
signal \N__8639\ : std_logic;
signal \N__8636\ : std_logic;
signal \N__8633\ : std_logic;
signal \N__8630\ : std_logic;
signal \N__8629\ : std_logic;
signal \N__8628\ : std_logic;
signal \N__8621\ : std_logic;
signal \N__8618\ : std_logic;
signal \N__8615\ : std_logic;
signal \N__8614\ : std_logic;
signal \N__8609\ : std_logic;
signal \N__8606\ : std_logic;
signal \N__8603\ : std_logic;
signal \N__8600\ : std_logic;
signal \N__8597\ : std_logic;
signal \N__8594\ : std_logic;
signal \N__8593\ : std_logic;
signal \N__8588\ : std_logic;
signal \N__8585\ : std_logic;
signal \N__8582\ : std_logic;
signal \N__8579\ : std_logic;
signal \N__8576\ : std_logic;
signal \N__8573\ : std_logic;
signal \N__8572\ : std_logic;
signal \N__8569\ : std_logic;
signal \N__8566\ : std_logic;
signal \N__8563\ : std_logic;
signal \N__8560\ : std_logic;
signal \N__8551\ : std_logic;
signal \N__8548\ : std_logic;
signal \N__8545\ : std_logic;
signal \N__8544\ : std_logic;
signal \N__8541\ : std_logic;
signal \N__8538\ : std_logic;
signal \N__8537\ : std_logic;
signal \N__8534\ : std_logic;
signal \N__8533\ : std_logic;
signal \N__8532\ : std_logic;
signal \N__8529\ : std_logic;
signal \N__8526\ : std_logic;
signal \N__8523\ : std_logic;
signal \N__8520\ : std_logic;
signal \N__8517\ : std_logic;
signal \N__8516\ : std_logic;
signal \N__8513\ : std_logic;
signal \N__8510\ : std_logic;
signal \N__8505\ : std_logic;
signal \N__8502\ : std_logic;
signal \N__8501\ : std_logic;
signal \N__8500\ : std_logic;
signal \N__8497\ : std_logic;
signal \N__8494\ : std_logic;
signal \N__8491\ : std_logic;
signal \N__8488\ : std_logic;
signal \N__8485\ : std_logic;
signal \N__8482\ : std_logic;
signal \N__8479\ : std_logic;
signal \N__8476\ : std_logic;
signal \N__8473\ : std_logic;
signal \N__8470\ : std_logic;
signal \N__8467\ : std_logic;
signal \N__8462\ : std_logic;
signal \N__8459\ : std_logic;
signal \N__8456\ : std_logic;
signal \N__8453\ : std_logic;
signal \N__8448\ : std_logic;
signal \N__8443\ : std_logic;
signal \N__8440\ : std_logic;
signal \N__8431\ : std_logic;
signal \N__8430\ : std_logic;
signal \N__8427\ : std_logic;
signal \N__8424\ : std_logic;
signal \N__8421\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8414\ : std_logic;
signal \N__8411\ : std_logic;
signal \N__8410\ : std_logic;
signal \N__8407\ : std_logic;
signal \N__8402\ : std_logic;
signal \N__8399\ : std_logic;
signal \N__8396\ : std_logic;
signal \N__8395\ : std_logic;
signal \N__8390\ : std_logic;
signal \N__8389\ : std_logic;
signal \N__8386\ : std_logic;
signal \N__8383\ : std_logic;
signal \N__8382\ : std_logic;
signal \N__8379\ : std_logic;
signal \N__8376\ : std_logic;
signal \N__8371\ : std_logic;
signal \N__8368\ : std_logic;
signal \N__8363\ : std_logic;
signal \N__8358\ : std_logic;
signal \N__8357\ : std_logic;
signal \N__8354\ : std_logic;
signal \N__8351\ : std_logic;
signal \N__8348\ : std_logic;
signal \N__8345\ : std_logic;
signal \N__8340\ : std_logic;
signal \N__8337\ : std_logic;
signal \N__8334\ : std_logic;
signal \N__8329\ : std_logic;
signal \N__8326\ : std_logic;
signal \N__8325\ : std_logic;
signal \N__8322\ : std_logic;
signal \N__8321\ : std_logic;
signal \N__8318\ : std_logic;
signal \N__8315\ : std_logic;
signal \N__8314\ : std_logic;
signal \N__8311\ : std_logic;
signal \N__8308\ : std_logic;
signal \N__8307\ : std_logic;
signal \N__8304\ : std_logic;
signal \N__8301\ : std_logic;
signal \N__8298\ : std_logic;
signal \N__8295\ : std_logic;
signal \N__8292\ : std_logic;
signal \N__8291\ : std_logic;
signal \N__8286\ : std_logic;
signal \N__8285\ : std_logic;
signal \N__8282\ : std_logic;
signal \N__8277\ : std_logic;
signal \N__8274\ : std_logic;
signal \N__8271\ : std_logic;
signal \N__8268\ : std_logic;
signal \N__8265\ : std_logic;
signal \N__8260\ : std_logic;
signal \N__8255\ : std_logic;
signal \N__8254\ : std_logic;
signal \N__8251\ : std_logic;
signal \N__8248\ : std_logic;
signal \N__8245\ : std_logic;
signal \N__8242\ : std_logic;
signal \N__8237\ : std_logic;
signal \N__8232\ : std_logic;
signal \N__8229\ : std_logic;
signal \N__8226\ : std_logic;
signal \N__8221\ : std_logic;
signal \N__8218\ : std_logic;
signal \N__8215\ : std_logic;
signal \N__8214\ : std_logic;
signal \N__8213\ : std_logic;
signal \N__8212\ : std_logic;
signal \N__8209\ : std_logic;
signal \N__8206\ : std_logic;
signal \N__8205\ : std_logic;
signal \N__8202\ : std_logic;
signal \N__8201\ : std_logic;
signal \N__8198\ : std_logic;
signal \N__8193\ : std_logic;
signal \N__8190\ : std_logic;
signal \N__8187\ : std_logic;
signal \N__8184\ : std_logic;
signal \N__8181\ : std_logic;
signal \N__8176\ : std_logic;
signal \N__8173\ : std_logic;
signal \N__8170\ : std_logic;
signal \N__8169\ : std_logic;
signal \N__8166\ : std_logic;
signal \N__8163\ : std_logic;
signal \N__8160\ : std_logic;
signal \N__8157\ : std_logic;
signal \N__8154\ : std_logic;
signal \N__8151\ : std_logic;
signal \N__8148\ : std_logic;
signal \N__8145\ : std_logic;
signal \N__8142\ : std_logic;
signal \N__8139\ : std_logic;
signal \N__8138\ : std_logic;
signal \N__8135\ : std_logic;
signal \N__8132\ : std_logic;
signal \N__8125\ : std_logic;
signal \N__8122\ : std_logic;
signal \N__8119\ : std_logic;
signal \N__8116\ : std_logic;
signal \N__8113\ : std_logic;
signal \N__8110\ : std_logic;
signal \N__8107\ : std_logic;
signal \N__8104\ : std_logic;
signal \N__8101\ : std_logic;
signal \N__8098\ : std_logic;
signal \N__8089\ : std_logic;
signal \N__8088\ : std_logic;
signal \N__8085\ : std_logic;
signal \N__8082\ : std_logic;
signal \N__8081\ : std_logic;
signal \N__8078\ : std_logic;
signal \N__8075\ : std_logic;
signal \N__8072\ : std_logic;
signal \N__8071\ : std_logic;
signal \N__8068\ : std_logic;
signal \N__8065\ : std_logic;
signal \N__8062\ : std_logic;
signal \N__8061\ : std_logic;
signal \N__8058\ : std_logic;
signal \N__8057\ : std_logic;
signal \N__8056\ : std_logic;
signal \N__8053\ : std_logic;
signal \N__8050\ : std_logic;
signal \N__8047\ : std_logic;
signal \N__8044\ : std_logic;
signal \N__8041\ : std_logic;
signal \N__8038\ : std_logic;
signal \N__8037\ : std_logic;
signal \N__8034\ : std_logic;
signal \N__8029\ : std_logic;
signal \N__8026\ : std_logic;
signal \N__8023\ : std_logic;
signal \N__8020\ : std_logic;
signal \N__8017\ : std_logic;
signal \N__8014\ : std_logic;
signal \N__8011\ : std_logic;
signal \N__8006\ : std_logic;
signal \N__8003\ : std_logic;
signal \N__7996\ : std_logic;
signal \N__7993\ : std_logic;
signal \N__7988\ : std_logic;
signal \N__7985\ : std_logic;
signal \N__7982\ : std_logic;
signal \TVP_VIDEO_c_3\ : std_logic;
signal \VCCG0\ : std_logic;
signal \TVP_VIDEO_c_5\ : std_logic;
signal \TVP_VIDEO_c_4\ : std_logic;
signal \TVP_VIDEO_c_7\ : std_logic;
signal \TVP_VIDEO_c_6\ : std_logic;
signal \TVP_VIDEO_c_8\ : std_logic;
signal \TVP_VIDEO_c_9\ : std_logic;
signal \TVP_VIDEO_c_2\ : std_logic;
signal \GNDG0\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_3\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_2\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_4\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_9\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_87\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_89\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_88\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_90\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_91\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_77\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_92\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_93\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_95\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_94\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_8\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_7\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_10\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_6\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_5\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_15\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_12\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_11\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_14\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_13\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_64\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_65\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_41\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_63\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_74\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_76\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_75\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_73\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_48\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_47\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_46\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_42\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_96\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_45\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_44\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_43\ : std_logic;
signal \transmit_module.video_signal_controller.n3788_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.n2876\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_0\ : std_logic;
signal \bfn_10_15_0_\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_1\ : std_logic;
signal \transmit_module.video_signal_controller.n3279\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_2\ : std_logic;
signal \transmit_module.video_signal_controller.n3280\ : std_logic;
signal \transmit_module.video_signal_controller.n3281\ : std_logic;
signal \transmit_module.video_signal_controller.n3282\ : std_logic;
signal \transmit_module.video_signal_controller.n3283\ : std_logic;
signal \transmit_module.video_signal_controller.n3284\ : std_logic;
signal \transmit_module.video_signal_controller.n3285\ : std_logic;
signal \transmit_module.video_signal_controller.n3286\ : std_logic;
signal \bfn_10_16_0_\ : std_logic;
signal \transmit_module.video_signal_controller.n3287\ : std_logic;
signal \transmit_module.video_signal_controller.n3288\ : std_logic;
signal \transmit_module.video_signal_controller.n3289\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_55\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_54\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_40\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_56\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_97\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_36\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_62\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_66\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_53\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_52\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_51\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_81\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_50\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_49\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_35\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_34\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_72\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_82\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_69\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_78\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_80\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_79\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_71\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_70\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_68\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_67\ : std_logic;
signal \transmit_module.video_signal_controller.n2886\ : std_logic;
signal \transmit_module.video_signal_controller.n1983_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.n2926\ : std_logic;
signal \transmit_module.video_signal_controller.n2010_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.n1983\ : std_logic;
signal \transmit_module.video_signal_controller.n3789\ : std_logic;
signal \transmit_module.video_signal_controller.n3467\ : std_logic;
signal \transmit_module.video_signal_controller.n18_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_3\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_5\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_8\ : std_logic;
signal \transmit_module.video_signal_controller.n4_adj_617_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_6\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_9\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_10\ : std_logic;
signal \transmit_module.video_signal_controller.n4\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_7\ : std_logic;
signal \transmit_module.video_signal_controller.n3794_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_4\ : std_logic;
signal \transmit_module.video_signal_controller.n3618\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_61\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_37\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_39\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_38\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_58\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_57\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_60\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_59\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_98\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_86\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_85\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_84\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_83\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_99\ : std_logic;
signal \bfn_12_13_0_\ : std_logic;
signal \transmit_module.video_signal_controller.n3290\ : std_logic;
signal \transmit_module.video_signal_controller.n3291\ : std_logic;
signal \transmit_module.video_signal_controller.n3292\ : std_logic;
signal \transmit_module.video_signal_controller.n3293\ : std_logic;
signal \transmit_module.video_signal_controller.n3294\ : std_logic;
signal \transmit_module.video_signal_controller.n3295\ : std_logic;
signal \transmit_module.video_signal_controller.n3296\ : std_logic;
signal \transmit_module.video_signal_controller.n3297\ : std_logic;
signal \bfn_12_14_0_\ : std_logic;
signal \transmit_module.video_signal_controller.n3298\ : std_logic;
signal \transmit_module.video_signal_controller.n3299\ : std_logic;
signal \transmit_module.video_signal_controller.n3300\ : std_logic;
signal \transmit_module.video_signal_controller.n2010\ : std_logic;
signal \transmit_module.video_signal_controller.n2361\ : std_logic;
signal \transmit_module.n3787_cascade_\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_7\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_6\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_5\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_4\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_3\ : std_logic;
signal \line_buffer.n578\ : std_logic;
signal \line_buffer.n570\ : std_logic;
signal \line_buffer.n577\ : std_logic;
signal \line_buffer.n569\ : std_logic;
signal \bfn_13_10_0_\ : std_logic;
signal \receive_module.rx_counter.n3271\ : std_logic;
signal \receive_module.rx_counter.n3272\ : std_logic;
signal \receive_module.rx_counter.n3273\ : std_logic;
signal \receive_module.rx_counter.n3274\ : std_logic;
signal \receive_module.rx_counter.n3275\ : std_logic;
signal \receive_module.rx_counter.n3276\ : std_logic;
signal \receive_module.rx_counter.n3277\ : std_logic;
signal \receive_module.rx_counter.n3278\ : std_logic;
signal \bfn_13_11_0_\ : std_logic;
signal \transmit_module.video_signal_controller.n3786_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.n8\ : std_logic;
signal \transmit_module.video_signal_controller.n7_adj_615_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.n2_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.n3785\ : std_logic;
signal \transmit_module.video_signal_controller.n3577_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.n3485\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_9\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_6\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_11\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_7\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_5\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_2\ : std_logic;
signal \transmit_module.n3798\ : std_logic;
signal \transmit_module.n112_cascade_\ : std_logic;
signal n24 : std_logic;
signal \transmit_module.old_VGA_HS\ : std_logic;
signal \transmit_module.VGA_VISIBLE_Y\ : std_logic;
signal \ADV_HSYNC_c\ : std_logic;
signal \transmit_module.video_signal_controller.n3486\ : std_logic;
signal \transmit_module.video_signal_controller.n7\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_11\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_VISIBLE_N_578\ : std_logic;
signal \transmit_module.n111_cascade_\ : std_logic;
signal n23 : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_4\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_5\ : std_logic;
signal \line_buffer.n571\ : std_logic;
signal \line_buffer.n563\ : std_logic;
signal \line_buffer.n514\ : std_logic;
signal \line_buffer.n506\ : std_logic;
signal \line_buffer.n3764\ : std_logic;
signal \line_buffer.n513\ : std_logic;
signal \line_buffer.n505\ : std_logic;
signal \line_buffer.n3646_cascade_\ : std_logic;
signal \line_buffer.n3647\ : std_logic;
signal \receive_module.rx_counter.Y_3\ : std_logic;
signal \receive_module.rx_counter.Y_2\ : std_logic;
signal \receive_module.rx_counter.Y_1\ : std_logic;
signal \receive_module.rx_counter.Y_5\ : std_logic;
signal \receive_module.rx_counter.Y_6\ : std_logic;
signal \receive_module.rx_counter.n4_adj_604\ : std_logic;
signal \receive_module.rx_counter.n5_cascade_\ : std_logic;
signal \receive_module.rx_counter.n3548\ : std_logic;
signal \receive_module.rx_counter.Y_0\ : std_logic;
signal \receive_module.rx_counter.n14_adj_611\ : std_logic;
signal \receive_module.rx_counter.n10_adj_610\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_7\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_1\ : std_logic;
signal \transmit_module.n2093\ : std_logic;
signal \transmit_module.n2147\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_4\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_8\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_0\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_3\ : std_logic;
signal \transmit_module.video_signal_controller.n3626_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_1\ : std_logic;
signal \transmit_module.n111\ : std_logic;
signal \transmit_module.n143\ : std_logic;
signal \transmit_module.n143_cascade_\ : std_logic;
signal \transmit_module.n112\ : std_logic;
signal \transmit_module.n142\ : std_logic;
signal \transmit_module.n141_cascade_\ : std_logic;
signal \transmit_module.n137_cascade_\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_1\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_10\ : std_logic;
signal \transmit_module.video_signal_controller.n3632\ : std_logic;
signal \transmit_module.video_signal_controller.n18_adj_616\ : std_logic;
signal \transmit_module.video_signal_controller.n3614\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_10\ : std_logic;
signal \transmit_module.n146\ : std_logic;
signal \transmit_module.n146_cascade_\ : std_logic;
signal \transmit_module.n115\ : std_logic;
signal n27 : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_2\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_1\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_9\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_8\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_10\ : std_logic;
signal \line_buffer.n507\ : std_logic;
signal \line_buffer.n499\ : std_logic;
signal \line_buffer.n3752\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_6\ : std_logic;
signal \transmit_module.n106\ : std_logic;
signal \transmit_module.n137\ : std_logic;
signal n18 : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_0\ : std_logic;
signal \line_buffer.n3722\ : std_logic;
signal \TX_DATA_6\ : std_logic;
signal n1792 : std_logic;
signal n1798 : std_logic;
signal \line_buffer.n448\ : std_logic;
signal \line_buffer.n440\ : std_logic;
signal \line_buffer.n3679\ : std_logic;
signal \transmit_module.n116\ : std_logic;
signal \transmit_module.n147\ : std_logic;
signal n28 : std_logic;
signal \transmit_module.n110\ : std_logic;
signal \transmit_module.n141\ : std_logic;
signal n22 : std_logic;
signal \transmit_module.n109\ : std_logic;
signal \transmit_module.n140\ : std_logic;
signal n21 : std_logic;
signal \LED_c\ : std_logic;
signal \receive_module.rx_counter.n3628_cascade_\ : std_logic;
signal \receive_module.rx_counter.n7_adj_609\ : std_logic;
signal \receive_module.rx_counter.n11\ : std_logic;
signal \receive_module.rx_counter.n11_cascade_\ : std_logic;
signal \receive_module.rx_counter.old_VS\ : std_logic;
signal \line_buffer.n543\ : std_logic;
signal \line_buffer.n535\ : std_logic;
signal \receive_module.rx_counter.Y_7\ : std_logic;
signal \receive_module.rx_counter.n3791\ : std_logic;
signal \receive_module.rx_counter.Y_4\ : std_logic;
signal \receive_module.rx_counter.n3551\ : std_logic;
signal \receive_module.rx_counter.n2045\ : std_logic;
signal \receive_module.rx_counter.old_HS\ : std_logic;
signal \bfn_15_11_0_\ : std_logic;
signal \receive_module.n3245\ : std_logic;
signal \receive_module.n3246\ : std_logic;
signal \receive_module.n3247\ : std_logic;
signal \receive_module.n3248\ : std_logic;
signal \receive_module.n3249\ : std_logic;
signal \receive_module.n3250\ : std_logic;
signal \receive_module.n3251\ : std_logic;
signal \receive_module.n3252\ : std_logic;
signal \bfn_15_12_0_\ : std_logic;
signal \receive_module.n3253\ : std_logic;
signal \receive_module.n3254\ : std_logic;
signal \receive_module.n3255\ : std_logic;
signal \receive_module.n3256\ : std_logic;
signal \receive_module.n3257\ : std_logic;
signal \transmit_module.TX_ADDR_0\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_0\ : std_logic;
signal \transmit_module.n132\ : std_logic;
signal \bfn_15_13_0_\ : std_logic;
signal \transmit_module.TX_ADDR_1\ : std_logic;
signal \transmit_module.n131\ : std_logic;
signal \transmit_module.n3258\ : std_logic;
signal \transmit_module.n3259\ : std_logic;
signal \transmit_module.n3260\ : std_logic;
signal \transmit_module.TX_ADDR_4\ : std_logic;
signal \transmit_module.n128\ : std_logic;
signal \transmit_module.n3261\ : std_logic;
signal \transmit_module.TX_ADDR_5\ : std_logic;
signal \transmit_module.n127\ : std_logic;
signal \transmit_module.n3262\ : std_logic;
signal \transmit_module.TX_ADDR_6\ : std_logic;
signal \transmit_module.n126\ : std_logic;
signal \transmit_module.n3263\ : std_logic;
signal \transmit_module.TX_ADDR_7\ : std_logic;
signal \transmit_module.n125\ : std_logic;
signal \transmit_module.n3264\ : std_logic;
signal \transmit_module.n3265\ : std_logic;
signal \bfn_15_14_0_\ : std_logic;
signal \transmit_module.n3266\ : std_logic;
signal \transmit_module.TX_ADDR_10\ : std_logic;
signal \transmit_module.n122\ : std_logic;
signal \transmit_module.n3267\ : std_logic;
signal \transmit_module.n3268\ : std_logic;
signal \transmit_module.n3269\ : std_logic;
signal \transmit_module.n3270\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_9\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_12\ : std_logic;
signal \transmit_module.n120\ : std_logic;
signal \transmit_module.n119\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_11\ : std_logic;
signal \transmit_module.n121\ : std_logic;
signal \transmit_module.n2039\ : std_logic;
signal \transmit_module.n130\ : std_logic;
signal \line_buffer.n3755\ : std_logic;
signal \TX_DATA_0\ : std_logic;
signal \receive_module.n134\ : std_logic;
signal \RX_ADDR_2\ : std_logic;
signal \line_buffer.n545\ : std_logic;
signal \line_buffer.n537\ : std_logic;
signal \line_buffer.n3680\ : std_logic;
signal \receive_module.n126\ : std_logic;
signal \RX_ADDR_10\ : std_logic;
signal \receive_module.n132\ : std_logic;
signal \RX_ADDR_4\ : std_logic;
signal \receive_module.n131\ : std_logic;
signal \RX_ADDR_5\ : std_logic;
signal \receive_module.n130\ : std_logic;
signal \RX_ADDR_6\ : std_logic;
signal \receive_module.n129\ : std_logic;
signal \RX_ADDR_7\ : std_logic;
signal \receive_module.n128\ : std_logic;
signal \RX_ADDR_8\ : std_logic;
signal \receive_module.n127\ : std_logic;
signal \RX_ADDR_9\ : std_logic;
signal \receive_module.rx_counter.FRAME_COUNTER_0\ : std_logic;
signal \bfn_16_5_0_\ : std_logic;
signal \receive_module.rx_counter.FRAME_COUNTER_1\ : std_logic;
signal \receive_module.rx_counter.n3310\ : std_logic;
signal \receive_module.rx_counter.FRAME_COUNTER_2\ : std_logic;
signal \receive_module.rx_counter.n3311\ : std_logic;
signal \receive_module.rx_counter.FRAME_COUNTER_3\ : std_logic;
signal \receive_module.rx_counter.n3312\ : std_logic;
signal \receive_module.rx_counter.FRAME_COUNTER_4\ : std_logic;
signal \receive_module.rx_counter.n3313\ : std_logic;
signal \receive_module.rx_counter.n3314\ : std_logic;
signal \receive_module.rx_counter.FRAME_COUNTER_5\ : std_logic;
signal \receive_module.rx_counter.n3792\ : std_logic;
signal \receive_module.rx_counter.n2517\ : std_logic;
signal \receive_module.n136\ : std_logic;
signal \RX_ADDR_0\ : std_logic;
signal \receive_module.n135\ : std_logic;
signal \RX_ADDR_1\ : std_logic;
signal \line_buffer.n511\ : std_logic;
signal \line_buffer.n503\ : std_logic;
signal \line_buffer.n509\ : std_logic;
signal \line_buffer.n501\ : std_logic;
signal \receive_module.rx_counter.n4_cascade_\ : std_logic;
signal \receive_module.rx_counter.n6_cascade_\ : std_logic;
signal \receive_module.rx_counter.n3534\ : std_logic;
signal \receive_module.rx_counter.n3581\ : std_logic;
signal \line_buffer.n517\ : std_logic;
signal \line_buffer.n452\ : std_logic;
signal \line_buffer.n548\ : std_logic;
signal \receive_module.n3795\ : std_logic;
signal \line_buffer.n451\ : std_logic;
signal \line_buffer.n549\ : std_logic;
signal \line_buffer.n516\ : std_logic;
signal \receive_module.rx_counter.n3575\ : std_logic;
signal \receive_module.rx_counter.n4_adj_606\ : std_logic;
signal \receive_module.rx_counter.Y_8\ : std_logic;
signal \receive_module.rx_counter.n55_adj_607\ : std_logic;
signal \line_buffer.n581\ : std_logic;
signal \RX_ADDR_12\ : std_logic;
signal \RX_ADDR_13\ : std_logic;
signal \RX_ADDR_11\ : std_logic;
signal \line_buffer.n580\ : std_logic;
signal \RX_TX_SYNC_BUFF\ : std_logic;
signal \RX_TX_SYNC\ : std_logic;
signal \sync_buffer.BUFFER_0\ : std_logic;
signal \sync_buffer.BUFFER_1\ : std_logic;
signal \INVsync_buffer.WIRE_OUT_8C_net\ : std_logic;
signal \transmit_module.n124\ : std_logic;
signal \transmit_module.n139_cascade_\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_8\ : std_logic;
signal \transmit_module.TX_ADDR_8\ : std_logic;
signal \transmit_module.TX_ADDR_9\ : std_logic;
signal \transmit_module.n123\ : std_logic;
signal \transmit_module.n138\ : std_logic;
signal \transmit_module.n138_cascade_\ : std_logic;
signal \transmit_module.n107\ : std_logic;
signal n19 : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_13\ : std_logic;
signal \line_buffer.n3634\ : std_logic;
signal \line_buffer.n442\ : std_logic;
signal \line_buffer.n434\ : std_logic;
signal \line_buffer.n3749\ : std_logic;
signal \line_buffer.n541\ : std_logic;
signal \line_buffer.n533\ : std_logic;
signal \line_buffer.n3676\ : std_logic;
signal \line_buffer.n3674\ : std_logic;
signal \line_buffer.n3716\ : std_logic;
signal \line_buffer.n446\ : std_logic;
signal \line_buffer.n438\ : std_logic;
signal \line_buffer.n3728\ : std_logic;
signal \line_buffer.n3640_cascade_\ : std_logic;
signal \line_buffer.n3641\ : std_logic;
signal \transmit_module.n114\ : std_logic;
signal \transmit_module.n145\ : std_logic;
signal n26 : std_logic;
signal \transmit_module.VGA_VISIBLE\ : std_logic;
signal \transmit_module.n129\ : std_logic;
signal \transmit_module.n144\ : std_logic;
signal \transmit_module.n144_cascade_\ : std_logic;
signal n25 : std_logic;
signal \transmit_module.TX_ADDR_2\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_2\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_0\ : std_logic;
signal \transmit_module.n113\ : std_logic;
signal \transmit_module.TX_ADDR_3\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_3\ : std_logic;
signal \transmit_module.n2061\ : std_logic;
signal \TX_DATA_4\ : std_logic;
signal n1794 : std_logic;
signal \TX_DATA_2\ : std_logic;
signal n1796 : std_logic;
signal \line_buffer.n444\ : std_logic;
signal \line_buffer.n436\ : std_logic;
signal \line_buffer.n3673\ : std_logic;
signal \transmit_module.n3787\ : std_logic;
signal \transmit_module.n108\ : std_logic;
signal \transmit_module.n139\ : std_logic;
signal n20 : std_logic;
signal \GB_BUFFER_TVP_CLK_c_THRU_CO\ : std_logic;
signal \TVP_HSYNC_c\ : std_logic;
signal \receive_module.rx_counter.n10\ : std_logic;
signal \bfn_17_10_0_\ : std_logic;
signal \receive_module.rx_counter.n9\ : std_logic;
signal \receive_module.rx_counter.n3301\ : std_logic;
signal \receive_module.rx_counter.n8\ : std_logic;
signal \receive_module.rx_counter.n3302\ : std_logic;
signal \receive_module.rx_counter.X_3\ : std_logic;
signal \receive_module.rx_counter.n3303\ : std_logic;
signal \receive_module.rx_counter.X_4\ : std_logic;
signal \receive_module.rx_counter.n3304\ : std_logic;
signal \receive_module.rx_counter.X_5\ : std_logic;
signal \receive_module.rx_counter.n3305\ : std_logic;
signal \receive_module.rx_counter.X_6\ : std_logic;
signal \receive_module.rx_counter.n3306\ : std_logic;
signal \receive_module.rx_counter.X_7\ : std_logic;
signal \receive_module.rx_counter.n3307\ : std_logic;
signal \receive_module.rx_counter.n3308\ : std_logic;
signal \receive_module.rx_counter.X_8\ : std_logic;
signal \bfn_17_11_0_\ : std_logic;
signal \receive_module.rx_counter.n3309\ : std_logic;
signal \receive_module.rx_counter.X_9\ : std_logic;
signal \receive_module.rx_counter.n3790\ : std_logic;
signal \line_buffer.n576\ : std_logic;
signal \line_buffer.n568\ : std_logic;
signal \line_buffer.n504\ : std_logic;
signal \line_buffer.n512\ : std_logic;
signal \line_buffer.n3734_cascade_\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_12\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_11\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_25\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_26\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_13\ : std_logic;
signal \line_buffer.n539\ : std_logic;
signal \line_buffer.n531\ : std_logic;
signal \line_buffer.n3746\ : std_logic;
signal \line_buffer.n573\ : std_logic;
signal \line_buffer.n565\ : std_logic;
signal \line_buffer.n3677\ : std_logic;
signal \line_buffer.n567\ : std_logic;
signal \line_buffer.n575\ : std_logic;
signal \line_buffer.n3635\ : std_logic;
signal \line_buffer.n3737\ : std_logic;
signal \line_buffer.n447\ : std_logic;
signal \line_buffer.n439\ : std_logic;
signal \line_buffer.n3701\ : std_logic;
signal \TX_DATA_5\ : std_logic;
signal n1793 : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_33\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_27\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_28\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_29\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_30\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_32\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_31\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_22\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_24\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_23\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_16\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_17\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_19\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_18\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_15\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_14\ : std_logic;
signal n1797 : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_21\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_20\ : std_logic;
signal \transmit_module.n3797\ : std_logic;
signal \ADV_VSYNC_c\ : std_logic;
signal \line_buffer.n544\ : std_logic;
signal \line_buffer.n536\ : std_logic;
signal \line_buffer.n3698\ : std_logic;
signal \line_buffer.n508\ : std_logic;
signal \line_buffer.n500\ : std_logic;
signal \line_buffer.n3695_cascade_\ : std_logic;
signal \TX_DATA_1\ : std_logic;
signal \line_buffer.n572\ : std_logic;
signal \line_buffer.n564\ : std_logic;
signal \line_buffer.n3692\ : std_logic;
signal \RX_WE\ : std_logic;
signal \receive_module.n133\ : std_logic;
signal \TVP_VSYNC_c\ : std_logic;
signal \RX_ADDR_3\ : std_logic;
signal \TVP_CLK_c\ : std_logic;
signal \receive_module.n3793\ : std_logic;
signal \line_buffer.n542\ : std_logic;
signal \line_buffer.n534\ : std_logic;
signal \line_buffer.n445\ : std_logic;
signal \line_buffer.n437\ : std_logic;
signal \line_buffer.n3710\ : std_logic;
signal \line_buffer.n566\ : std_logic;
signal \line_buffer.n574\ : std_logic;
signal \line_buffer.n502\ : std_logic;
signal \line_buffer.n510\ : std_logic;
signal \line_buffer.n3758_cascade_\ : std_logic;
signal \line_buffer.n540\ : std_logic;
signal \line_buffer.n532\ : std_logic;
signal \line_buffer.n435\ : std_logic;
signal \line_buffer.n443\ : std_logic;
signal \line_buffer.n3740_cascade_\ : std_logic;
signal \line_buffer.n3743\ : std_logic;
signal \line_buffer.n3761\ : std_logic;
signal \line_buffer.n3713\ : std_logic;
signal \TX_ADDR_13\ : std_logic;
signal \line_buffer.n3767\ : std_logic;
signal \TX_ADDR_11\ : std_logic;
signal \line_buffer.n546\ : std_logic;
signal \line_buffer.n538\ : std_logic;
signal \TX_DATA_3\ : std_logic;
signal n1795 : std_logic;
signal \TX_DATA_7\ : std_logic;
signal \ADV_B_c\ : std_logic;
signal \ADV_CLK_c\ : std_logic;
signal \transmit_module.n2354\ : std_logic;
signal \line_buffer.n449\ : std_logic;
signal \TX_ADDR_12\ : std_logic;
signal \line_buffer.n441\ : std_logic;
signal \line_buffer.n3704\ : std_logic;
signal \line_buffer.n3707\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \TVP_CLK_wire\ : std_logic;
signal \ADV_CLK_wire\ : std_logic;
signal \TVP_VIDEO_wire\ : std_logic_vector(9 downto 0);
signal \ADV_G_wire\ : std_logic_vector(7 downto 0);
signal \ADV_R_wire\ : std_logic_vector(7 downto 0);
signal \ADV_B_wire\ : std_logic_vector(7 downto 0);
signal \ADV_SYNC_N_wire\ : std_logic;
signal \TVP_HSYNC_wire\ : std_logic;
signal \TVP_VSYNC_wire\ : std_logic;
signal \ADV_BLANK_N_wire\ : std_logic;
signal \LED_wire\ : std_logic;
signal \ADV_HSYNC_wire\ : std_logic;
signal \ADV_VSYNC_wire\ : std_logic;
signal \tx_pll.TX_PLL_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);
signal \line_buffer.mem2_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem2_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem2_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem2_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem2_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem14_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem14_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem14_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem14_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem14_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem5_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem5_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem5_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem5_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem5_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem11_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem11_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem11_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem11_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem11_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem21_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem21_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem21_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem21_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem21_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem12_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem12_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem12_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem12_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem12_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem18_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem18_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem18_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem18_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem18_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem24_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem24_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem24_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem24_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem24_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem15_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem15_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem15_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem15_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem15_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem27_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem27_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem27_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem27_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem27_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem4_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem4_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem4_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem4_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem4_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem16_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem16_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem16_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem16_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem16_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem30_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem30_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem30_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem30_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem30_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem7_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem7_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem7_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem7_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem7_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem20_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem20_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem20_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem20_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem20_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem13_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem13_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem13_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem13_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem13_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem19_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem19_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem19_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem19_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem19_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem23_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem23_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem23_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem23_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem23_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem26_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem26_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem26_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem26_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem26_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem3_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem3_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem3_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem3_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem3_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem17_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem17_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem17_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem17_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem17_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem31_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem31_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem31_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem31_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem31_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem9_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem9_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem9_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem9_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem9_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem29_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem29_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem29_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem29_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem29_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem6_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem6_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem6_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem6_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem6_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem10_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem10_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem10_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem10_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem10_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem22_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem22_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem22_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem22_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem22_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem25_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem25_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem25_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem25_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem25_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem8_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem8_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem8_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem8_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem8_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem28_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem28_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem28_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem28_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem28_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    \TVP_CLK_wire\ <= TVP_CLK;
    ADV_CLK <= \ADV_CLK_wire\;
    \TVP_VIDEO_wire\ <= TVP_VIDEO;
    ADV_G <= \ADV_G_wire\;
    ADV_R <= \ADV_R_wire\;
    ADV_B <= \ADV_B_wire\;
    ADV_SYNC_N <= \ADV_SYNC_N_wire\;
    \TVP_HSYNC_wire\ <= TVP_HSYNC;
    \TVP_VSYNC_wire\ <= TVP_VSYNC;
    ADV_BLANK_N <= \ADV_BLANK_N_wire\;
    LED <= \LED_wire\;
    ADV_HSYNC <= \ADV_HSYNC_wire\;
    ADV_VSYNC <= \ADV_VSYNC_wire\;
    \tx_pll.TX_PLL_inst_DYNAMICDELAY_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.n449\ <= \line_buffer.mem2_physical_RDATA_wire\(11);
    \line_buffer.n448\ <= \line_buffer.mem2_physical_RDATA_wire\(3);
    \line_buffer.mem2_physical_RADDR_wire\ <= \N__12333\&\N__17139\&\N__18750\&\N__12621\&\N__12885\&\N__10308\&\N__10683\&\N__18051\&\N__18399\&\N__11649\&\N__11892\;
    \line_buffer.mem2_physical_WADDR_wire\ <= \N__15513\&\N__13995\&\N__14256\&\N__14505\&\N__14760\&\N__15021\&\N__15258\&\N__20280\&\N__13641\&\N__15816\&\N__16071\;
    \line_buffer.mem2_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem2_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8614\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8739\&'0'&'0'&'0';
    \line_buffer.n536\ <= \line_buffer.mem14_physical_RDATA_wire\(11);
    \line_buffer.n535\ <= \line_buffer.mem14_physical_RDATA_wire\(3);
    \line_buffer.mem14_physical_RADDR_wire\ <= \N__12405\&\N__17211\&\N__18822\&\N__12693\&\N__12957\&\N__10380\&\N__10755\&\N__18123\&\N__18471\&\N__11721\&\N__11964\;
    \line_buffer.mem14_physical_WADDR_wire\ <= \N__15585\&\N__14067\&\N__14328\&\N__14577\&\N__14832\&\N__15093\&\N__15330\&\N__20352\&\N__13713\&\N__15888\&\N__16143\;
    \line_buffer.mem14_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem14_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8537\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8410\&'0'&'0'&'0';
    \line_buffer.n546\ <= \line_buffer.mem5_physical_RDATA_wire\(11);
    \line_buffer.n545\ <= \line_buffer.mem5_physical_RDATA_wire\(3);
    \line_buffer.mem5_physical_RADDR_wire\ <= \N__12336\&\N__17154\&\N__18753\&\N__12630\&\N__12882\&\N__10299\&\N__10710\&\N__18060\&\N__18402\&\N__11652\&\N__11895\;
    \line_buffer.mem5_physical_WADDR_wire\ <= \N__15534\&\N__14016\&\N__14259\&\N__14514\&\N__14763\&\N__15030\&\N__15267\&\N__20289\&\N__13650\&\N__15825\&\N__16092\;
    \line_buffer.mem5_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem5_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8639\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8753\&'0'&'0'&'0';
    \line_buffer.n504\ <= \line_buffer.mem11_physical_RDATA_wire\(11);
    \line_buffer.n503\ <= \line_buffer.mem11_physical_RDATA_wire\(3);
    \line_buffer.mem11_physical_RADDR_wire\ <= \N__12441\&\N__17247\&\N__18858\&\N__12729\&\N__12993\&\N__10416\&\N__10791\&\N__18159\&\N__18507\&\N__11757\&\N__12000\;
    \line_buffer.mem11_physical_WADDR_wire\ <= \N__15621\&\N__14103\&\N__14364\&\N__14613\&\N__14868\&\N__15129\&\N__15366\&\N__20388\&\N__13749\&\N__15924\&\N__16179\;
    \line_buffer.mem11_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem11_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8501\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8389\&'0'&'0'&'0';
    \line_buffer.n566\ <= \line_buffer.mem21_physical_RDATA_wire\(11);
    \line_buffer.n565\ <= \line_buffer.mem21_physical_RDATA_wire\(3);
    \line_buffer.mem21_physical_RADDR_wire\ <= \N__12309\&\N__17115\&\N__18726\&\N__12597\&\N__12861\&\N__10284\&\N__10659\&\N__18027\&\N__18375\&\N__11625\&\N__11868\;
    \line_buffer.mem21_physical_WADDR_wire\ <= \N__15489\&\N__13970\&\N__14232\&\N__14481\&\N__14736\&\N__14997\&\N__15234\&\N__20256\&\N__13617\&\N__15792\&\N__16047\;
    \line_buffer.mem21_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem21_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8321\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8221\&'0'&'0'&'0';
    \line_buffer.n502\ <= \line_buffer.mem12_physical_RDATA_wire\(11);
    \line_buffer.n501\ <= \line_buffer.mem12_physical_RDATA_wire\(3);
    \line_buffer.mem12_physical_RADDR_wire\ <= \N__12429\&\N__17235\&\N__18846\&\N__12717\&\N__12981\&\N__10404\&\N__10779\&\N__18147\&\N__18495\&\N__11745\&\N__11988\;
    \line_buffer.mem12_physical_WADDR_wire\ <= \N__15609\&\N__14091\&\N__14352\&\N__14601\&\N__14856\&\N__15117\&\N__15354\&\N__20376\&\N__13737\&\N__15912\&\N__16167\;
    \line_buffer.mem12_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem12_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8291\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8213\&'0'&'0'&'0';
    \line_buffer.n445\ <= \line_buffer.mem18_physical_RDATA_wire\(11);
    \line_buffer.n444\ <= \line_buffer.mem18_physical_RDATA_wire\(3);
    \line_buffer.mem18_physical_RADDR_wire\ <= \N__12357\&\N__17163\&\N__18774\&\N__12645\&\N__12909\&\N__10332\&\N__10707\&\N__18075\&\N__18423\&\N__11673\&\N__11916\;
    \line_buffer.mem18_physical_WADDR_wire\ <= \N__15537\&\N__14019\&\N__14280\&\N__14529\&\N__14784\&\N__15045\&\N__15282\&\N__20304\&\N__13665\&\N__15840\&\N__16095\;
    \line_buffer.mem18_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem18_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8325\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8214\&'0'&'0'&'0';
    \line_buffer.n510\ <= \line_buffer.mem24_physical_RDATA_wire\(11);
    \line_buffer.n509\ <= \line_buffer.mem24_physical_RDATA_wire\(3);
    \line_buffer.mem24_physical_RADDR_wire\ <= \N__12456\&\N__17274\&\N__18873\&\N__12750\&\N__13002\&\N__10419\&\N__10828\&\N__18180\&\N__18522\&\N__11772\&\N__12015\;
    \line_buffer.mem24_physical_WADDR_wire\ <= \N__15654\&\N__14136\&\N__14379\&\N__14634\&\N__14883\&\N__15150\&\N__15387\&\N__20409\&\N__13770\&\N__15945\&\N__16212\;
    \line_buffer.mem24_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem24_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8254\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8138\&'0'&'0'&'0';
    \line_buffer.n538\ <= \line_buffer.mem1_physical_RDATA_wire\(11);
    \line_buffer.n537\ <= \line_buffer.mem1_physical_RDATA_wire\(3);
    \line_buffer.mem1_physical_RADDR_wire\ <= \N__12465\&\N__17271\&\N__18882\&\N__12753\&\N__13015\&\N__10435\&\N__10815\&\N__18183\&\N__18531\&\N__11781\&\N__12024\;
    \line_buffer.mem1_physical_WADDR_wire\ <= \N__15645\&\N__14127\&\N__14388\&\N__14637\&\N__14892\&\N__15153\&\N__15390\&\N__20412\&\N__13773\&\N__15948\&\N__16203\;
    \line_buffer.mem1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8593\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8712\&'0'&'0'&'0';
    \line_buffer.n534\ <= \line_buffer.mem15_physical_RDATA_wire\(11);
    \line_buffer.n533\ <= \line_buffer.mem15_physical_RDATA_wire\(3);
    \line_buffer.mem15_physical_RADDR_wire\ <= \N__12393\&\N__17199\&\N__18810\&\N__12681\&\N__12945\&\N__10368\&\N__10743\&\N__18111\&\N__18459\&\N__11709\&\N__11952\;
    \line_buffer.mem15_physical_WADDR_wire\ <= \N__15573\&\N__14055\&\N__14316\&\N__14565\&\N__14820\&\N__15081\&\N__15318\&\N__20340\&\N__13701\&\N__15876\&\N__16131\;
    \line_buffer.mem15_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem15_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8307\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8205\&'0'&'0'&'0';
    \line_buffer.n542\ <= \line_buffer.mem27_physical_RDATA_wire\(11);
    \line_buffer.n541\ <= \line_buffer.mem27_physical_RDATA_wire\(3);
    \line_buffer.mem27_physical_RADDR_wire\ <= \N__12420\&\N__17238\&\N__18837\&\N__12714\&\N__12966\&\N__10383\&\N__10794\&\N__18144\&\N__18486\&\N__11736\&\N__11979\;
    \line_buffer.mem27_physical_WADDR_wire\ <= \N__15618\&\N__14100\&\N__14343\&\N__14598\&\N__14847\&\N__15114\&\N__15351\&\N__20373\&\N__13734\&\N__15909\&\N__16176\;
    \line_buffer.mem27_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem27_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8285\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8169\&'0'&'0'&'0';
    \line_buffer.n514\ <= \line_buffer.mem4_physical_RDATA_wire\(11);
    \line_buffer.n513\ <= \line_buffer.mem4_physical_RDATA_wire\(3);
    \line_buffer.mem4_physical_RADDR_wire\ <= \N__12348\&\N__17166\&\N__18765\&\N__12642\&\N__12894\&\N__10311\&\N__10722\&\N__18072\&\N__18414\&\N__11664\&\N__11907\;
    \line_buffer.mem4_physical_WADDR_wire\ <= \N__15546\&\N__14028\&\N__14271\&\N__14526\&\N__14775\&\N__15042\&\N__15279\&\N__20301\&\N__13662\&\N__15837\&\N__16104\;
    \line_buffer.mem4_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem4_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8629\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8740\&'0'&'0'&'0';
    \line_buffer.n532\ <= \line_buffer.mem16_physical_RDATA_wire\(11);
    \line_buffer.n531\ <= \line_buffer.mem16_physical_RDATA_wire\(3);
    \line_buffer.mem16_physical_RADDR_wire\ <= \N__12381\&\N__17187\&\N__18798\&\N__12669\&\N__12933\&\N__10356\&\N__10731\&\N__18099\&\N__18447\&\N__11697\&\N__11940\;
    \line_buffer.mem16_physical_WADDR_wire\ <= \N__15561\&\N__14043\&\N__14304\&\N__14553\&\N__14808\&\N__15069\&\N__15306\&\N__20328\&\N__13689\&\N__15864\&\N__16119\;
    \line_buffer.mem16_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem16_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8088\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8862\&'0'&'0'&'0';
    \line_buffer.n574\ <= \line_buffer.mem30_physical_RDATA_wire\(11);
    \line_buffer.n573\ <= \line_buffer.mem30_physical_RDATA_wire\(3);
    \line_buffer.mem30_physical_RADDR_wire\ <= \N__12372\&\N__17190\&\N__18789\&\N__12666\&\N__12918\&\N__10335\&\N__10746\&\N__18096\&\N__18438\&\N__11688\&\N__11931\;
    \line_buffer.mem30_physical_WADDR_wire\ <= \N__15570\&\N__14052\&\N__14295\&\N__14550\&\N__14799\&\N__15066\&\N__15303\&\N__20325\&\N__13686\&\N__15861\&\N__16128\;
    \line_buffer.mem30_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem30_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8314\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8201\&'0'&'0'&'0';
    \line_buffer.n441\ <= \line_buffer.mem7_physical_RDATA_wire\(11);
    \line_buffer.n440\ <= \line_buffer.mem7_physical_RDATA_wire\(3);
    \line_buffer.mem7_physical_RADDR_wire\ <= \N__12312\&\N__17130\&\N__18729\&\N__12606\&\N__12858\&\N__10275\&\N__10686\&\N__18036\&\N__18378\&\N__11628\&\N__11871\;
    \line_buffer.mem7_physical_WADDR_wire\ <= \N__15510\&\N__13992\&\N__14235\&\N__14490\&\N__14739\&\N__15006\&\N__15243\&\N__20265\&\N__13626\&\N__15801\&\N__16068\;
    \line_buffer.mem7_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem7_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8644\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8755\&'0'&'0'&'0';
    \line_buffer.n568\ <= \line_buffer.mem20_physical_RDATA_wire\(11);
    \line_buffer.n567\ <= \line_buffer.mem20_physical_RDATA_wire\(3);
    \line_buffer.mem20_physical_RADDR_wire\ <= \N__12321\&\N__17127\&\N__18738\&\N__12609\&\N__12873\&\N__10296\&\N__10671\&\N__18039\&\N__18387\&\N__11637\&\N__11880\;
    \line_buffer.mem20_physical_WADDR_wire\ <= \N__15501\&\N__13983\&\N__14244\&\N__14493\&\N__14748\&\N__15009\&\N__15246\&\N__20268\&\N__13629\&\N__15804\&\N__16059\;
    \line_buffer.mem20_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem20_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8544\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8431\&'0'&'0'&'0';
    \line_buffer.n500\ <= \line_buffer.mem13_physical_RDATA_wire\(11);
    \line_buffer.n499\ <= \line_buffer.mem13_physical_RDATA_wire\(3);
    \line_buffer.mem13_physical_RADDR_wire\ <= \N__12417\&\N__17223\&\N__18834\&\N__12705\&\N__12969\&\N__10392\&\N__10767\&\N__18135\&\N__18483\&\N__11733\&\N__11976\;
    \line_buffer.mem13_physical_WADDR_wire\ <= \N__15597\&\N__14079\&\N__14340\&\N__14589\&\N__14844\&\N__15105\&\N__15342\&\N__20364\&\N__13725\&\N__15900\&\N__16155\;
    \line_buffer.mem13_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem13_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8057\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8855\&'0'&'0'&'0';
    \line_buffer.n443\ <= \line_buffer.mem19_physical_RDATA_wire\(11);
    \line_buffer.n442\ <= \line_buffer.mem19_physical_RDATA_wire\(3);
    \line_buffer.mem19_physical_RADDR_wire\ <= \N__12345\&\N__17151\&\N__18762\&\N__12633\&\N__12897\&\N__10320\&\N__10695\&\N__18063\&\N__18411\&\N__11661\&\N__11904\;
    \line_buffer.mem19_physical_WADDR_wire\ <= \N__15525\&\N__14007\&\N__14268\&\N__14517\&\N__14772\&\N__15033\&\N__15270\&\N__20292\&\N__13653\&\N__15828\&\N__16083\;
    \line_buffer.mem19_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem19_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8071\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8874\&'0'&'0'&'0';
    \line_buffer.n512\ <= \line_buffer.mem23_physical_RDATA_wire\(11);
    \line_buffer.n511\ <= \line_buffer.mem23_physical_RDATA_wire\(3);
    \line_buffer.mem23_physical_RADDR_wire\ <= \N__12468\&\N__17284\&\N__18885\&\N__12762\&\N__13014\&\N__10431\&\N__10834\&\N__18192\&\N__18534\&\N__11784\&\N__12027\;
    \line_buffer.mem23_physical_WADDR_wire\ <= \N__15661\&\N__14143\&\N__14391\&\N__14646\&\N__14895\&\N__15162\&\N__15399\&\N__20421\&\N__13782\&\N__15957\&\N__16219\;
    \line_buffer.mem23_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem23_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8516\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8357\&'0'&'0'&'0';
    \line_buffer.n506\ <= \line_buffer.mem0_physical_RDATA_wire\(11);
    \line_buffer.n505\ <= \line_buffer.mem0_physical_RDATA_wire\(3);
    \line_buffer.mem0_physical_RADDR_wire\ <= \N__12472\&\N__17283\&\N__18889\&\N__12763\&\N__13021\&\N__10441\&\N__10827\&\N__18193\&\N__18538\&\N__11788\&\N__12031\;
    \line_buffer.mem0_physical_WADDR_wire\ <= \N__15657\&\N__14139\&\N__14395\&\N__14647\&\N__14899\&\N__15163\&\N__15400\&\N__20422\&\N__13783\&\N__15958\&\N__16215\;
    \line_buffer.mem0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8572\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8711\&'0'&'0'&'0';
    \line_buffer.n544\ <= \line_buffer.mem26_physical_RDATA_wire\(11);
    \line_buffer.n543\ <= \line_buffer.mem26_physical_RDATA_wire\(3);
    \line_buffer.mem26_physical_RADDR_wire\ <= \N__12432\&\N__17250\&\N__18849\&\N__12726\&\N__12978\&\N__10395\&\N__10806\&\N__18156\&\N__18498\&\N__11748\&\N__11991\;
    \line_buffer.mem26_physical_WADDR_wire\ <= \N__15630\&\N__14112\&\N__14355\&\N__14610\&\N__14859\&\N__15126\&\N__15363\&\N__20385\&\N__13746\&\N__15921\&\N__16188\;
    \line_buffer.mem26_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem26_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8500\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8382\&'0'&'0'&'0';
    \line_buffer.n570\ <= \line_buffer.mem3_physical_RDATA_wire\(11);
    \line_buffer.n569\ <= \line_buffer.mem3_physical_RDATA_wire\(3);
    \line_buffer.mem3_physical_RADDR_wire\ <= \N__12384\&\N__17202\&\N__18801\&\N__12678\&\N__12930\&\N__10347\&\N__10758\&\N__18108\&\N__18450\&\N__11700\&\N__11943\;
    \line_buffer.mem3_physical_WADDR_wire\ <= \N__15582\&\N__14064\&\N__14307\&\N__14562\&\N__14811\&\N__15078\&\N__15315\&\N__20337\&\N__13698\&\N__15873\&\N__16140\;
    \line_buffer.mem3_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem3_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8628\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8727\&'0'&'0'&'0';
    \line_buffer.n447\ <= \line_buffer.mem17_physical_RDATA_wire\(11);
    \line_buffer.n446\ <= \line_buffer.mem17_physical_RDATA_wire\(3);
    \line_buffer.mem17_physical_RADDR_wire\ <= \N__12369\&\N__17175\&\N__18786\&\N__12657\&\N__12921\&\N__10344\&\N__10719\&\N__18087\&\N__18435\&\N__11685\&\N__11928\;
    \line_buffer.mem17_physical_WADDR_wire\ <= \N__15549\&\N__14031\&\N__14292\&\N__14541\&\N__14796\&\N__15057\&\N__15294\&\N__20316\&\N__13677\&\N__15852\&\N__16107\;
    \line_buffer.mem17_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem17_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8532\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8420\&'0'&'0'&'0';
    \line_buffer.n572\ <= \line_buffer.mem31_physical_RDATA_wire\(11);
    \line_buffer.n571\ <= \line_buffer.mem31_physical_RDATA_wire\(3);
    \line_buffer.mem31_physical_RADDR_wire\ <= \N__12360\&\N__17178\&\N__18777\&\N__12654\&\N__12906\&\N__10323\&\N__10734\&\N__18084\&\N__18426\&\N__11676\&\N__11919\;
    \line_buffer.mem31_physical_WADDR_wire\ <= \N__15558\&\N__14040\&\N__14283\&\N__14538\&\N__14787\&\N__15054\&\N__15291\&\N__20313\&\N__13674\&\N__15849\&\N__16116\;
    \line_buffer.mem31_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem31_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8061\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8840\&'0'&'0'&'0';
    \line_buffer.n437\ <= \line_buffer.mem9_physical_RDATA_wire\(11);
    \line_buffer.n436\ <= \line_buffer.mem9_physical_RDATA_wire\(3);
    \line_buffer.mem9_physical_RADDR_wire\ <= \N__12288\&\N__17106\&\N__18705\&\N__12582\&\N__12834\&\N__10251\&\N__10662\&\N__18012\&\N__18354\&\N__11604\&\N__11847\;
    \line_buffer.mem9_physical_WADDR_wire\ <= \N__15486\&\N__13964\&\N__14211\&\N__14466\&\N__14715\&\N__14978\&\N__15219\&\N__20241\&\N__13602\&\N__15777\&\N__16044\;
    \line_buffer.mem9_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem9_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8329\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8212\&'0'&'0'&'0';
    \line_buffer.n576\ <= \line_buffer.mem29_physical_RDATA_wire\(11);
    \line_buffer.n575\ <= \line_buffer.mem29_physical_RDATA_wire\(3);
    \line_buffer.mem29_physical_RADDR_wire\ <= \N__12396\&\N__17214\&\N__18813\&\N__12690\&\N__12942\&\N__10359\&\N__10770\&\N__18120\&\N__18462\&\N__11712\&\N__11955\;
    \line_buffer.mem29_physical_WADDR_wire\ <= \N__15594\&\N__14076\&\N__14319\&\N__14574\&\N__14823\&\N__15090\&\N__15327\&\N__20349\&\N__13710\&\N__15885\&\N__16152\;
    \line_buffer.mem29_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem29_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8533\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8395\&'0'&'0'&'0';
    \line_buffer.n578\ <= \line_buffer.mem6_physical_RDATA_wire\(11);
    \line_buffer.n577\ <= \line_buffer.mem6_physical_RDATA_wire\(3);
    \line_buffer.mem6_physical_RADDR_wire\ <= \N__12324\&\N__17142\&\N__18741\&\N__12618\&\N__12870\&\N__10287\&\N__10698\&\N__18048\&\N__18390\&\N__11640\&\N__11883\;
    \line_buffer.mem6_physical_WADDR_wire\ <= \N__15522\&\N__14004\&\N__14247\&\N__14502\&\N__14751\&\N__15018\&\N__15255\&\N__20277\&\N__13638\&\N__15813\&\N__16080\;
    \line_buffer.mem6_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem6_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8640\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8754\&'0'&'0'&'0';
    \line_buffer.n435\ <= \line_buffer.mem10_physical_RDATA_wire\(11);
    \line_buffer.n434\ <= \line_buffer.mem10_physical_RDATA_wire\(3);
    \line_buffer.mem10_physical_RADDR_wire\ <= \N__12453\&\N__17259\&\N__18870\&\N__12741\&\N__13005\&\N__10428\&\N__10803\&\N__18171\&\N__18519\&\N__11769\&\N__12012\;
    \line_buffer.mem10_physical_WADDR_wire\ <= \N__15633\&\N__14115\&\N__14376\&\N__14625\&\N__14880\&\N__15141\&\N__15378\&\N__20400\&\N__13761\&\N__15936\&\N__16191\;
    \line_buffer.mem10_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem10_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8081\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8841\&'0'&'0'&'0';
    \line_buffer.n564\ <= \line_buffer.mem22_physical_RDATA_wire\(11);
    \line_buffer.n563\ <= \line_buffer.mem22_physical_RDATA_wire\(3);
    \line_buffer.mem22_physical_RADDR_wire\ <= \N__12297\&\N__17103\&\N__18714\&\N__12585\&\N__12849\&\N__10272\&\N__10647\&\N__18015\&\N__18363\&\N__11613\&\N__11856\;
    \line_buffer.mem22_physical_WADDR_wire\ <= \N__15476\&\N__13952\&\N__14220\&\N__14469\&\N__14724\&\N__14984\&\N__15222\&\N__20244\&\N__13605\&\N__15780\&\N__16035\;
    \line_buffer.mem22_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem22_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8089\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8881\&'0'&'0'&'0';
    \line_buffer.n508\ <= \line_buffer.mem25_physical_RDATA_wire\(11);
    \line_buffer.n507\ <= \line_buffer.mem25_physical_RDATA_wire\(3);
    \line_buffer.mem25_physical_RADDR_wire\ <= \N__12444\&\N__17262\&\N__18861\&\N__12738\&\N__12990\&\N__10407\&\N__10818\&\N__18168\&\N__18510\&\N__11760\&\N__12003\;
    \line_buffer.mem25_physical_WADDR_wire\ <= \N__15642\&\N__14124\&\N__14367\&\N__14622\&\N__14871\&\N__15138\&\N__15375\&\N__20397\&\N__13758\&\N__15933\&\N__16200\;
    \line_buffer.mem25_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem25_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8056\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8809\&'0'&'0'&'0';
    \line_buffer.n439\ <= \line_buffer.mem8_physical_RDATA_wire\(11);
    \line_buffer.n438\ <= \line_buffer.mem8_physical_RDATA_wire\(3);
    \line_buffer.mem8_physical_RADDR_wire\ <= \N__12300\&\N__17118\&\N__18717\&\N__12594\&\N__12846\&\N__10263\&\N__10674\&\N__18024\&\N__18366\&\N__11616\&\N__11859\;
    \line_buffer.mem8_physical_WADDR_wire\ <= \N__15498\&\N__13980\&\N__14223\&\N__14478\&\N__14727\&\N__14994\&\N__15231\&\N__20253\&\N__13614\&\N__15789\&\N__16056\;
    \line_buffer.mem8_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem8_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8551\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8430\&'0'&'0'&'0';
    \line_buffer.n540\ <= \line_buffer.mem28_physical_RDATA_wire\(11);
    \line_buffer.n539\ <= \line_buffer.mem28_physical_RDATA_wire\(3);
    \line_buffer.mem28_physical_RADDR_wire\ <= \N__12408\&\N__17226\&\N__18825\&\N__12702\&\N__12954\&\N__10371\&\N__10782\&\N__18132\&\N__18474\&\N__11724\&\N__11967\;
    \line_buffer.mem28_physical_WADDR_wire\ <= \N__15606\&\N__14088\&\N__14331\&\N__14586\&\N__14835\&\N__15102\&\N__15339\&\N__20361\&\N__13722\&\N__15897\&\N__16164\;
    \line_buffer.mem28_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem28_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8037\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8822\&'0'&'0'&'0';

    \tx_pll.TX_PLL_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "010",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "100",
            DIVF => "0100110",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            LATCHINPUTVALUE => '0',
            SCLK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => \ADV_CLK_c\,
            REFERENCECLK => \N__18664\,
            RESETB => \N__19656\,
            BYPASS => \GNDG0\,
            SDI => '0',
            DYNAMICDELAY => \tx_pll.TX_PLL_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => OPEN
        );

    \line_buffer.mem2_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_E => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_D => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_C => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_B => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_A => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_9 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_8 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_7 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_6 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_5 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_4 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_3 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_2 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_1 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_0 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001"
        )
    port map (
            RDATA => \line_buffer.mem2_physical_RDATA_wire\,
            RADDR => \line_buffer.mem2_physical_RADDR_wire\,
            WADDR => \line_buffer.mem2_physical_WADDR_wire\,
            MASK => \line_buffer.mem2_physical_MASK_wire\,
            WDATA => \line_buffer.mem2_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22913\,
            RE => \N__19629\,
            WCLKE => 'H',
            WCLK => \N__20171\,
            WE => \N__16447\
        );

    \line_buffer.mem14_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_E => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_D => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_C => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_B => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_A => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_9 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_8 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_7 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_6 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_5 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_4 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_3 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011",
            INIT_2 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011",
            INIT_1 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011",
            INIT_0 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011"
        )
    port map (
            RDATA => \line_buffer.mem14_physical_RDATA_wire\,
            RADDR => \line_buffer.mem14_physical_RADDR_wire\,
            WADDR => \line_buffer.mem14_physical_WADDR_wire\,
            MASK => \line_buffer.mem14_physical_MASK_wire\,
            WDATA => \line_buffer.mem14_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23251\,
            RE => \N__19791\,
            WCLKE => 'H',
            WCLK => \N__20154\,
            WE => \N__16397\
        );

    \line_buffer.mem5_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_E => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_D => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_C => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_B => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_A => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_9 => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_8 => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_7 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_6 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_5 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_4 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_3 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110",
            INIT_2 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110",
            INIT_1 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110",
            INIT_0 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110"
        )
    port map (
            RDATA => \line_buffer.mem5_physical_RDATA_wire\,
            RADDR => \line_buffer.mem5_physical_RADDR_wire\,
            WADDR => \line_buffer.mem5_physical_WADDR_wire\,
            MASK => \line_buffer.mem5_physical_MASK_wire\,
            WDATA => \line_buffer.mem5_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22497\,
            RE => \N__19705\,
            WCLKE => 'H',
            WCLK => \N__20166\,
            WE => \N__16987\
        );

    \line_buffer.mem11_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_E => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_D => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_C => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_B => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_A => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_9 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_8 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_7 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_6 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_5 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_4 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_3 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_2 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_1 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_0 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100"
        )
    port map (
            RDATA => \line_buffer.mem11_physical_RDATA_wire\,
            RADDR => \line_buffer.mem11_physical_RADDR_wire\,
            WADDR => \line_buffer.mem11_physical_WADDR_wire\,
            MASK => \line_buffer.mem11_physical_MASK_wire\,
            WDATA => \line_buffer.mem11_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23293\,
            RE => \N__19819\,
            WCLKE => 'H',
            WCLK => \N__20146\,
            WE => \N__16935\
        );

    \line_buffer.mem21_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_E => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_D => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_C => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_B => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_A => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_9 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_8 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_7 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_6 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_5 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_4 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_3 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_2 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_1 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_0 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011"
        )
    port map (
            RDATA => \line_buffer.mem21_physical_RDATA_wire\,
            RADDR => \line_buffer.mem21_physical_RADDR_wire\,
            WADDR => \line_buffer.mem21_physical_WADDR_wire\,
            MASK => \line_buffer.mem21_physical_MASK_wire\,
            WDATA => \line_buffer.mem21_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22770\,
            RE => \N__19700\,
            WCLKE => 'H',
            WCLK => \N__20175\,
            WE => \N__16638\
        );

    \line_buffer.mem12_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_E => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_D => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_C => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_B => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_A => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_9 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_8 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_7 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_6 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_5 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_4 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_3 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_2 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_1 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_0 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100"
        )
    port map (
            RDATA => \line_buffer.mem12_physical_RDATA_wire\,
            RADDR => \line_buffer.mem12_physical_RADDR_wire\,
            WADDR => \line_buffer.mem12_physical_WADDR_wire\,
            MASK => \line_buffer.mem12_physical_MASK_wire\,
            WDATA => \line_buffer.mem12_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23279\,
            RE => \N__19818\,
            WCLKE => 'H',
            WCLK => \N__20148\,
            WE => \N__16928\
        );

    \line_buffer.mem18_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_E => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_D => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_C => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_B => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_A => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_9 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_8 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_7 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_6 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_5 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_4 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_3 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_2 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_1 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_0 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001"
        )
    port map (
            RDATA => \line_buffer.mem18_physical_RDATA_wire\,
            RADDR => \line_buffer.mem18_physical_RADDR_wire\,
            WADDR => \line_buffer.mem18_physical_WADDR_wire\,
            MASK => \line_buffer.mem18_physical_MASK_wire\,
            WDATA => \line_buffer.mem18_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23027\,
            RE => \N__19723\,
            WCLKE => 'H',
            WCLK => \N__20163\,
            WE => \N__16439\
        );

    \line_buffer.mem24_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_E => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_D => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_C => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_B => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_A => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_9 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_8 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_7 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_6 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_5 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_4 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_3 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_2 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_1 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_0 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001"
        )
    port map (
            RDATA => \line_buffer.mem24_physical_RDATA_wire\,
            RADDR => \line_buffer.mem24_physical_RADDR_wire\,
            WADDR => \line_buffer.mem24_physical_WADDR_wire\,
            MASK => \line_buffer.mem24_physical_MASK_wire\,
            WDATA => \line_buffer.mem24_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23271\,
            RE => \N__19855\,
            WCLKE => 'H',
            WCLK => \N__20138\,
            WE => \N__16491\
        );

    \line_buffer.mem1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_E => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_D => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_C => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_B => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_A => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_9 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_8 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_7 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_6 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_5 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_4 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_3 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011",
            INIT_2 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011",
            INIT_1 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011",
            INIT_0 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011"
        )
    port map (
            RDATA => \line_buffer.mem1_physical_RDATA_wire\,
            RADDR => \line_buffer.mem1_physical_RADDR_wire\,
            WADDR => \line_buffer.mem1_physical_WADDR_wire\,
            MASK => \line_buffer.mem1_physical_MASK_wire\,
            WDATA => \line_buffer.mem1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23301\,
            RE => \N__19839\,
            WCLKE => 'H',
            WCLK => \N__20136\,
            WE => \N__16396\
        );

    \line_buffer.mem15_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_E => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_D => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_C => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_B => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_A => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_9 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_8 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_7 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_6 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_5 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_4 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_3 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011",
            INIT_2 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011",
            INIT_1 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011",
            INIT_0 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011"
        )
    port map (
            RDATA => \line_buffer.mem15_physical_RDATA_wire\,
            RADDR => \line_buffer.mem15_physical_RADDR_wire\,
            WADDR => \line_buffer.mem15_physical_WADDR_wire\,
            MASK => \line_buffer.mem15_physical_MASK_wire\,
            WDATA => \line_buffer.mem15_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23200\,
            RE => \N__19759\,
            WCLKE => 'H',
            WCLK => \N__20156\,
            WE => \N__16404\
        );

    \line_buffer.mem27_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_E => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_D => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_C => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_B => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_A => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_9 => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_8 => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_7 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_6 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_5 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_4 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_3 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110",
            INIT_2 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110",
            INIT_1 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110",
            INIT_0 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110"
        )
    port map (
            RDATA => \line_buffer.mem27_physical_RDATA_wire\,
            RADDR => \line_buffer.mem27_physical_RADDR_wire\,
            WADDR => \line_buffer.mem27_physical_WADDR_wire\,
            MASK => \line_buffer.mem27_physical_MASK_wire\,
            WDATA => \line_buffer.mem27_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23270\,
            RE => \N__19829\,
            WCLKE => 'H',
            WCLK => \N__20149\,
            WE => \N__16976\
        );

    \line_buffer.mem4_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_E => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_D => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_C => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_B => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_A => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_9 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_8 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_7 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_6 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_5 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_4 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_3 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_2 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_1 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_0 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001"
        )
    port map (
            RDATA => \line_buffer.mem4_physical_RDATA_wire\,
            RADDR => \line_buffer.mem4_physical_RADDR_wire\,
            WADDR => \line_buffer.mem4_physical_WADDR_wire\,
            MASK => \line_buffer.mem4_physical_MASK_wire\,
            WDATA => \line_buffer.mem4_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22882\,
            RE => \N__19743\,
            WCLKE => 'H',
            WCLK => \N__20164\,
            WE => \N__16490\
        );

    \line_buffer.mem16_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_E => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_D => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_C => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_B => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_A => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_9 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_8 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_7 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_6 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_5 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_4 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_3 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011",
            INIT_2 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011",
            INIT_1 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011",
            INIT_0 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011"
        )
    port map (
            RDATA => \line_buffer.mem16_physical_RDATA_wire\,
            RADDR => \line_buffer.mem16_physical_RADDR_wire\,
            WADDR => \line_buffer.mem16_physical_WADDR_wire\,
            MASK => \line_buffer.mem16_physical_MASK_wire\,
            WDATA => \line_buffer.mem16_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23159\,
            RE => \N__19758\,
            WCLKE => 'H',
            WCLK => \N__20159\,
            WE => \N__16405\
        );

    \line_buffer.mem30_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_E => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_D => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_C => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_B => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_A => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_9 => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_8 => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_7 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_6 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_5 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_4 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_3 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110",
            INIT_2 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110",
            INIT_1 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110",
            INIT_0 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110"
        )
    port map (
            RDATA => \line_buffer.mem30_physical_RDATA_wire\,
            RADDR => \line_buffer.mem30_physical_RADDR_wire\,
            WADDR => \line_buffer.mem30_physical_WADDR_wire\,
            MASK => \line_buffer.mem30_physical_MASK_wire\,
            WDATA => \line_buffer.mem30_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23152\,
            RE => \N__19807\,
            WCLKE => 'H',
            WCLK => \N__20160\,
            WE => \N__16817\
        );

    \line_buffer.mem7_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_E => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_D => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_C => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_B => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_A => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_9 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_8 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_7 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_6 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_5 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_4 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_3 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_2 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_1 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_0 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000"
        )
    port map (
            RDATA => \line_buffer.mem7_physical_RDATA_wire\,
            RADDR => \line_buffer.mem7_physical_RADDR_wire\,
            WADDR => \line_buffer.mem7_physical_WADDR_wire\,
            MASK => \line_buffer.mem7_physical_MASK_wire\,
            WDATA => \line_buffer.mem7_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22530\,
            RE => \N__19718\,
            WCLKE => 'H',
            WCLK => \N__20174\,
            WE => \N__17033\
        );

    \line_buffer.mem20_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_E => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_D => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_C => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_B => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_A => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_9 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_8 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_7 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_6 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_5 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_4 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_3 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_2 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_1 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_0 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011"
        )
    port map (
            RDATA => \line_buffer.mem20_physical_RDATA_wire\,
            RADDR => \line_buffer.mem20_physical_RADDR_wire\,
            WADDR => \line_buffer.mem20_physical_WADDR_wire\,
            MASK => \line_buffer.mem20_physical_MASK_wire\,
            WDATA => \line_buffer.mem20_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22912\,
            RE => \N__19699\,
            WCLKE => 'H',
            WCLK => \N__20173\,
            WE => \N__16634\
        );

    \line_buffer.mem13_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_E => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_D => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_C => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_B => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_A => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_9 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_8 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_7 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_6 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_5 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_4 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_3 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_2 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_1 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_0 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100"
        )
    port map (
            RDATA => \line_buffer.mem13_physical_RDATA_wire\,
            RADDR => \line_buffer.mem13_physical_RADDR_wire\,
            WADDR => \line_buffer.mem13_physical_WADDR_wire\,
            MASK => \line_buffer.mem13_physical_MASK_wire\,
            WDATA => \line_buffer.mem13_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23278\,
            RE => \N__19792\,
            WCLKE => 'H',
            WCLK => \N__20150\,
            WE => \N__16908\
        );

    \line_buffer.mem19_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_E => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_D => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_C => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_B => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_A => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_9 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_8 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_7 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_6 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_5 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_4 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_3 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_2 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_1 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_0 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001"
        )
    port map (
            RDATA => \line_buffer.mem19_physical_RDATA_wire\,
            RADDR => \line_buffer.mem19_physical_RADDR_wire\,
            WADDR => \line_buffer.mem19_physical_WADDR_wire\,
            MASK => \line_buffer.mem19_physical_MASK_wire\,
            WDATA => \line_buffer.mem19_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23026\,
            RE => \N__19680\,
            WCLKE => 'H',
            WCLK => \N__20165\,
            WE => \N__16446\
        );

    \line_buffer.mem23_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_E => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_D => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_C => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_B => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_A => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_9 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_8 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_7 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_6 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_5 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_4 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_3 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_2 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_1 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_0 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001"
        )
    port map (
            RDATA => \line_buffer.mem23_physical_RDATA_wire\,
            RADDR => \line_buffer.mem23_physical_RADDR_wire\,
            WADDR => \line_buffer.mem23_physical_WADDR_wire\,
            MASK => \line_buffer.mem23_physical_MASK_wire\,
            WDATA => \line_buffer.mem23_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23272\,
            RE => \N__19704\,
            WCLKE => 'H',
            WCLK => \N__20134\,
            WE => \N__16492\
        );

    \line_buffer.mem0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_E => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_D => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_C => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_B => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_A => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_9 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_8 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_7 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_6 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_5 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_4 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_3 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_2 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_1 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_0 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100"
        )
    port map (
            RDATA => \line_buffer.mem0_physical_RDATA_wire\,
            RADDR => \line_buffer.mem0_physical_RADDR_wire\,
            WADDR => \line_buffer.mem0_physical_WADDR_wire\,
            MASK => \line_buffer.mem0_physical_MASK_wire\,
            WDATA => \line_buffer.mem0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23302\,
            RE => \N__19850\,
            WCLKE => 'H',
            WCLK => \N__20132\,
            WE => \N__16939\
        );

    \line_buffer.mem26_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_E => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_D => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_C => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_B => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_A => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_9 => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_8 => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_7 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_6 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_5 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_4 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_3 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110",
            INIT_2 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110",
            INIT_1 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110",
            INIT_0 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110"
        )
    port map (
            RDATA => \line_buffer.mem26_physical_RDATA_wire\,
            RADDR => \line_buffer.mem26_physical_RADDR_wire\,
            WADDR => \line_buffer.mem26_physical_WADDR_wire\,
            MASK => \line_buffer.mem26_physical_MASK_wire\,
            WDATA => \line_buffer.mem26_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22649\,
            RE => \N__19843\,
            WCLKE => 'H',
            WCLK => \N__20147\,
            WE => \N__16986\
        );

    \line_buffer.mem3_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_E => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_D => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_C => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_B => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_A => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_9 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_8 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_7 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_6 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_5 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_4 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_3 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_2 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_1 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_0 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011"
        )
    port map (
            RDATA => \line_buffer.mem3_physical_RDATA_wire\,
            RADDR => \line_buffer.mem3_physical_RADDR_wire\,
            WADDR => \line_buffer.mem3_physical_WADDR_wire\,
            MASK => \line_buffer.mem3_physical_MASK_wire\,
            WDATA => \line_buffer.mem3_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23078\,
            RE => \N__19808\,
            WCLKE => 'H',
            WCLK => \N__20157\,
            WE => \N__16624\
        );

    \line_buffer.mem17_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_E => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_D => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_C => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_B => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_A => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_9 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_8 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_7 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_6 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_5 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_4 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_3 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_2 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_1 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_0 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001"
        )
    port map (
            RDATA => \line_buffer.mem17_physical_RDATA_wire\,
            RADDR => \line_buffer.mem17_physical_RADDR_wire\,
            WADDR => \line_buffer.mem17_physical_WADDR_wire\,
            MASK => \line_buffer.mem17_physical_MASK_wire\,
            WDATA => \line_buffer.mem17_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23106\,
            RE => \N__19724\,
            WCLKE => 'H',
            WCLK => \N__20161\,
            WE => \N__16438\
        );

    \line_buffer.mem31_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_E => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_D => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_C => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_B => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_A => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_9 => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_8 => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_7 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_6 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_5 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_4 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_3 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110",
            INIT_2 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110",
            INIT_1 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110",
            INIT_0 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110"
        )
    port map (
            RDATA => \line_buffer.mem31_physical_RDATA_wire\,
            RADDR => \line_buffer.mem31_physical_RADDR_wire\,
            WADDR => \line_buffer.mem31_physical_WADDR_wire\,
            MASK => \line_buffer.mem31_physical_MASK_wire\,
            WDATA => \line_buffer.mem31_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22545\,
            RE => \N__19776\,
            WCLKE => 'H',
            WCLK => \N__20162\,
            WE => \N__16824\
        );

    \line_buffer.mem9_physical\ : SB_RAM40_4K
    generic map (
            INIT_0 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_E => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_D => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_C => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_B => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_A => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_9 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_8 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_7 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_6 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_5 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_4 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_3 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_2 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_1 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000"
        )
    port map (
            RDATA => \line_buffer.mem9_physical_RDATA_wire\,
            RADDR => \line_buffer.mem9_physical_RADDR_wire\,
            WADDR => \line_buffer.mem9_physical_WADDR_wire\,
            MASK => \line_buffer.mem9_physical_MASK_wire\,
            WDATA => \line_buffer.mem9_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22461\,
            RE => \N__19757\,
            WCLKE => 'H',
            WCLK => \N__20178\,
            WE => \N__17041\
        );

    \line_buffer.mem29_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_E => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_D => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_C => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_B => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_A => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_9 => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_8 => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_7 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_6 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_5 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_4 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_3 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110",
            INIT_2 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110",
            INIT_1 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110",
            INIT_0 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110"
        )
    port map (
            RDATA => \line_buffer.mem29_physical_RDATA_wire\,
            RADDR => \line_buffer.mem29_physical_RADDR_wire\,
            WADDR => \line_buffer.mem29_physical_WADDR_wire\,
            MASK => \line_buffer.mem29_physical_MASK_wire\,
            WDATA => \line_buffer.mem29_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23202\,
            RE => \N__19652\,
            WCLKE => 'H',
            WCLK => \N__20155\,
            WE => \N__16808\
        );

    \line_buffer.mem6_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_E => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_D => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_C => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_B => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_A => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_9 => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_8 => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_7 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_6 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_5 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_4 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_3 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110",
            INIT_2 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110",
            INIT_1 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110",
            INIT_0 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110"
        )
    port map (
            RDATA => \line_buffer.mem6_physical_RDATA_wire\,
            RADDR => \line_buffer.mem6_physical_RADDR_wire\,
            WADDR => \line_buffer.mem6_physical_WADDR_wire\,
            MASK => \line_buffer.mem6_physical_MASK_wire\,
            WDATA => \line_buffer.mem6_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22746\,
            RE => \N__19602\,
            WCLKE => 'H',
            WCLK => \N__20172\,
            WE => \N__16828\
        );

    \line_buffer.mem10_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_E => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_D => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_C => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_B => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_A => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_9 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_8 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_7 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_6 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_5 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_4 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_3 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_2 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_1 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_0 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000"
        )
    port map (
            RDATA => \line_buffer.mem10_physical_RDATA_wire\,
            RADDR => \line_buffer.mem10_physical_RADDR_wire\,
            WADDR => \line_buffer.mem10_physical_WADDR_wire\,
            MASK => \line_buffer.mem10_physical_MASK_wire\,
            WDATA => \line_buffer.mem10_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23294\,
            RE => \N__19838\,
            WCLKE => 'H',
            WCLK => \N__20140\,
            WE => \N__17024\
        );

    \line_buffer.mem22_physical\ : SB_RAM40_4K
    generic map (
            INIT_0 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_E => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_D => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_C => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_B => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_A => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_9 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_8 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_7 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_6 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_5 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_4 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_3 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_2 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_1 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011"
        )
    port map (
            RDATA => \line_buffer.mem22_physical_RDATA_wire\,
            RADDR => \line_buffer.mem22_physical_RADDR_wire\,
            WADDR => \line_buffer.mem22_physical_WADDR_wire\,
            MASK => \line_buffer.mem22_physical_MASK_wire\,
            WDATA => \line_buffer.mem22_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22531\,
            RE => \N__19742\,
            WCLKE => 'H',
            WCLK => \N__20177\,
            WE => \N__16639\
        );

    \line_buffer.mem25_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_E => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_D => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_C => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_B => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_A => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_9 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_8 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_7 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_6 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_5 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_4 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_3 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_2 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_1 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_0 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001"
        )
    port map (
            RDATA => \line_buffer.mem25_physical_RDATA_wire\,
            RADDR => \line_buffer.mem25_physical_RADDR_wire\,
            WADDR => \line_buffer.mem25_physical_WADDR_wire\,
            MASK => \line_buffer.mem25_physical_MASK_wire\,
            WDATA => \line_buffer.mem25_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23235\,
            RE => \N__19851\,
            WCLKE => 'H',
            WCLK => \N__20144\,
            WE => \N__16483\
        );

    \line_buffer.mem8_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_E => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_D => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_C => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_B => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_A => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_9 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_8 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_7 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_6 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_5 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_4 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_3 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_2 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_1 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_0 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000"
        )
    port map (
            RDATA => \line_buffer.mem8_physical_RDATA_wire\,
            RADDR => \line_buffer.mem8_physical_RADDR_wire\,
            WADDR => \line_buffer.mem8_physical_WADDR_wire\,
            MASK => \line_buffer.mem8_physical_MASK_wire\,
            WDATA => \line_buffer.mem8_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22610\,
            RE => \N__19719\,
            WCLKE => 'H',
            WCLK => \N__20176\,
            WE => \N__17040\
        );

    \line_buffer.mem28_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_E => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_D => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_C => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_B => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_A => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_9 => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_8 => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_7 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_6 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_5 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_4 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_3 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110",
            INIT_2 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110",
            INIT_1 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110",
            INIT_0 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110"
        )
    port map (
            RDATA => \line_buffer.mem28_physical_RDATA_wire\,
            RADDR => \line_buffer.mem28_physical_RADDR_wire\,
            WADDR => \line_buffer.mem28_physical_WADDR_wire\,
            MASK => \line_buffer.mem28_physical_MASK_wire\,
            WDATA => \line_buffer.mem28_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23269\,
            RE => \N__19809\,
            WCLKE => 'H',
            WCLK => \N__20151\,
            WE => \N__16972\
        );

    \TVP_CLK_pad_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__24119\,
            GLOBALBUFFEROUTPUT => \TVP_CLK_c\
        );

    \TVP_CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24121\,
            DIN => \N__24120\,
            DOUT => \N__24119\,
            PACKAGEPIN => \TVP_CLK_wire\
        );

    \TVP_CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24121\,
            PADOUT => \N__24120\,
            PADIN => \N__24119\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24110\,
            DIN => \N__24109\,
            DOUT => \N__24108\,
            PACKAGEPIN => \ADV_CLK_wire\
        );

    \ADV_CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24110\,
            PADOUT => \N__24109\,
            PADIN => \N__24108\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__22632\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24101\,
            DIN => \N__24100\,
            DOUT => \N__24099\,
            PACKAGEPIN => DEBUG(3)
        );

    \DEBUG_pad_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24101\,
            PADOUT => \N__24100\,
            PADIN => \N__24099\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_VIDEO_pad_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24092\,
            DIN => \N__24091\,
            DOUT => \N__24090\,
            PACKAGEPIN => \TVP_VIDEO_wire\(2)
        );

    \TVP_VIDEO_pad_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24092\,
            PADOUT => \N__24091\,
            PADIN => \N__24090\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_VIDEO_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24083\,
            DIN => \N__24082\,
            DOUT => \N__24081\,
            PACKAGEPIN => \ADV_G_wire\(5)
        );

    \ADV_G_pad_5_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24083\,
            PADOUT => \N__24082\,
            PADIN => \N__24081\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__19905\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24074\,
            DIN => \N__24073\,
            DOUT => \N__24072\,
            PACKAGEPIN => \ADV_R_wire\(3)
        );

    \ADV_R_pad_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24074\,
            PADOUT => \N__24073\,
            PADIN => \N__24072\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__23424\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24065\,
            DIN => \N__24064\,
            DOUT => \N__24063\,
            PACKAGEPIN => DEBUG(7)
        );

    \DEBUG_pad_7_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24065\,
            PADOUT => \N__24064\,
            PADIN => \N__24063\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_VIDEO_pad_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24056\,
            DIN => \N__24055\,
            DOUT => \N__24054\,
            PACKAGEPIN => \TVP_VIDEO_wire\(6)
        );

    \TVP_VIDEO_pad_6_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24056\,
            PADOUT => \N__24055\,
            PADIN => \N__24054\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_VIDEO_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24047\,
            DIN => \N__24046\,
            DOUT => \N__24045\,
            PACKAGEPIN => \ADV_G_wire\(1)
        );

    \ADV_G_pad_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24047\,
            PADOUT => \N__24046\,
            PADIN => \N__24045\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__21559\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24038\,
            DIN => \N__24037\,
            DOUT => \N__24036\,
            PACKAGEPIN => \ADV_R_wire\(0)
        );

    \ADV_R_pad_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24038\,
            PADOUT => \N__24037\,
            PADIN => \N__24036\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12172\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24029\,
            DIN => \N__24028\,
            DOUT => \N__24027\,
            PACKAGEPIN => DEBUG(2)
        );

    \DEBUG_pad_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24029\,
            PADOUT => \N__24028\,
            PADIN => \N__24027\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_VIDEO_pad_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24020\,
            DIN => \N__24019\,
            DOUT => \N__24018\,
            PACKAGEPIN => \TVP_VIDEO_wire\(3)
        );

    \TVP_VIDEO_pad_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24020\,
            PADOUT => \N__24019\,
            PADIN => \N__24018\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_VIDEO_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24011\,
            DIN => \N__24010\,
            DOUT => \N__24009\,
            PACKAGEPIN => \ADV_G_wire\(4)
        );

    \ADV_G_pad_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24011\,
            PADOUT => \N__24010\,
            PADIN => \N__24009\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__17693\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24002\,
            DIN => \N__24001\,
            DOUT => \N__24000\,
            PACKAGEPIN => \ADV_R_wire\(5)
        );

    \ADV_R_pad_5_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24002\,
            PADOUT => \N__24001\,
            PADIN => \N__24000\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__19898\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_VIDEO_pad_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__23993\,
            DIN => \N__23992\,
            DOUT => \N__23991\,
            PACKAGEPIN => \TVP_VIDEO_wire\(9)
        );

    \TVP_VIDEO_pad_9_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23993\,
            PADOUT => \N__23992\,
            PADIN => \N__23991\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_VIDEO_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__23984\,
            DIN => \N__23983\,
            DOUT => \N__23982\,
            PACKAGEPIN => DEBUG(1)
        );

    \DEBUG_pad_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23984\,
            PADOUT => \N__23983\,
            PADIN => \N__23982\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23975\,
            DIN => \N__23974\,
            DOUT => \N__23973\,
            PACKAGEPIN => \ADV_B_wire\(1)
        );

    \ADV_B_pad_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23975\,
            PADOUT => \N__23974\,
            PADIN => \N__23973\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__21545\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_SYNC_N_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__23966\,
            DIN => \N__23965\,
            DOUT => \N__23964\,
            PACKAGEPIN => \ADV_SYNC_N_wire\
        );

    \ADV_SYNC_N_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23966\,
            PADOUT => \N__23965\,
            PADIN => \N__23964\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23957\,
            DIN => \N__23956\,
            DOUT => \N__23955\,
            PACKAGEPIN => \ADV_B_wire\(6)
        );

    \ADV_B_pad_6_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23957\,
            PADOUT => \N__23956\,
            PADIN => \N__23955\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12223\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__23948\,
            DIN => \N__23947\,
            DOUT => \N__23946\,
            PACKAGEPIN => DEBUG(6)
        );

    \DEBUG_pad_6_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23948\,
            PADOUT => \N__23947\,
            PADIN => \N__23946\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_VIDEO_pad_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__23939\,
            DIN => \N__23938\,
            DOUT => \N__23937\,
            PACKAGEPIN => \TVP_VIDEO_wire\(7)
        );

    \TVP_VIDEO_pad_7_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23939\,
            PADOUT => \N__23938\,
            PADIN => \N__23937\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_VIDEO_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23930\,
            DIN => \N__23929\,
            DOUT => \N__23928\,
            PACKAGEPIN => \ADV_G_wire\(0)
        );

    \ADV_G_pad_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23930\,
            PADOUT => \N__23929\,
            PADIN => \N__23928\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12167\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23921\,
            DIN => \N__23920\,
            DOUT => \N__23919\,
            PACKAGEPIN => \ADV_R_wire\(1)
        );

    \ADV_R_pad_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23921\,
            PADOUT => \N__23920\,
            PADIN => \N__23919\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__21558\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__23912\,
            DIN => \N__23911\,
            DOUT => \N__23910\,
            PACKAGEPIN => DEBUG(5)
        );

    \DEBUG_pad_5_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23912\,
            PADOUT => \N__23911\,
            PADIN => \N__23910\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_HSYNC_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__23903\,
            DIN => \N__23902\,
            DOUT => \N__23901\,
            PACKAGEPIN => \TVP_HSYNC_wire\
        );

    \TVP_HSYNC_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23903\,
            PADOUT => \N__23902\,
            PADIN => \N__23901\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_HSYNC_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23894\,
            DIN => \N__23893\,
            DOUT => \N__23892\,
            PACKAGEPIN => \ADV_G_wire\(7)
        );

    \ADV_G_pad_7_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23894\,
            PADOUT => \N__23893\,
            PADIN => \N__23892\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__23357\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23885\,
            DIN => \N__23884\,
            DOUT => \N__23883\,
            PACKAGEPIN => \ADV_R_wire\(6)
        );

    \ADV_R_pad_6_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23885\,
            PADOUT => \N__23884\,
            PADIN => \N__23883\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12215\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_VSYNC_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__23876\,
            DIN => \N__23875\,
            DOUT => \N__23874\,
            PACKAGEPIN => \TVP_VSYNC_wire\
        );

    \TVP_VSYNC_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23876\,
            PADOUT => \N__23875\,
            PADIN => \N__23874\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_VSYNC_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_BLANK_N_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__23867\,
            DIN => \N__23866\,
            DOUT => \N__23865\,
            PACKAGEPIN => \ADV_BLANK_N_wire\
        );

    \ADV_BLANK_N_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23867\,
            PADOUT => \N__23866\,
            PADIN => \N__23865\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__19657\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__23858\,
            DIN => \N__23857\,
            DOUT => \N__23856\,
            PACKAGEPIN => DEBUG(0)
        );

    \DEBUG_pad_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23858\,
            PADOUT => \N__23857\,
            PADIN => \N__23856\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23849\,
            DIN => \N__23848\,
            DOUT => \N__23847\,
            PACKAGEPIN => \ADV_B_wire\(2)
        );

    \ADV_B_pad_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23849\,
            PADOUT => \N__23848\,
            PADIN => \N__23847\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__17624\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23840\,
            DIN => \N__23839\,
            DOUT => \N__23838\,
            PACKAGEPIN => \ADV_B_wire\(7)
        );

    \ADV_B_pad_7_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23840\,
            PADOUT => \N__23839\,
            PADIN => \N__23838\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__23364\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LED_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__23831\,
            DIN => \N__23830\,
            DOUT => \N__23829\,
            PACKAGEPIN => \LED_wire\
        );

    \LED_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23831\,
            PADOUT => \N__23830\,
            PADIN => \N__23829\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12553\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_VIDEO_pad_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__23822\,
            DIN => \N__23821\,
            DOUT => \N__23820\,
            PACKAGEPIN => \TVP_VIDEO_wire\(4)
        );

    \TVP_VIDEO_pad_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23822\,
            PADOUT => \N__23821\,
            PADIN => \N__23820\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_VIDEO_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23813\,
            DIN => \N__23812\,
            DOUT => \N__23811\,
            PACKAGEPIN => \ADV_G_wire\(3)
        );

    \ADV_G_pad_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23813\,
            PADOUT => \N__23812\,
            PADIN => \N__23811\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__23434\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_HSYNC_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23804\,
            DIN => \N__23803\,
            DOUT => \N__23802\,
            PACKAGEPIN => \ADV_HSYNC_wire\
        );

    \ADV_HSYNC_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23804\,
            PADOUT => \N__23803\,
            PADIN => \N__23802\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10570\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23795\,
            DIN => \N__23794\,
            DOUT => \N__23793\,
            PACKAGEPIN => \ADV_R_wire\(2)
        );

    \ADV_R_pad_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23795\,
            PADOUT => \N__23794\,
            PADIN => \N__23793\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__17629\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23786\,
            DIN => \N__23785\,
            DOUT => \N__23784\,
            PACKAGEPIN => \ADV_B_wire\(4)
        );

    \ADV_B_pad_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23786\,
            PADOUT => \N__23785\,
            PADIN => \N__23784\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__17697\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__23777\,
            DIN => \N__23776\,
            DOUT => \N__23775\,
            PACKAGEPIN => DEBUG(4)
        );

    \DEBUG_pad_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23777\,
            PADOUT => \N__23776\,
            PADIN => \N__23775\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23768\,
            DIN => \N__23767\,
            DOUT => \N__23766\,
            PACKAGEPIN => \ADV_G_wire\(6)
        );

    \ADV_G_pad_6_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23768\,
            PADOUT => \N__23767\,
            PADIN => \N__23766\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12219\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23759\,
            DIN => \N__23758\,
            DOUT => \N__23757\,
            PACKAGEPIN => \ADV_R_wire\(7)
        );

    \ADV_R_pad_7_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23759\,
            PADOUT => \N__23758\,
            PADIN => \N__23757\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__23365\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23750\,
            DIN => \N__23749\,
            DOUT => \N__23748\,
            PACKAGEPIN => \ADV_B_wire\(3)
        );

    \ADV_B_pad_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23750\,
            PADOUT => \N__23749\,
            PADIN => \N__23748\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__23417\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23741\,
            DIN => \N__23740\,
            DOUT => \N__23739\,
            PACKAGEPIN => \ADV_R_wire\(4)
        );

    \ADV_R_pad_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23741\,
            PADOUT => \N__23740\,
            PADIN => \N__23739\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__17698\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_VIDEO_pad_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__23732\,
            DIN => \N__23731\,
            DOUT => \N__23730\,
            PACKAGEPIN => \TVP_VIDEO_wire\(8)
        );

    \TVP_VIDEO_pad_8_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23732\,
            PADOUT => \N__23731\,
            PADIN => \N__23730\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_VIDEO_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23723\,
            DIN => \N__23722\,
            DOUT => \N__23721\,
            PACKAGEPIN => \ADV_B_wire\(0)
        );

    \ADV_B_pad_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23723\,
            PADOUT => \N__23722\,
            PADIN => \N__23721\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12168\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_VIDEO_pad_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__23714\,
            DIN => \N__23713\,
            DOUT => \N__23712\,
            PACKAGEPIN => \TVP_VIDEO_wire\(5)
        );

    \TVP_VIDEO_pad_5_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23714\,
            PADOUT => \N__23713\,
            PADIN => \N__23712\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_VIDEO_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23705\,
            DIN => \N__23704\,
            DOUT => \N__23703\,
            PACKAGEPIN => \ADV_G_wire\(2)
        );

    \ADV_G_pad_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23705\,
            PADOUT => \N__23704\,
            PADIN => \N__23703\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__17628\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_VSYNC_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23696\,
            DIN => \N__23695\,
            DOUT => \N__23694\,
            PACKAGEPIN => \ADV_VSYNC_wire\
        );

    \ADV_VSYNC_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23696\,
            PADOUT => \N__23695\,
            PADIN => \N__23694\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__21352\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23687\,
            DIN => \N__23686\,
            DOUT => \N__23685\,
            PACKAGEPIN => \ADV_B_wire\(5)
        );

    \ADV_B_pad_5_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23687\,
            PADOUT => \N__23686\,
            PADIN => \N__23685\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__19909\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__5727\ : InMux
    port map (
            O => \N__23668\,
            I => \N__23660\
        );

    \I__5726\ : InMux
    port map (
            O => \N__23667\,
            I => \N__23656\
        );

    \I__5725\ : CascadeMux
    port map (
            O => \N__23666\,
            I => \N__23650\
        );

    \I__5724\ : InMux
    port map (
            O => \N__23665\,
            I => \N__23644\
        );

    \I__5723\ : InMux
    port map (
            O => \N__23664\,
            I => \N__23641\
        );

    \I__5722\ : InMux
    port map (
            O => \N__23663\,
            I => \N__23634\
        );

    \I__5721\ : LocalMux
    port map (
            O => \N__23660\,
            I => \N__23631\
        );

    \I__5720\ : InMux
    port map (
            O => \N__23659\,
            I => \N__23626\
        );

    \I__5719\ : LocalMux
    port map (
            O => \N__23656\,
            I => \N__23623\
        );

    \I__5718\ : InMux
    port map (
            O => \N__23655\,
            I => \N__23620\
        );

    \I__5717\ : InMux
    port map (
            O => \N__23654\,
            I => \N__23617\
        );

    \I__5716\ : InMux
    port map (
            O => \N__23653\,
            I => \N__23614\
        );

    \I__5715\ : InMux
    port map (
            O => \N__23650\,
            I => \N__23609\
        );

    \I__5714\ : InMux
    port map (
            O => \N__23649\,
            I => \N__23609\
        );

    \I__5713\ : InMux
    port map (
            O => \N__23648\,
            I => \N__23606\
        );

    \I__5712\ : InMux
    port map (
            O => \N__23647\,
            I => \N__23603\
        );

    \I__5711\ : LocalMux
    port map (
            O => \N__23644\,
            I => \N__23596\
        );

    \I__5710\ : LocalMux
    port map (
            O => \N__23641\,
            I => \N__23596\
        );

    \I__5709\ : InMux
    port map (
            O => \N__23640\,
            I => \N__23593\
        );

    \I__5708\ : InMux
    port map (
            O => \N__23639\,
            I => \N__23590\
        );

    \I__5707\ : InMux
    port map (
            O => \N__23638\,
            I => \N__23587\
        );

    \I__5706\ : InMux
    port map (
            O => \N__23637\,
            I => \N__23584\
        );

    \I__5705\ : LocalMux
    port map (
            O => \N__23634\,
            I => \N__23581\
        );

    \I__5704\ : Span4Mux_h
    port map (
            O => \N__23631\,
            I => \N__23578\
        );

    \I__5703\ : InMux
    port map (
            O => \N__23630\,
            I => \N__23575\
        );

    \I__5702\ : InMux
    port map (
            O => \N__23629\,
            I => \N__23571\
        );

    \I__5701\ : LocalMux
    port map (
            O => \N__23626\,
            I => \N__23564\
        );

    \I__5700\ : Span4Mux_h
    port map (
            O => \N__23623\,
            I => \N__23564\
        );

    \I__5699\ : LocalMux
    port map (
            O => \N__23620\,
            I => \N__23564\
        );

    \I__5698\ : LocalMux
    port map (
            O => \N__23617\,
            I => \N__23561\
        );

    \I__5697\ : LocalMux
    port map (
            O => \N__23614\,
            I => \N__23554\
        );

    \I__5696\ : LocalMux
    port map (
            O => \N__23609\,
            I => \N__23554\
        );

    \I__5695\ : LocalMux
    port map (
            O => \N__23606\,
            I => \N__23554\
        );

    \I__5694\ : LocalMux
    port map (
            O => \N__23603\,
            I => \N__23551\
        );

    \I__5693\ : InMux
    port map (
            O => \N__23602\,
            I => \N__23548\
        );

    \I__5692\ : InMux
    port map (
            O => \N__23601\,
            I => \N__23545\
        );

    \I__5691\ : Span4Mux_h
    port map (
            O => \N__23596\,
            I => \N__23536\
        );

    \I__5690\ : LocalMux
    port map (
            O => \N__23593\,
            I => \N__23536\
        );

    \I__5689\ : LocalMux
    port map (
            O => \N__23590\,
            I => \N__23536\
        );

    \I__5688\ : LocalMux
    port map (
            O => \N__23587\,
            I => \N__23529\
        );

    \I__5687\ : LocalMux
    port map (
            O => \N__23584\,
            I => \N__23529\
        );

    \I__5686\ : Span4Mux_h
    port map (
            O => \N__23581\,
            I => \N__23529\
        );

    \I__5685\ : Span4Mux_v
    port map (
            O => \N__23578\,
            I => \N__23524\
        );

    \I__5684\ : LocalMux
    port map (
            O => \N__23575\,
            I => \N__23524\
        );

    \I__5683\ : InMux
    port map (
            O => \N__23574\,
            I => \N__23521\
        );

    \I__5682\ : LocalMux
    port map (
            O => \N__23571\,
            I => \N__23516\
        );

    \I__5681\ : Span4Mux_v
    port map (
            O => \N__23564\,
            I => \N__23516\
        );

    \I__5680\ : Span4Mux_v
    port map (
            O => \N__23561\,
            I => \N__23507\
        );

    \I__5679\ : Span4Mux_v
    port map (
            O => \N__23554\,
            I => \N__23507\
        );

    \I__5678\ : Span4Mux_v
    port map (
            O => \N__23551\,
            I => \N__23507\
        );

    \I__5677\ : LocalMux
    port map (
            O => \N__23548\,
            I => \N__23507\
        );

    \I__5676\ : LocalMux
    port map (
            O => \N__23545\,
            I => \N__23504\
        );

    \I__5675\ : InMux
    port map (
            O => \N__23544\,
            I => \N__23501\
        );

    \I__5674\ : InMux
    port map (
            O => \N__23543\,
            I => \N__23498\
        );

    \I__5673\ : Span4Mux_v
    port map (
            O => \N__23536\,
            I => \N__23489\
        );

    \I__5672\ : Span4Mux_v
    port map (
            O => \N__23529\,
            I => \N__23489\
        );

    \I__5671\ : Span4Mux_v
    port map (
            O => \N__23524\,
            I => \N__23489\
        );

    \I__5670\ : LocalMux
    port map (
            O => \N__23521\,
            I => \N__23489\
        );

    \I__5669\ : Span4Mux_v
    port map (
            O => \N__23516\,
            I => \N__23484\
        );

    \I__5668\ : Span4Mux_h
    port map (
            O => \N__23507\,
            I => \N__23484\
        );

    \I__5667\ : Odrv4
    port map (
            O => \N__23504\,
            I => \TX_ADDR_11\
        );

    \I__5666\ : LocalMux
    port map (
            O => \N__23501\,
            I => \TX_ADDR_11\
        );

    \I__5665\ : LocalMux
    port map (
            O => \N__23498\,
            I => \TX_ADDR_11\
        );

    \I__5664\ : Odrv4
    port map (
            O => \N__23489\,
            I => \TX_ADDR_11\
        );

    \I__5663\ : Odrv4
    port map (
            O => \N__23484\,
            I => \TX_ADDR_11\
        );

    \I__5662\ : InMux
    port map (
            O => \N__23473\,
            I => \N__23470\
        );

    \I__5661\ : LocalMux
    port map (
            O => \N__23470\,
            I => \N__23467\
        );

    \I__5660\ : Span12Mux_v
    port map (
            O => \N__23467\,
            I => \N__23464\
        );

    \I__5659\ : Span12Mux_h
    port map (
            O => \N__23464\,
            I => \N__23461\
        );

    \I__5658\ : Odrv12
    port map (
            O => \N__23461\,
            I => \line_buffer.n546\
        );

    \I__5657\ : InMux
    port map (
            O => \N__23458\,
            I => \N__23455\
        );

    \I__5656\ : LocalMux
    port map (
            O => \N__23455\,
            I => \N__23452\
        );

    \I__5655\ : Span12Mux_h
    port map (
            O => \N__23452\,
            I => \N__23449\
        );

    \I__5654\ : Span12Mux_v
    port map (
            O => \N__23449\,
            I => \N__23446\
        );

    \I__5653\ : Odrv12
    port map (
            O => \N__23446\,
            I => \line_buffer.n538\
        );

    \I__5652\ : InMux
    port map (
            O => \N__23443\,
            I => \N__23440\
        );

    \I__5651\ : LocalMux
    port map (
            O => \N__23440\,
            I => \N__23437\
        );

    \I__5650\ : Odrv4
    port map (
            O => \N__23437\,
            I => \TX_DATA_3\
        );

    \I__5649\ : IoInMux
    port map (
            O => \N__23434\,
            I => \N__23431\
        );

    \I__5648\ : LocalMux
    port map (
            O => \N__23431\,
            I => \N__23428\
        );

    \I__5647\ : IoSpan4Mux
    port map (
            O => \N__23428\,
            I => \N__23425\
        );

    \I__5646\ : IoSpan4Mux
    port map (
            O => \N__23425\,
            I => \N__23421\
        );

    \I__5645\ : IoInMux
    port map (
            O => \N__23424\,
            I => \N__23418\
        );

    \I__5644\ : IoSpan4Mux
    port map (
            O => \N__23421\,
            I => \N__23412\
        );

    \I__5643\ : LocalMux
    port map (
            O => \N__23418\,
            I => \N__23412\
        );

    \I__5642\ : IoInMux
    port map (
            O => \N__23417\,
            I => \N__23409\
        );

    \I__5641\ : Span4Mux_s3_h
    port map (
            O => \N__23412\,
            I => \N__23406\
        );

    \I__5640\ : LocalMux
    port map (
            O => \N__23409\,
            I => \N__23403\
        );

    \I__5639\ : Span4Mux_h
    port map (
            O => \N__23406\,
            I => \N__23400\
        );

    \I__5638\ : IoSpan4Mux
    port map (
            O => \N__23403\,
            I => \N__23397\
        );

    \I__5637\ : Span4Mux_h
    port map (
            O => \N__23400\,
            I => \N__23394\
        );

    \I__5636\ : IoSpan4Mux
    port map (
            O => \N__23397\,
            I => \N__23391\
        );

    \I__5635\ : Span4Mux_h
    port map (
            O => \N__23394\,
            I => \N__23388\
        );

    \I__5634\ : Span4Mux_s2_v
    port map (
            O => \N__23391\,
            I => \N__23385\
        );

    \I__5633\ : Span4Mux_h
    port map (
            O => \N__23388\,
            I => \N__23382\
        );

    \I__5632\ : Sp12to4
    port map (
            O => \N__23385\,
            I => \N__23379\
        );

    \I__5631\ : Odrv4
    port map (
            O => \N__23382\,
            I => n1795
        );

    \I__5630\ : Odrv12
    port map (
            O => \N__23379\,
            I => n1795
        );

    \I__5629\ : InMux
    port map (
            O => \N__23374\,
            I => \N__23371\
        );

    \I__5628\ : LocalMux
    port map (
            O => \N__23371\,
            I => \N__23368\
        );

    \I__5627\ : Odrv12
    port map (
            O => \N__23368\,
            I => \TX_DATA_7\
        );

    \I__5626\ : IoInMux
    port map (
            O => \N__23365\,
            I => \N__23361\
        );

    \I__5625\ : IoInMux
    port map (
            O => \N__23364\,
            I => \N__23358\
        );

    \I__5624\ : LocalMux
    port map (
            O => \N__23361\,
            I => \N__23354\
        );

    \I__5623\ : LocalMux
    port map (
            O => \N__23358\,
            I => \N__23351\
        );

    \I__5622\ : IoInMux
    port map (
            O => \N__23357\,
            I => \N__23348\
        );

    \I__5621\ : Span4Mux_s2_h
    port map (
            O => \N__23354\,
            I => \N__23345\
        );

    \I__5620\ : Span4Mux_s2_v
    port map (
            O => \N__23351\,
            I => \N__23342\
        );

    \I__5619\ : LocalMux
    port map (
            O => \N__23348\,
            I => \N__23339\
        );

    \I__5618\ : Span4Mux_v
    port map (
            O => \N__23345\,
            I => \N__23336\
        );

    \I__5617\ : Span4Mux_h
    port map (
            O => \N__23342\,
            I => \N__23333\
        );

    \I__5616\ : IoSpan4Mux
    port map (
            O => \N__23339\,
            I => \N__23330\
        );

    \I__5615\ : Span4Mux_v
    port map (
            O => \N__23336\,
            I => \N__23327\
        );

    \I__5614\ : Span4Mux_v
    port map (
            O => \N__23333\,
            I => \N__23324\
        );

    \I__5613\ : Span4Mux_s3_v
    port map (
            O => \N__23330\,
            I => \N__23321\
        );

    \I__5612\ : Sp12to4
    port map (
            O => \N__23327\,
            I => \N__23318\
        );

    \I__5611\ : Span4Mux_v
    port map (
            O => \N__23324\,
            I => \N__23315\
        );

    \I__5610\ : Sp12to4
    port map (
            O => \N__23321\,
            I => \N__23312\
        );

    \I__5609\ : Span12Mux_h
    port map (
            O => \N__23318\,
            I => \N__23305\
        );

    \I__5608\ : Sp12to4
    port map (
            O => \N__23315\,
            I => \N__23305\
        );

    \I__5607\ : Span12Mux_s10_v
    port map (
            O => \N__23312\,
            I => \N__23305\
        );

    \I__5606\ : Odrv12
    port map (
            O => \N__23305\,
            I => \ADV_B_c\
        );

    \I__5605\ : ClkMux
    port map (
            O => \N__23302\,
            I => \N__23298\
        );

    \I__5604\ : ClkMux
    port map (
            O => \N__23301\,
            I => \N__23295\
        );

    \I__5603\ : LocalMux
    port map (
            O => \N__23298\,
            I => \N__23289\
        );

    \I__5602\ : LocalMux
    port map (
            O => \N__23295\,
            I => \N__23286\
        );

    \I__5601\ : ClkMux
    port map (
            O => \N__23294\,
            I => \N__23283\
        );

    \I__5600\ : ClkMux
    port map (
            O => \N__23293\,
            I => \N__23280\
        );

    \I__5599\ : ClkMux
    port map (
            O => \N__23292\,
            I => \N__23275\
        );

    \I__5598\ : Span4Mux_s2_v
    port map (
            O => \N__23289\,
            I => \N__23261\
        );

    \I__5597\ : Span4Mux_h
    port map (
            O => \N__23286\,
            I => \N__23261\
        );

    \I__5596\ : LocalMux
    port map (
            O => \N__23283\,
            I => \N__23261\
        );

    \I__5595\ : LocalMux
    port map (
            O => \N__23280\,
            I => \N__23258\
        );

    \I__5594\ : ClkMux
    port map (
            O => \N__23279\,
            I => \N__23255\
        );

    \I__5593\ : ClkMux
    port map (
            O => \N__23278\,
            I => \N__23252\
        );

    \I__5592\ : LocalMux
    port map (
            O => \N__23275\,
            I => \N__23248\
        );

    \I__5591\ : ClkMux
    port map (
            O => \N__23274\,
            I => \N__23245\
        );

    \I__5590\ : ClkMux
    port map (
            O => \N__23273\,
            I => \N__23242\
        );

    \I__5589\ : ClkMux
    port map (
            O => \N__23272\,
            I => \N__23239\
        );

    \I__5588\ : ClkMux
    port map (
            O => \N__23271\,
            I => \N__23236\
        );

    \I__5587\ : ClkMux
    port map (
            O => \N__23270\,
            I => \N__23232\
        );

    \I__5586\ : ClkMux
    port map (
            O => \N__23269\,
            I => \N__23229\
        );

    \I__5585\ : ClkMux
    port map (
            O => \N__23268\,
            I => \N__23226\
        );

    \I__5584\ : Span4Mux_v
    port map (
            O => \N__23261\,
            I => \N__23217\
        );

    \I__5583\ : Span4Mux_h
    port map (
            O => \N__23258\,
            I => \N__23217\
        );

    \I__5582\ : LocalMux
    port map (
            O => \N__23255\,
            I => \N__23217\
        );

    \I__5581\ : LocalMux
    port map (
            O => \N__23252\,
            I => \N__23214\
        );

    \I__5580\ : ClkMux
    port map (
            O => \N__23251\,
            I => \N__23211\
        );

    \I__5579\ : Span4Mux_h
    port map (
            O => \N__23248\,
            I => \N__23204\
        );

    \I__5578\ : LocalMux
    port map (
            O => \N__23245\,
            I => \N__23204\
        );

    \I__5577\ : LocalMux
    port map (
            O => \N__23242\,
            I => \N__23204\
        );

    \I__5576\ : LocalMux
    port map (
            O => \N__23239\,
            I => \N__23194\
        );

    \I__5575\ : LocalMux
    port map (
            O => \N__23236\,
            I => \N__23194\
        );

    \I__5574\ : ClkMux
    port map (
            O => \N__23235\,
            I => \N__23191\
        );

    \I__5573\ : LocalMux
    port map (
            O => \N__23232\,
            I => \N__23182\
        );

    \I__5572\ : LocalMux
    port map (
            O => \N__23229\,
            I => \N__23182\
        );

    \I__5571\ : LocalMux
    port map (
            O => \N__23226\,
            I => \N__23182\
        );

    \I__5570\ : ClkMux
    port map (
            O => \N__23225\,
            I => \N__23179\
        );

    \I__5569\ : ClkMux
    port map (
            O => \N__23224\,
            I => \N__23176\
        );

    \I__5568\ : Span4Mux_v
    port map (
            O => \N__23217\,
            I => \N__23167\
        );

    \I__5567\ : Span4Mux_h
    port map (
            O => \N__23214\,
            I => \N__23167\
        );

    \I__5566\ : LocalMux
    port map (
            O => \N__23211\,
            I => \N__23167\
        );

    \I__5565\ : Span4Mux_v
    port map (
            O => \N__23204\,
            I => \N__23164\
        );

    \I__5564\ : ClkMux
    port map (
            O => \N__23203\,
            I => \N__23161\
        );

    \I__5563\ : ClkMux
    port map (
            O => \N__23202\,
            I => \N__23156\
        );

    \I__5562\ : ClkMux
    port map (
            O => \N__23201\,
            I => \N__23153\
        );

    \I__5561\ : ClkMux
    port map (
            O => \N__23200\,
            I => \N__23148\
        );

    \I__5560\ : ClkMux
    port map (
            O => \N__23199\,
            I => \N__23145\
        );

    \I__5559\ : Span4Mux_s3_v
    port map (
            O => \N__23194\,
            I => \N__23138\
        );

    \I__5558\ : LocalMux
    port map (
            O => \N__23191\,
            I => \N__23138\
        );

    \I__5557\ : ClkMux
    port map (
            O => \N__23190\,
            I => \N__23135\
        );

    \I__5556\ : ClkMux
    port map (
            O => \N__23189\,
            I => \N__23131\
        );

    \I__5555\ : Span4Mux_v
    port map (
            O => \N__23182\,
            I => \N__23125\
        );

    \I__5554\ : LocalMux
    port map (
            O => \N__23179\,
            I => \N__23125\
        );

    \I__5553\ : LocalMux
    port map (
            O => \N__23176\,
            I => \N__23122\
        );

    \I__5552\ : ClkMux
    port map (
            O => \N__23175\,
            I => \N__23119\
        );

    \I__5551\ : ClkMux
    port map (
            O => \N__23174\,
            I => \N__23116\
        );

    \I__5550\ : Span4Mux_v
    port map (
            O => \N__23167\,
            I => \N__23113\
        );

    \I__5549\ : Span4Mux_v
    port map (
            O => \N__23164\,
            I => \N__23108\
        );

    \I__5548\ : LocalMux
    port map (
            O => \N__23161\,
            I => \N__23108\
        );

    \I__5547\ : ClkMux
    port map (
            O => \N__23160\,
            I => \N__23102\
        );

    \I__5546\ : ClkMux
    port map (
            O => \N__23159\,
            I => \N__23097\
        );

    \I__5545\ : LocalMux
    port map (
            O => \N__23156\,
            I => \N__23091\
        );

    \I__5544\ : LocalMux
    port map (
            O => \N__23153\,
            I => \N__23091\
        );

    \I__5543\ : ClkMux
    port map (
            O => \N__23152\,
            I => \N__23088\
        );

    \I__5542\ : ClkMux
    port map (
            O => \N__23151\,
            I => \N__23083\
        );

    \I__5541\ : LocalMux
    port map (
            O => \N__23148\,
            I => \N__23074\
        );

    \I__5540\ : LocalMux
    port map (
            O => \N__23145\,
            I => \N__23070\
        );

    \I__5539\ : ClkMux
    port map (
            O => \N__23144\,
            I => \N__23067\
        );

    \I__5538\ : ClkMux
    port map (
            O => \N__23143\,
            I => \N__23064\
        );

    \I__5537\ : Span4Mux_v
    port map (
            O => \N__23138\,
            I => \N__23059\
        );

    \I__5536\ : LocalMux
    port map (
            O => \N__23135\,
            I => \N__23059\
        );

    \I__5535\ : ClkMux
    port map (
            O => \N__23134\,
            I => \N__23056\
        );

    \I__5534\ : LocalMux
    port map (
            O => \N__23131\,
            I => \N__23052\
        );

    \I__5533\ : ClkMux
    port map (
            O => \N__23130\,
            I => \N__23049\
        );

    \I__5532\ : Span4Mux_v
    port map (
            O => \N__23125\,
            I => \N__23042\
        );

    \I__5531\ : Span4Mux_h
    port map (
            O => \N__23122\,
            I => \N__23042\
        );

    \I__5530\ : LocalMux
    port map (
            O => \N__23119\,
            I => \N__23042\
        );

    \I__5529\ : LocalMux
    port map (
            O => \N__23116\,
            I => \N__23039\
        );

    \I__5528\ : Span4Mux_h
    port map (
            O => \N__23113\,
            I => \N__23034\
        );

    \I__5527\ : Span4Mux_h
    port map (
            O => \N__23108\,
            I => \N__23034\
        );

    \I__5526\ : ClkMux
    port map (
            O => \N__23107\,
            I => \N__23031\
        );

    \I__5525\ : ClkMux
    port map (
            O => \N__23106\,
            I => \N__23028\
        );

    \I__5524\ : ClkMux
    port map (
            O => \N__23105\,
            I => \N__23023\
        );

    \I__5523\ : LocalMux
    port map (
            O => \N__23102\,
            I => \N__23020\
        );

    \I__5522\ : ClkMux
    port map (
            O => \N__23101\,
            I => \N__23017\
        );

    \I__5521\ : ClkMux
    port map (
            O => \N__23100\,
            I => \N__23014\
        );

    \I__5520\ : LocalMux
    port map (
            O => \N__23097\,
            I => \N__23011\
        );

    \I__5519\ : ClkMux
    port map (
            O => \N__23096\,
            I => \N__23008\
        );

    \I__5518\ : Span4Mux_h
    port map (
            O => \N__23091\,
            I => \N__23005\
        );

    \I__5517\ : LocalMux
    port map (
            O => \N__23088\,
            I => \N__23002\
        );

    \I__5516\ : ClkMux
    port map (
            O => \N__23087\,
            I => \N__22999\
        );

    \I__5515\ : ClkMux
    port map (
            O => \N__23086\,
            I => \N__22991\
        );

    \I__5514\ : LocalMux
    port map (
            O => \N__23083\,
            I => \N__22986\
        );

    \I__5513\ : ClkMux
    port map (
            O => \N__23082\,
            I => \N__22983\
        );

    \I__5512\ : ClkMux
    port map (
            O => \N__23081\,
            I => \N__22976\
        );

    \I__5511\ : ClkMux
    port map (
            O => \N__23080\,
            I => \N__22973\
        );

    \I__5510\ : ClkMux
    port map (
            O => \N__23079\,
            I => \N__22969\
        );

    \I__5509\ : ClkMux
    port map (
            O => \N__23078\,
            I => \N__22965\
        );

    \I__5508\ : ClkMux
    port map (
            O => \N__23077\,
            I => \N__22962\
        );

    \I__5507\ : Span4Mux_h
    port map (
            O => \N__23074\,
            I => \N__22958\
        );

    \I__5506\ : ClkMux
    port map (
            O => \N__23073\,
            I => \N__22955\
        );

    \I__5505\ : Span4Mux_v
    port map (
            O => \N__23070\,
            I => \N__22948\
        );

    \I__5504\ : LocalMux
    port map (
            O => \N__23067\,
            I => \N__22948\
        );

    \I__5503\ : LocalMux
    port map (
            O => \N__23064\,
            I => \N__22948\
        );

    \I__5502\ : Span4Mux_v
    port map (
            O => \N__23059\,
            I => \N__22942\
        );

    \I__5501\ : LocalMux
    port map (
            O => \N__23056\,
            I => \N__22942\
        );

    \I__5500\ : ClkMux
    port map (
            O => \N__23055\,
            I => \N__22939\
        );

    \I__5499\ : Span4Mux_h
    port map (
            O => \N__23052\,
            I => \N__22933\
        );

    \I__5498\ : LocalMux
    port map (
            O => \N__23049\,
            I => \N__22933\
        );

    \I__5497\ : Span4Mux_h
    port map (
            O => \N__23042\,
            I => \N__22923\
        );

    \I__5496\ : Span4Mux_h
    port map (
            O => \N__23039\,
            I => \N__22923\
        );

    \I__5495\ : Span4Mux_h
    port map (
            O => \N__23034\,
            I => \N__22923\
        );

    \I__5494\ : LocalMux
    port map (
            O => \N__23031\,
            I => \N__22923\
        );

    \I__5493\ : LocalMux
    port map (
            O => \N__23028\,
            I => \N__22920\
        );

    \I__5492\ : ClkMux
    port map (
            O => \N__23027\,
            I => \N__22917\
        );

    \I__5491\ : ClkMux
    port map (
            O => \N__23026\,
            I => \N__22914\
        );

    \I__5490\ : LocalMux
    port map (
            O => \N__23023\,
            I => \N__22909\
        );

    \I__5489\ : Span4Mux_h
    port map (
            O => \N__23020\,
            I => \N__22902\
        );

    \I__5488\ : LocalMux
    port map (
            O => \N__23017\,
            I => \N__22902\
        );

    \I__5487\ : LocalMux
    port map (
            O => \N__23014\,
            I => \N__22902\
        );

    \I__5486\ : Span4Mux_h
    port map (
            O => \N__23011\,
            I => \N__22897\
        );

    \I__5485\ : LocalMux
    port map (
            O => \N__23008\,
            I => \N__22897\
        );

    \I__5484\ : Span4Mux_v
    port map (
            O => \N__23005\,
            I => \N__22890\
        );

    \I__5483\ : Span4Mux_h
    port map (
            O => \N__23002\,
            I => \N__22890\
        );

    \I__5482\ : LocalMux
    port map (
            O => \N__22999\,
            I => \N__22890\
        );

    \I__5481\ : ClkMux
    port map (
            O => \N__22998\,
            I => \N__22887\
        );

    \I__5480\ : ClkMux
    port map (
            O => \N__22997\,
            I => \N__22884\
        );

    \I__5479\ : ClkMux
    port map (
            O => \N__22996\,
            I => \N__22879\
        );

    \I__5478\ : ClkMux
    port map (
            O => \N__22995\,
            I => \N__22876\
        );

    \I__5477\ : ClkMux
    port map (
            O => \N__22994\,
            I => \N__22873\
        );

    \I__5476\ : LocalMux
    port map (
            O => \N__22991\,
            I => \N__22869\
        );

    \I__5475\ : ClkMux
    port map (
            O => \N__22990\,
            I => \N__22866\
        );

    \I__5474\ : ClkMux
    port map (
            O => \N__22989\,
            I => \N__22863\
        );

    \I__5473\ : Span4Mux_h
    port map (
            O => \N__22986\,
            I => \N__22858\
        );

    \I__5472\ : LocalMux
    port map (
            O => \N__22983\,
            I => \N__22858\
        );

    \I__5471\ : ClkMux
    port map (
            O => \N__22982\,
            I => \N__22855\
        );

    \I__5470\ : ClkMux
    port map (
            O => \N__22981\,
            I => \N__22850\
        );

    \I__5469\ : ClkMux
    port map (
            O => \N__22980\,
            I => \N__22847\
        );

    \I__5468\ : ClkMux
    port map (
            O => \N__22979\,
            I => \N__22844\
        );

    \I__5467\ : LocalMux
    port map (
            O => \N__22976\,
            I => \N__22840\
        );

    \I__5466\ : LocalMux
    port map (
            O => \N__22973\,
            I => \N__22837\
        );

    \I__5465\ : ClkMux
    port map (
            O => \N__22972\,
            I => \N__22834\
        );

    \I__5464\ : LocalMux
    port map (
            O => \N__22969\,
            I => \N__22829\
        );

    \I__5463\ : ClkMux
    port map (
            O => \N__22968\,
            I => \N__22826\
        );

    \I__5462\ : LocalMux
    port map (
            O => \N__22965\,
            I => \N__22821\
        );

    \I__5461\ : LocalMux
    port map (
            O => \N__22962\,
            I => \N__22818\
        );

    \I__5460\ : ClkMux
    port map (
            O => \N__22961\,
            I => \N__22815\
        );

    \I__5459\ : Span4Mux_h
    port map (
            O => \N__22958\,
            I => \N__22810\
        );

    \I__5458\ : LocalMux
    port map (
            O => \N__22955\,
            I => \N__22810\
        );

    \I__5457\ : Span4Mux_h
    port map (
            O => \N__22948\,
            I => \N__22806\
        );

    \I__5456\ : ClkMux
    port map (
            O => \N__22947\,
            I => \N__22803\
        );

    \I__5455\ : Span4Mux_h
    port map (
            O => \N__22942\,
            I => \N__22800\
        );

    \I__5454\ : LocalMux
    port map (
            O => \N__22939\,
            I => \N__22797\
        );

    \I__5453\ : ClkMux
    port map (
            O => \N__22938\,
            I => \N__22794\
        );

    \I__5452\ : Span4Mux_h
    port map (
            O => \N__22933\,
            I => \N__22791\
        );

    \I__5451\ : ClkMux
    port map (
            O => \N__22932\,
            I => \N__22788\
        );

    \I__5450\ : Span4Mux_h
    port map (
            O => \N__22923\,
            I => \N__22785\
        );

    \I__5449\ : Span4Mux_h
    port map (
            O => \N__22920\,
            I => \N__22780\
        );

    \I__5448\ : LocalMux
    port map (
            O => \N__22917\,
            I => \N__22780\
        );

    \I__5447\ : LocalMux
    port map (
            O => \N__22914\,
            I => \N__22777\
        );

    \I__5446\ : ClkMux
    port map (
            O => \N__22913\,
            I => \N__22774\
        );

    \I__5445\ : ClkMux
    port map (
            O => \N__22912\,
            I => \N__22771\
        );

    \I__5444\ : Span4Mux_h
    port map (
            O => \N__22909\,
            I => \N__22765\
        );

    \I__5443\ : Span4Mux_h
    port map (
            O => \N__22902\,
            I => \N__22765\
        );

    \I__5442\ : Span4Mux_h
    port map (
            O => \N__22897\,
            I => \N__22758\
        );

    \I__5441\ : Span4Mux_h
    port map (
            O => \N__22890\,
            I => \N__22758\
        );

    \I__5440\ : LocalMux
    port map (
            O => \N__22887\,
            I => \N__22758\
        );

    \I__5439\ : LocalMux
    port map (
            O => \N__22884\,
            I => \N__22755\
        );

    \I__5438\ : ClkMux
    port map (
            O => \N__22883\,
            I => \N__22752\
        );

    \I__5437\ : ClkMux
    port map (
            O => \N__22882\,
            I => \N__22748\
        );

    \I__5436\ : LocalMux
    port map (
            O => \N__22879\,
            I => \N__22743\
        );

    \I__5435\ : LocalMux
    port map (
            O => \N__22876\,
            I => \N__22738\
        );

    \I__5434\ : LocalMux
    port map (
            O => \N__22873\,
            I => \N__22738\
        );

    \I__5433\ : ClkMux
    port map (
            O => \N__22872\,
            I => \N__22735\
        );

    \I__5432\ : Span4Mux_v
    port map (
            O => \N__22869\,
            I => \N__22728\
        );

    \I__5431\ : LocalMux
    port map (
            O => \N__22866\,
            I => \N__22728\
        );

    \I__5430\ : LocalMux
    port map (
            O => \N__22863\,
            I => \N__22728\
        );

    \I__5429\ : Span4Mux_h
    port map (
            O => \N__22858\,
            I => \N__22723\
        );

    \I__5428\ : LocalMux
    port map (
            O => \N__22855\,
            I => \N__22723\
        );

    \I__5427\ : ClkMux
    port map (
            O => \N__22854\,
            I => \N__22720\
        );

    \I__5426\ : ClkMux
    port map (
            O => \N__22853\,
            I => \N__22717\
        );

    \I__5425\ : LocalMux
    port map (
            O => \N__22850\,
            I => \N__22714\
        );

    \I__5424\ : LocalMux
    port map (
            O => \N__22847\,
            I => \N__22711\
        );

    \I__5423\ : LocalMux
    port map (
            O => \N__22844\,
            I => \N__22708\
        );

    \I__5422\ : ClkMux
    port map (
            O => \N__22843\,
            I => \N__22705\
        );

    \I__5421\ : Span4Mux_v
    port map (
            O => \N__22840\,
            I => \N__22698\
        );

    \I__5420\ : Span4Mux_h
    port map (
            O => \N__22837\,
            I => \N__22698\
        );

    \I__5419\ : LocalMux
    port map (
            O => \N__22834\,
            I => \N__22698\
        );

    \I__5418\ : ClkMux
    port map (
            O => \N__22833\,
            I => \N__22695\
        );

    \I__5417\ : ClkMux
    port map (
            O => \N__22832\,
            I => \N__22691\
        );

    \I__5416\ : Span4Mux_v
    port map (
            O => \N__22829\,
            I => \N__22685\
        );

    \I__5415\ : LocalMux
    port map (
            O => \N__22826\,
            I => \N__22685\
        );

    \I__5414\ : ClkMux
    port map (
            O => \N__22825\,
            I => \N__22682\
        );

    \I__5413\ : ClkMux
    port map (
            O => \N__22824\,
            I => \N__22679\
        );

    \I__5412\ : Span4Mux_h
    port map (
            O => \N__22821\,
            I => \N__22670\
        );

    \I__5411\ : Span4Mux_v
    port map (
            O => \N__22818\,
            I => \N__22670\
        );

    \I__5410\ : LocalMux
    port map (
            O => \N__22815\,
            I => \N__22670\
        );

    \I__5409\ : Span4Mux_h
    port map (
            O => \N__22810\,
            I => \N__22670\
        );

    \I__5408\ : ClkMux
    port map (
            O => \N__22809\,
            I => \N__22667\
        );

    \I__5407\ : Span4Mux_v
    port map (
            O => \N__22806\,
            I => \N__22662\
        );

    \I__5406\ : LocalMux
    port map (
            O => \N__22803\,
            I => \N__22662\
        );

    \I__5405\ : Span4Mux_v
    port map (
            O => \N__22800\,
            I => \N__22651\
        );

    \I__5404\ : Span4Mux_h
    port map (
            O => \N__22797\,
            I => \N__22651\
        );

    \I__5403\ : LocalMux
    port map (
            O => \N__22794\,
            I => \N__22651\
        );

    \I__5402\ : Span4Mux_h
    port map (
            O => \N__22791\,
            I => \N__22651\
        );

    \I__5401\ : LocalMux
    port map (
            O => \N__22788\,
            I => \N__22651\
        );

    \I__5400\ : Span4Mux_v
    port map (
            O => \N__22785\,
            I => \N__22646\
        );

    \I__5399\ : Span4Mux_v
    port map (
            O => \N__22780\,
            I => \N__22639\
        );

    \I__5398\ : Span4Mux_h
    port map (
            O => \N__22777\,
            I => \N__22639\
        );

    \I__5397\ : LocalMux
    port map (
            O => \N__22774\,
            I => \N__22639\
        );

    \I__5396\ : LocalMux
    port map (
            O => \N__22771\,
            I => \N__22636\
        );

    \I__5395\ : ClkMux
    port map (
            O => \N__22770\,
            I => \N__22633\
        );

    \I__5394\ : Span4Mux_v
    port map (
            O => \N__22765\,
            I => \N__22623\
        );

    \I__5393\ : Span4Mux_h
    port map (
            O => \N__22758\,
            I => \N__22623\
        );

    \I__5392\ : Span4Mux_v
    port map (
            O => \N__22755\,
            I => \N__22623\
        );

    \I__5391\ : LocalMux
    port map (
            O => \N__22752\,
            I => \N__22623\
        );

    \I__5390\ : ClkMux
    port map (
            O => \N__22751\,
            I => \N__22620\
        );

    \I__5389\ : LocalMux
    port map (
            O => \N__22748\,
            I => \N__22617\
        );

    \I__5388\ : ClkMux
    port map (
            O => \N__22747\,
            I => \N__22614\
        );

    \I__5387\ : ClkMux
    port map (
            O => \N__22746\,
            I => \N__22611\
        );

    \I__5386\ : Span4Mux_h
    port map (
            O => \N__22743\,
            I => \N__22603\
        );

    \I__5385\ : Span4Mux_h
    port map (
            O => \N__22738\,
            I => \N__22603\
        );

    \I__5384\ : LocalMux
    port map (
            O => \N__22735\,
            I => \N__22603\
        );

    \I__5383\ : Span4Mux_h
    port map (
            O => \N__22728\,
            I => \N__22594\
        );

    \I__5382\ : Span4Mux_v
    port map (
            O => \N__22723\,
            I => \N__22594\
        );

    \I__5381\ : LocalMux
    port map (
            O => \N__22720\,
            I => \N__22594\
        );

    \I__5380\ : LocalMux
    port map (
            O => \N__22717\,
            I => \N__22594\
        );

    \I__5379\ : Span4Mux_h
    port map (
            O => \N__22714\,
            I => \N__22585\
        );

    \I__5378\ : Span4Mux_v
    port map (
            O => \N__22711\,
            I => \N__22585\
        );

    \I__5377\ : Span4Mux_h
    port map (
            O => \N__22708\,
            I => \N__22585\
        );

    \I__5376\ : LocalMux
    port map (
            O => \N__22705\,
            I => \N__22585\
        );

    \I__5375\ : Span4Mux_v
    port map (
            O => \N__22698\,
            I => \N__22580\
        );

    \I__5374\ : LocalMux
    port map (
            O => \N__22695\,
            I => \N__22580\
        );

    \I__5373\ : ClkMux
    port map (
            O => \N__22694\,
            I => \N__22577\
        );

    \I__5372\ : LocalMux
    port map (
            O => \N__22691\,
            I => \N__22574\
        );

    \I__5371\ : ClkMux
    port map (
            O => \N__22690\,
            I => \N__22571\
        );

    \I__5370\ : Span4Mux_h
    port map (
            O => \N__22685\,
            I => \N__22566\
        );

    \I__5369\ : LocalMux
    port map (
            O => \N__22682\,
            I => \N__22566\
        );

    \I__5368\ : LocalMux
    port map (
            O => \N__22679\,
            I => \N__22559\
        );

    \I__5367\ : Span4Mux_h
    port map (
            O => \N__22670\,
            I => \N__22559\
        );

    \I__5366\ : LocalMux
    port map (
            O => \N__22667\,
            I => \N__22559\
        );

    \I__5365\ : Span4Mux_h
    port map (
            O => \N__22662\,
            I => \N__22552\
        );

    \I__5364\ : Span4Mux_h
    port map (
            O => \N__22651\,
            I => \N__22552\
        );

    \I__5363\ : ClkMux
    port map (
            O => \N__22650\,
            I => \N__22549\
        );

    \I__5362\ : ClkMux
    port map (
            O => \N__22649\,
            I => \N__22546\
        );

    \I__5361\ : Span4Mux_v
    port map (
            O => \N__22646\,
            I => \N__22542\
        );

    \I__5360\ : Span4Mux_v
    port map (
            O => \N__22639\,
            I => \N__22535\
        );

    \I__5359\ : Span4Mux_h
    port map (
            O => \N__22636\,
            I => \N__22535\
        );

    \I__5358\ : LocalMux
    port map (
            O => \N__22633\,
            I => \N__22535\
        );

    \I__5357\ : IoInMux
    port map (
            O => \N__22632\,
            I => \N__22532\
        );

    \I__5356\ : Span4Mux_v
    port map (
            O => \N__22623\,
            I => \N__22525\
        );

    \I__5355\ : LocalMux
    port map (
            O => \N__22620\,
            I => \N__22525\
        );

    \I__5354\ : Span4Mux_h
    port map (
            O => \N__22617\,
            I => \N__22520\
        );

    \I__5353\ : LocalMux
    port map (
            O => \N__22614\,
            I => \N__22520\
        );

    \I__5352\ : LocalMux
    port map (
            O => \N__22611\,
            I => \N__22517\
        );

    \I__5351\ : ClkMux
    port map (
            O => \N__22610\,
            I => \N__22514\
        );

    \I__5350\ : Span4Mux_v
    port map (
            O => \N__22603\,
            I => \N__22503\
        );

    \I__5349\ : Span4Mux_v
    port map (
            O => \N__22594\,
            I => \N__22503\
        );

    \I__5348\ : Span4Mux_h
    port map (
            O => \N__22585\,
            I => \N__22503\
        );

    \I__5347\ : Span4Mux_h
    port map (
            O => \N__22580\,
            I => \N__22503\
        );

    \I__5346\ : LocalMux
    port map (
            O => \N__22577\,
            I => \N__22503\
        );

    \I__5345\ : Span4Mux_h
    port map (
            O => \N__22574\,
            I => \N__22498\
        );

    \I__5344\ : LocalMux
    port map (
            O => \N__22571\,
            I => \N__22498\
        );

    \I__5343\ : Span4Mux_v
    port map (
            O => \N__22566\,
            I => \N__22492\
        );

    \I__5342\ : Span4Mux_h
    port map (
            O => \N__22559\,
            I => \N__22492\
        );

    \I__5341\ : ClkMux
    port map (
            O => \N__22558\,
            I => \N__22489\
        );

    \I__5340\ : ClkMux
    port map (
            O => \N__22557\,
            I => \N__22486\
        );

    \I__5339\ : Span4Mux_v
    port map (
            O => \N__22552\,
            I => \N__22483\
        );

    \I__5338\ : LocalMux
    port map (
            O => \N__22549\,
            I => \N__22480\
        );

    \I__5337\ : LocalMux
    port map (
            O => \N__22546\,
            I => \N__22477\
        );

    \I__5336\ : ClkMux
    port map (
            O => \N__22545\,
            I => \N__22474\
        );

    \I__5335\ : Span4Mux_v
    port map (
            O => \N__22542\,
            I => \N__22471\
        );

    \I__5334\ : Span4Mux_v
    port map (
            O => \N__22535\,
            I => \N__22468\
        );

    \I__5333\ : LocalMux
    port map (
            O => \N__22532\,
            I => \N__22465\
        );

    \I__5332\ : ClkMux
    port map (
            O => \N__22531\,
            I => \N__22462\
        );

    \I__5331\ : ClkMux
    port map (
            O => \N__22530\,
            I => \N__22458\
        );

    \I__5330\ : Span4Mux_h
    port map (
            O => \N__22525\,
            I => \N__22453\
        );

    \I__5329\ : Span4Mux_h
    port map (
            O => \N__22520\,
            I => \N__22453\
        );

    \I__5328\ : Span4Mux_h
    port map (
            O => \N__22517\,
            I => \N__22450\
        );

    \I__5327\ : LocalMux
    port map (
            O => \N__22514\,
            I => \N__22447\
        );

    \I__5326\ : Span4Mux_v
    port map (
            O => \N__22503\,
            I => \N__22442\
        );

    \I__5325\ : Span4Mux_h
    port map (
            O => \N__22498\,
            I => \N__22442\
        );

    \I__5324\ : ClkMux
    port map (
            O => \N__22497\,
            I => \N__22439\
        );

    \I__5323\ : Span4Mux_v
    port map (
            O => \N__22492\,
            I => \N__22434\
        );

    \I__5322\ : LocalMux
    port map (
            O => \N__22489\,
            I => \N__22434\
        );

    \I__5321\ : LocalMux
    port map (
            O => \N__22486\,
            I => \N__22431\
        );

    \I__5320\ : Span4Mux_v
    port map (
            O => \N__22483\,
            I => \N__22426\
        );

    \I__5319\ : Span4Mux_h
    port map (
            O => \N__22480\,
            I => \N__22426\
        );

    \I__5318\ : Span12Mux_h
    port map (
            O => \N__22477\,
            I => \N__22423\
        );

    \I__5317\ : LocalMux
    port map (
            O => \N__22474\,
            I => \N__22420\
        );

    \I__5316\ : Span4Mux_v
    port map (
            O => \N__22471\,
            I => \N__22415\
        );

    \I__5315\ : Span4Mux_h
    port map (
            O => \N__22468\,
            I => \N__22415\
        );

    \I__5314\ : Span4Mux_s1_v
    port map (
            O => \N__22465\,
            I => \N__22412\
        );

    \I__5313\ : LocalMux
    port map (
            O => \N__22462\,
            I => \N__22409\
        );

    \I__5312\ : ClkMux
    port map (
            O => \N__22461\,
            I => \N__22406\
        );

    \I__5311\ : LocalMux
    port map (
            O => \N__22458\,
            I => \N__22403\
        );

    \I__5310\ : Span4Mux_v
    port map (
            O => \N__22453\,
            I => \N__22400\
        );

    \I__5309\ : Span4Mux_v
    port map (
            O => \N__22450\,
            I => \N__22395\
        );

    \I__5308\ : Span4Mux_h
    port map (
            O => \N__22447\,
            I => \N__22395\
        );

    \I__5307\ : Span4Mux_v
    port map (
            O => \N__22442\,
            I => \N__22392\
        );

    \I__5306\ : LocalMux
    port map (
            O => \N__22439\,
            I => \N__22389\
        );

    \I__5305\ : Span4Mux_v
    port map (
            O => \N__22434\,
            I => \N__22384\
        );

    \I__5304\ : Span4Mux_h
    port map (
            O => \N__22431\,
            I => \N__22384\
        );

    \I__5303\ : Span4Mux_v
    port map (
            O => \N__22426\,
            I => \N__22381\
        );

    \I__5302\ : Span12Mux_v
    port map (
            O => \N__22423\,
            I => \N__22376\
        );

    \I__5301\ : Span12Mux_h
    port map (
            O => \N__22420\,
            I => \N__22376\
        );

    \I__5300\ : Sp12to4
    port map (
            O => \N__22415\,
            I => \N__22369\
        );

    \I__5299\ : Sp12to4
    port map (
            O => \N__22412\,
            I => \N__22369\
        );

    \I__5298\ : Sp12to4
    port map (
            O => \N__22409\,
            I => \N__22369\
        );

    \I__5297\ : LocalMux
    port map (
            O => \N__22406\,
            I => \N__22366\
        );

    \I__5296\ : Span12Mux_h
    port map (
            O => \N__22403\,
            I => \N__22363\
        );

    \I__5295\ : Span4Mux_v
    port map (
            O => \N__22400\,
            I => \N__22358\
        );

    \I__5294\ : Span4Mux_h
    port map (
            O => \N__22395\,
            I => \N__22358\
        );

    \I__5293\ : Span4Mux_v
    port map (
            O => \N__22392\,
            I => \N__22355\
        );

    \I__5292\ : Span12Mux_h
    port map (
            O => \N__22389\,
            I => \N__22350\
        );

    \I__5291\ : Sp12to4
    port map (
            O => \N__22384\,
            I => \N__22350\
        );

    \I__5290\ : Span4Mux_v
    port map (
            O => \N__22381\,
            I => \N__22347\
        );

    \I__5289\ : Span12Mux_v
    port map (
            O => \N__22376\,
            I => \N__22340\
        );

    \I__5288\ : Span12Mux_h
    port map (
            O => \N__22369\,
            I => \N__22340\
        );

    \I__5287\ : Span12Mux_h
    port map (
            O => \N__22366\,
            I => \N__22340\
        );

    \I__5286\ : Odrv12
    port map (
            O => \N__22363\,
            I => \ADV_CLK_c\
        );

    \I__5285\ : Odrv4
    port map (
            O => \N__22358\,
            I => \ADV_CLK_c\
        );

    \I__5284\ : Odrv4
    port map (
            O => \N__22355\,
            I => \ADV_CLK_c\
        );

    \I__5283\ : Odrv12
    port map (
            O => \N__22350\,
            I => \ADV_CLK_c\
        );

    \I__5282\ : Odrv4
    port map (
            O => \N__22347\,
            I => \ADV_CLK_c\
        );

    \I__5281\ : Odrv12
    port map (
            O => \N__22340\,
            I => \ADV_CLK_c\
        );

    \I__5280\ : SRMux
    port map (
            O => \N__22327\,
            I => \N__22323\
        );

    \I__5279\ : SRMux
    port map (
            O => \N__22326\,
            I => \N__22316\
        );

    \I__5278\ : LocalMux
    port map (
            O => \N__22323\,
            I => \N__22312\
        );

    \I__5277\ : SRMux
    port map (
            O => \N__22322\,
            I => \N__22309\
        );

    \I__5276\ : SRMux
    port map (
            O => \N__22321\,
            I => \N__22306\
        );

    \I__5275\ : SRMux
    port map (
            O => \N__22320\,
            I => \N__22303\
        );

    \I__5274\ : SRMux
    port map (
            O => \N__22319\,
            I => \N__22300\
        );

    \I__5273\ : LocalMux
    port map (
            O => \N__22316\,
            I => \N__22297\
        );

    \I__5272\ : SRMux
    port map (
            O => \N__22315\,
            I => \N__22294\
        );

    \I__5271\ : Span4Mux_v
    port map (
            O => \N__22312\,
            I => \N__22289\
        );

    \I__5270\ : LocalMux
    port map (
            O => \N__22309\,
            I => \N__22289\
        );

    \I__5269\ : LocalMux
    port map (
            O => \N__22306\,
            I => \N__22286\
        );

    \I__5268\ : LocalMux
    port map (
            O => \N__22303\,
            I => \N__22283\
        );

    \I__5267\ : LocalMux
    port map (
            O => \N__22300\,
            I => \N__22280\
        );

    \I__5266\ : Span4Mux_h
    port map (
            O => \N__22297\,
            I => \N__22275\
        );

    \I__5265\ : LocalMux
    port map (
            O => \N__22294\,
            I => \N__22275\
        );

    \I__5264\ : Span4Mux_h
    port map (
            O => \N__22289\,
            I => \N__22272\
        );

    \I__5263\ : Span4Mux_v
    port map (
            O => \N__22286\,
            I => \N__22267\
        );

    \I__5262\ : Span4Mux_v
    port map (
            O => \N__22283\,
            I => \N__22267\
        );

    \I__5261\ : Span4Mux_h
    port map (
            O => \N__22280\,
            I => \N__22264\
        );

    \I__5260\ : Span4Mux_h
    port map (
            O => \N__22275\,
            I => \N__22261\
        );

    \I__5259\ : Odrv4
    port map (
            O => \N__22272\,
            I => \transmit_module.n2354\
        );

    \I__5258\ : Odrv4
    port map (
            O => \N__22267\,
            I => \transmit_module.n2354\
        );

    \I__5257\ : Odrv4
    port map (
            O => \N__22264\,
            I => \transmit_module.n2354\
        );

    \I__5256\ : Odrv4
    port map (
            O => \N__22261\,
            I => \transmit_module.n2354\
        );

    \I__5255\ : InMux
    port map (
            O => \N__22252\,
            I => \N__22249\
        );

    \I__5254\ : LocalMux
    port map (
            O => \N__22249\,
            I => \N__22246\
        );

    \I__5253\ : Span4Mux_v
    port map (
            O => \N__22246\,
            I => \N__22243\
        );

    \I__5252\ : Span4Mux_h
    port map (
            O => \N__22243\,
            I => \N__22240\
        );

    \I__5251\ : Odrv4
    port map (
            O => \N__22240\,
            I => \line_buffer.n449\
        );

    \I__5250\ : CascadeMux
    port map (
            O => \N__22237\,
            I => \N__22228\
        );

    \I__5249\ : CascadeMux
    port map (
            O => \N__22236\,
            I => \N__22222\
        );

    \I__5248\ : CascadeMux
    port map (
            O => \N__22235\,
            I => \N__22219\
        );

    \I__5247\ : InMux
    port map (
            O => \N__22234\,
            I => \N__22212\
        );

    \I__5246\ : CascadeMux
    port map (
            O => \N__22233\,
            I => \N__22209\
        );

    \I__5245\ : CascadeMux
    port map (
            O => \N__22232\,
            I => \N__22206\
        );

    \I__5244\ : InMux
    port map (
            O => \N__22231\,
            I => \N__22203\
        );

    \I__5243\ : InMux
    port map (
            O => \N__22228\,
            I => \N__22200\
        );

    \I__5242\ : InMux
    port map (
            O => \N__22227\,
            I => \N__22190\
        );

    \I__5241\ : InMux
    port map (
            O => \N__22226\,
            I => \N__22190\
        );

    \I__5240\ : InMux
    port map (
            O => \N__22225\,
            I => \N__22190\
        );

    \I__5239\ : InMux
    port map (
            O => \N__22222\,
            I => \N__22190\
        );

    \I__5238\ : InMux
    port map (
            O => \N__22219\,
            I => \N__22187\
        );

    \I__5237\ : CascadeMux
    port map (
            O => \N__22218\,
            I => \N__22183\
        );

    \I__5236\ : CascadeMux
    port map (
            O => \N__22217\,
            I => \N__22180\
        );

    \I__5235\ : CascadeMux
    port map (
            O => \N__22216\,
            I => \N__22175\
        );

    \I__5234\ : InMux
    port map (
            O => \N__22215\,
            I => \N__22169\
        );

    \I__5233\ : LocalMux
    port map (
            O => \N__22212\,
            I => \N__22166\
        );

    \I__5232\ : InMux
    port map (
            O => \N__22209\,
            I => \N__22163\
        );

    \I__5231\ : InMux
    port map (
            O => \N__22206\,
            I => \N__22160\
        );

    \I__5230\ : LocalMux
    port map (
            O => \N__22203\,
            I => \N__22155\
        );

    \I__5229\ : LocalMux
    port map (
            O => \N__22200\,
            I => \N__22155\
        );

    \I__5228\ : InMux
    port map (
            O => \N__22199\,
            I => \N__22152\
        );

    \I__5227\ : LocalMux
    port map (
            O => \N__22190\,
            I => \N__22149\
        );

    \I__5226\ : LocalMux
    port map (
            O => \N__22187\,
            I => \N__22146\
        );

    \I__5225\ : InMux
    port map (
            O => \N__22186\,
            I => \N__22143\
        );

    \I__5224\ : InMux
    port map (
            O => \N__22183\,
            I => \N__22140\
        );

    \I__5223\ : InMux
    port map (
            O => \N__22180\,
            I => \N__22137\
        );

    \I__5222\ : InMux
    port map (
            O => \N__22179\,
            I => \N__22134\
        );

    \I__5221\ : InMux
    port map (
            O => \N__22178\,
            I => \N__22129\
        );

    \I__5220\ : InMux
    port map (
            O => \N__22175\,
            I => \N__22129\
        );

    \I__5219\ : CascadeMux
    port map (
            O => \N__22174\,
            I => \N__22126\
        );

    \I__5218\ : InMux
    port map (
            O => \N__22173\,
            I => \N__22119\
        );

    \I__5217\ : InMux
    port map (
            O => \N__22172\,
            I => \N__22116\
        );

    \I__5216\ : LocalMux
    port map (
            O => \N__22169\,
            I => \N__22107\
        );

    \I__5215\ : Span4Mux_v
    port map (
            O => \N__22166\,
            I => \N__22107\
        );

    \I__5214\ : LocalMux
    port map (
            O => \N__22163\,
            I => \N__22107\
        );

    \I__5213\ : LocalMux
    port map (
            O => \N__22160\,
            I => \N__22107\
        );

    \I__5212\ : Span4Mux_v
    port map (
            O => \N__22155\,
            I => \N__22104\
        );

    \I__5211\ : LocalMux
    port map (
            O => \N__22152\,
            I => \N__22097\
        );

    \I__5210\ : Span4Mux_v
    port map (
            O => \N__22149\,
            I => \N__22097\
        );

    \I__5209\ : Span4Mux_v
    port map (
            O => \N__22146\,
            I => \N__22097\
        );

    \I__5208\ : LocalMux
    port map (
            O => \N__22143\,
            I => \N__22092\
        );

    \I__5207\ : LocalMux
    port map (
            O => \N__22140\,
            I => \N__22092\
        );

    \I__5206\ : LocalMux
    port map (
            O => \N__22137\,
            I => \N__22089\
        );

    \I__5205\ : LocalMux
    port map (
            O => \N__22134\,
            I => \N__22086\
        );

    \I__5204\ : LocalMux
    port map (
            O => \N__22129\,
            I => \N__22083\
        );

    \I__5203\ : InMux
    port map (
            O => \N__22126\,
            I => \N__22080\
        );

    \I__5202\ : InMux
    port map (
            O => \N__22125\,
            I => \N__22077\
        );

    \I__5201\ : InMux
    port map (
            O => \N__22124\,
            I => \N__22074\
        );

    \I__5200\ : InMux
    port map (
            O => \N__22123\,
            I => \N__22069\
        );

    \I__5199\ : InMux
    port map (
            O => \N__22122\,
            I => \N__22069\
        );

    \I__5198\ : LocalMux
    port map (
            O => \N__22119\,
            I => \N__22066\
        );

    \I__5197\ : LocalMux
    port map (
            O => \N__22116\,
            I => \N__22057\
        );

    \I__5196\ : Span4Mux_v
    port map (
            O => \N__22107\,
            I => \N__22057\
        );

    \I__5195\ : Span4Mux_h
    port map (
            O => \N__22104\,
            I => \N__22057\
        );

    \I__5194\ : Span4Mux_h
    port map (
            O => \N__22097\,
            I => \N__22057\
        );

    \I__5193\ : Span4Mux_v
    port map (
            O => \N__22092\,
            I => \N__22052\
        );

    \I__5192\ : Span4Mux_v
    port map (
            O => \N__22089\,
            I => \N__22052\
        );

    \I__5191\ : Span4Mux_v
    port map (
            O => \N__22086\,
            I => \N__22045\
        );

    \I__5190\ : Span4Mux_v
    port map (
            O => \N__22083\,
            I => \N__22045\
        );

    \I__5189\ : LocalMux
    port map (
            O => \N__22080\,
            I => \N__22045\
        );

    \I__5188\ : LocalMux
    port map (
            O => \N__22077\,
            I => \TX_ADDR_12\
        );

    \I__5187\ : LocalMux
    port map (
            O => \N__22074\,
            I => \TX_ADDR_12\
        );

    \I__5186\ : LocalMux
    port map (
            O => \N__22069\,
            I => \TX_ADDR_12\
        );

    \I__5185\ : Odrv4
    port map (
            O => \N__22066\,
            I => \TX_ADDR_12\
        );

    \I__5184\ : Odrv4
    port map (
            O => \N__22057\,
            I => \TX_ADDR_12\
        );

    \I__5183\ : Odrv4
    port map (
            O => \N__22052\,
            I => \TX_ADDR_12\
        );

    \I__5182\ : Odrv4
    port map (
            O => \N__22045\,
            I => \TX_ADDR_12\
        );

    \I__5181\ : CascadeMux
    port map (
            O => \N__22030\,
            I => \N__22027\
        );

    \I__5180\ : InMux
    port map (
            O => \N__22027\,
            I => \N__22024\
        );

    \I__5179\ : LocalMux
    port map (
            O => \N__22024\,
            I => \N__22021\
        );

    \I__5178\ : Span12Mux_h
    port map (
            O => \N__22021\,
            I => \N__22018\
        );

    \I__5177\ : Span12Mux_v
    port map (
            O => \N__22018\,
            I => \N__22015\
        );

    \I__5176\ : Span12Mux_h
    port map (
            O => \N__22015\,
            I => \N__22012\
        );

    \I__5175\ : Odrv12
    port map (
            O => \N__22012\,
            I => \line_buffer.n441\
        );

    \I__5174\ : InMux
    port map (
            O => \N__22009\,
            I => \N__22006\
        );

    \I__5173\ : LocalMux
    port map (
            O => \N__22006\,
            I => \line_buffer.n3704\
        );

    \I__5172\ : InMux
    port map (
            O => \N__22003\,
            I => \N__22000\
        );

    \I__5171\ : LocalMux
    port map (
            O => \N__22000\,
            I => \line_buffer.n3707\
        );

    \I__5170\ : SRMux
    port map (
            O => \N__21997\,
            I => \N__21994\
        );

    \I__5169\ : LocalMux
    port map (
            O => \N__21994\,
            I => \N__21991\
        );

    \I__5168\ : Span4Mux_h
    port map (
            O => \N__21991\,
            I => \N__21986\
        );

    \I__5167\ : SRMux
    port map (
            O => \N__21990\,
            I => \N__21983\
        );

    \I__5166\ : SRMux
    port map (
            O => \N__21989\,
            I => \N__21980\
        );

    \I__5165\ : Span4Mux_v
    port map (
            O => \N__21986\,
            I => \N__21976\
        );

    \I__5164\ : LocalMux
    port map (
            O => \N__21983\,
            I => \N__21973\
        );

    \I__5163\ : LocalMux
    port map (
            O => \N__21980\,
            I => \N__21970\
        );

    \I__5162\ : SRMux
    port map (
            O => \N__21979\,
            I => \N__21967\
        );

    \I__5161\ : Span4Mux_v
    port map (
            O => \N__21976\,
            I => \N__21962\
        );

    \I__5160\ : Span4Mux_h
    port map (
            O => \N__21973\,
            I => \N__21962\
        );

    \I__5159\ : Span4Mux_h
    port map (
            O => \N__21970\,
            I => \N__21957\
        );

    \I__5158\ : LocalMux
    port map (
            O => \N__21967\,
            I => \N__21957\
        );

    \I__5157\ : Span4Mux_v
    port map (
            O => \N__21962\,
            I => \N__21951\
        );

    \I__5156\ : Span4Mux_h
    port map (
            O => \N__21957\,
            I => \N__21951\
        );

    \I__5155\ : SRMux
    port map (
            O => \N__21956\,
            I => \N__21948\
        );

    \I__5154\ : Span4Mux_v
    port map (
            O => \N__21951\,
            I => \N__21943\
        );

    \I__5153\ : LocalMux
    port map (
            O => \N__21948\,
            I => \N__21940\
        );

    \I__5152\ : SRMux
    port map (
            O => \N__21947\,
            I => \N__21937\
        );

    \I__5151\ : SRMux
    port map (
            O => \N__21946\,
            I => \N__21934\
        );

    \I__5150\ : Span4Mux_v
    port map (
            O => \N__21943\,
            I => \N__21926\
        );

    \I__5149\ : Span4Mux_h
    port map (
            O => \N__21940\,
            I => \N__21926\
        );

    \I__5148\ : LocalMux
    port map (
            O => \N__21937\,
            I => \N__21926\
        );

    \I__5147\ : LocalMux
    port map (
            O => \N__21934\,
            I => \N__21923\
        );

    \I__5146\ : SRMux
    port map (
            O => \N__21933\,
            I => \N__21920\
        );

    \I__5145\ : Span4Mux_v
    port map (
            O => \N__21926\,
            I => \N__21917\
        );

    \I__5144\ : Span4Mux_v
    port map (
            O => \N__21923\,
            I => \N__21914\
        );

    \I__5143\ : LocalMux
    port map (
            O => \N__21920\,
            I => \N__21911\
        );

    \I__5142\ : Odrv4
    port map (
            O => \N__21917\,
            I => \receive_module.n3793\
        );

    \I__5141\ : Odrv4
    port map (
            O => \N__21914\,
            I => \receive_module.n3793\
        );

    \I__5140\ : Odrv12
    port map (
            O => \N__21911\,
            I => \receive_module.n3793\
        );

    \I__5139\ : InMux
    port map (
            O => \N__21904\,
            I => \N__21901\
        );

    \I__5138\ : LocalMux
    port map (
            O => \N__21901\,
            I => \N__21898\
        );

    \I__5137\ : Span12Mux_v
    port map (
            O => \N__21898\,
            I => \N__21895\
        );

    \I__5136\ : Odrv12
    port map (
            O => \N__21895\,
            I => \line_buffer.n542\
        );

    \I__5135\ : InMux
    port map (
            O => \N__21892\,
            I => \N__21889\
        );

    \I__5134\ : LocalMux
    port map (
            O => \N__21889\,
            I => \N__21886\
        );

    \I__5133\ : Odrv12
    port map (
            O => \N__21886\,
            I => \line_buffer.n534\
        );

    \I__5132\ : InMux
    port map (
            O => \N__21883\,
            I => \N__21880\
        );

    \I__5131\ : LocalMux
    port map (
            O => \N__21880\,
            I => \N__21877\
        );

    \I__5130\ : Span4Mux_v
    port map (
            O => \N__21877\,
            I => \N__21874\
        );

    \I__5129\ : Span4Mux_h
    port map (
            O => \N__21874\,
            I => \N__21871\
        );

    \I__5128\ : Odrv4
    port map (
            O => \N__21871\,
            I => \line_buffer.n445\
        );

    \I__5127\ : CascadeMux
    port map (
            O => \N__21868\,
            I => \N__21865\
        );

    \I__5126\ : InMux
    port map (
            O => \N__21865\,
            I => \N__21862\
        );

    \I__5125\ : LocalMux
    port map (
            O => \N__21862\,
            I => \N__21859\
        );

    \I__5124\ : Span4Mux_v
    port map (
            O => \N__21859\,
            I => \N__21856\
        );

    \I__5123\ : Span4Mux_v
    port map (
            O => \N__21856\,
            I => \N__21853\
        );

    \I__5122\ : Sp12to4
    port map (
            O => \N__21853\,
            I => \N__21850\
        );

    \I__5121\ : Span12Mux_h
    port map (
            O => \N__21850\,
            I => \N__21847\
        );

    \I__5120\ : Odrv12
    port map (
            O => \N__21847\,
            I => \line_buffer.n437\
        );

    \I__5119\ : InMux
    port map (
            O => \N__21844\,
            I => \N__21841\
        );

    \I__5118\ : LocalMux
    port map (
            O => \N__21841\,
            I => \line_buffer.n3710\
        );

    \I__5117\ : InMux
    port map (
            O => \N__21838\,
            I => \N__21835\
        );

    \I__5116\ : LocalMux
    port map (
            O => \N__21835\,
            I => \N__21832\
        );

    \I__5115\ : Span4Mux_v
    port map (
            O => \N__21832\,
            I => \N__21829\
        );

    \I__5114\ : Span4Mux_h
    port map (
            O => \N__21829\,
            I => \N__21826\
        );

    \I__5113\ : Sp12to4
    port map (
            O => \N__21826\,
            I => \N__21823\
        );

    \I__5112\ : Odrv12
    port map (
            O => \N__21823\,
            I => \line_buffer.n566\
        );

    \I__5111\ : InMux
    port map (
            O => \N__21820\,
            I => \N__21817\
        );

    \I__5110\ : LocalMux
    port map (
            O => \N__21817\,
            I => \N__21814\
        );

    \I__5109\ : Sp12to4
    port map (
            O => \N__21814\,
            I => \N__21811\
        );

    \I__5108\ : Odrv12
    port map (
            O => \N__21811\,
            I => \line_buffer.n574\
        );

    \I__5107\ : InMux
    port map (
            O => \N__21808\,
            I => \N__21805\
        );

    \I__5106\ : LocalMux
    port map (
            O => \N__21805\,
            I => \N__21802\
        );

    \I__5105\ : Span4Mux_h
    port map (
            O => \N__21802\,
            I => \N__21799\
        );

    \I__5104\ : Span4Mux_v
    port map (
            O => \N__21799\,
            I => \N__21796\
        );

    \I__5103\ : Span4Mux_v
    port map (
            O => \N__21796\,
            I => \N__21793\
        );

    \I__5102\ : Odrv4
    port map (
            O => \N__21793\,
            I => \line_buffer.n502\
        );

    \I__5101\ : InMux
    port map (
            O => \N__21790\,
            I => \N__21787\
        );

    \I__5100\ : LocalMux
    port map (
            O => \N__21787\,
            I => \N__21784\
        );

    \I__5099\ : Span4Mux_v
    port map (
            O => \N__21784\,
            I => \N__21781\
        );

    \I__5098\ : Sp12to4
    port map (
            O => \N__21781\,
            I => \N__21778\
        );

    \I__5097\ : Span12Mux_v
    port map (
            O => \N__21778\,
            I => \N__21775\
        );

    \I__5096\ : Odrv12
    port map (
            O => \N__21775\,
            I => \line_buffer.n510\
        );

    \I__5095\ : CascadeMux
    port map (
            O => \N__21772\,
            I => \line_buffer.n3758_cascade_\
        );

    \I__5094\ : InMux
    port map (
            O => \N__21769\,
            I => \N__21766\
        );

    \I__5093\ : LocalMux
    port map (
            O => \N__21766\,
            I => \N__21763\
        );

    \I__5092\ : Span12Mux_v
    port map (
            O => \N__21763\,
            I => \N__21760\
        );

    \I__5091\ : Odrv12
    port map (
            O => \N__21760\,
            I => \line_buffer.n540\
        );

    \I__5090\ : InMux
    port map (
            O => \N__21757\,
            I => \N__21754\
        );

    \I__5089\ : LocalMux
    port map (
            O => \N__21754\,
            I => \N__21751\
        );

    \I__5088\ : Odrv12
    port map (
            O => \N__21751\,
            I => \line_buffer.n532\
        );

    \I__5087\ : InMux
    port map (
            O => \N__21748\,
            I => \N__21745\
        );

    \I__5086\ : LocalMux
    port map (
            O => \N__21745\,
            I => \N__21742\
        );

    \I__5085\ : Span4Mux_h
    port map (
            O => \N__21742\,
            I => \N__21739\
        );

    \I__5084\ : Sp12to4
    port map (
            O => \N__21739\,
            I => \N__21736\
        );

    \I__5083\ : Span12Mux_v
    port map (
            O => \N__21736\,
            I => \N__21733\
        );

    \I__5082\ : Odrv12
    port map (
            O => \N__21733\,
            I => \line_buffer.n435\
        );

    \I__5081\ : InMux
    port map (
            O => \N__21730\,
            I => \N__21727\
        );

    \I__5080\ : LocalMux
    port map (
            O => \N__21727\,
            I => \N__21724\
        );

    \I__5079\ : Span4Mux_v
    port map (
            O => \N__21724\,
            I => \N__21721\
        );

    \I__5078\ : Span4Mux_h
    port map (
            O => \N__21721\,
            I => \N__21718\
        );

    \I__5077\ : Odrv4
    port map (
            O => \N__21718\,
            I => \line_buffer.n443\
        );

    \I__5076\ : CascadeMux
    port map (
            O => \N__21715\,
            I => \line_buffer.n3740_cascade_\
        );

    \I__5075\ : InMux
    port map (
            O => \N__21712\,
            I => \N__21709\
        );

    \I__5074\ : LocalMux
    port map (
            O => \N__21709\,
            I => \line_buffer.n3743\
        );

    \I__5073\ : InMux
    port map (
            O => \N__21706\,
            I => \N__21703\
        );

    \I__5072\ : LocalMux
    port map (
            O => \N__21703\,
            I => \line_buffer.n3761\
        );

    \I__5071\ : InMux
    port map (
            O => \N__21700\,
            I => \N__21697\
        );

    \I__5070\ : LocalMux
    port map (
            O => \N__21697\,
            I => \line_buffer.n3713\
        );

    \I__5069\ : CascadeMux
    port map (
            O => \N__21694\,
            I => \N__21688\
        );

    \I__5068\ : InMux
    port map (
            O => \N__21693\,
            I => \N__21685\
        );

    \I__5067\ : InMux
    port map (
            O => \N__21692\,
            I => \N__21679\
        );

    \I__5066\ : InMux
    port map (
            O => \N__21691\,
            I => \N__21676\
        );

    \I__5065\ : InMux
    port map (
            O => \N__21688\,
            I => \N__21671\
        );

    \I__5064\ : LocalMux
    port map (
            O => \N__21685\,
            I => \N__21668\
        );

    \I__5063\ : InMux
    port map (
            O => \N__21684\,
            I => \N__21665\
        );

    \I__5062\ : InMux
    port map (
            O => \N__21683\,
            I => \N__21662\
        );

    \I__5061\ : CascadeMux
    port map (
            O => \N__21682\,
            I => \N__21658\
        );

    \I__5060\ : LocalMux
    port map (
            O => \N__21679\,
            I => \N__21653\
        );

    \I__5059\ : LocalMux
    port map (
            O => \N__21676\,
            I => \N__21653\
        );

    \I__5058\ : CascadeMux
    port map (
            O => \N__21675\,
            I => \N__21649\
        );

    \I__5057\ : CascadeMux
    port map (
            O => \N__21674\,
            I => \N__21646\
        );

    \I__5056\ : LocalMux
    port map (
            O => \N__21671\,
            I => \N__21641\
        );

    \I__5055\ : Span4Mux_v
    port map (
            O => \N__21668\,
            I => \N__21636\
        );

    \I__5054\ : LocalMux
    port map (
            O => \N__21665\,
            I => \N__21636\
        );

    \I__5053\ : LocalMux
    port map (
            O => \N__21662\,
            I => \N__21633\
        );

    \I__5052\ : InMux
    port map (
            O => \N__21661\,
            I => \N__21628\
        );

    \I__5051\ : InMux
    port map (
            O => \N__21658\,
            I => \N__21628\
        );

    \I__5050\ : Span4Mux_v
    port map (
            O => \N__21653\,
            I => \N__21625\
        );

    \I__5049\ : InMux
    port map (
            O => \N__21652\,
            I => \N__21622\
        );

    \I__5048\ : InMux
    port map (
            O => \N__21649\,
            I => \N__21617\
        );

    \I__5047\ : InMux
    port map (
            O => \N__21646\,
            I => \N__21617\
        );

    \I__5046\ : InMux
    port map (
            O => \N__21645\,
            I => \N__21614\
        );

    \I__5045\ : InMux
    port map (
            O => \N__21644\,
            I => \N__21611\
        );

    \I__5044\ : Span4Mux_v
    port map (
            O => \N__21641\,
            I => \N__21606\
        );

    \I__5043\ : Span4Mux_h
    port map (
            O => \N__21636\,
            I => \N__21606\
        );

    \I__5042\ : Span12Mux_h
    port map (
            O => \N__21633\,
            I => \N__21603\
        );

    \I__5041\ : LocalMux
    port map (
            O => \N__21628\,
            I => \N__21594\
        );

    \I__5040\ : Span4Mux_h
    port map (
            O => \N__21625\,
            I => \N__21594\
        );

    \I__5039\ : LocalMux
    port map (
            O => \N__21622\,
            I => \N__21594\
        );

    \I__5038\ : LocalMux
    port map (
            O => \N__21617\,
            I => \N__21594\
        );

    \I__5037\ : LocalMux
    port map (
            O => \N__21614\,
            I => \N__21591\
        );

    \I__5036\ : LocalMux
    port map (
            O => \N__21611\,
            I => \TX_ADDR_13\
        );

    \I__5035\ : Odrv4
    port map (
            O => \N__21606\,
            I => \TX_ADDR_13\
        );

    \I__5034\ : Odrv12
    port map (
            O => \N__21603\,
            I => \TX_ADDR_13\
        );

    \I__5033\ : Odrv4
    port map (
            O => \N__21594\,
            I => \TX_ADDR_13\
        );

    \I__5032\ : Odrv4
    port map (
            O => \N__21591\,
            I => \TX_ADDR_13\
        );

    \I__5031\ : InMux
    port map (
            O => \N__21580\,
            I => \N__21577\
        );

    \I__5030\ : LocalMux
    port map (
            O => \N__21577\,
            I => \N__21574\
        );

    \I__5029\ : Odrv12
    port map (
            O => \N__21574\,
            I => \line_buffer.n3767\
        );

    \I__5028\ : InMux
    port map (
            O => \N__21571\,
            I => \N__21568\
        );

    \I__5027\ : LocalMux
    port map (
            O => \N__21568\,
            I => \transmit_module.Y_DELTA_PATTERN_15\
        );

    \I__5026\ : InMux
    port map (
            O => \N__21565\,
            I => \N__21562\
        );

    \I__5025\ : LocalMux
    port map (
            O => \N__21562\,
            I => \transmit_module.Y_DELTA_PATTERN_14\
        );

    \I__5024\ : IoInMux
    port map (
            O => \N__21559\,
            I => \N__21555\
        );

    \I__5023\ : IoInMux
    port map (
            O => \N__21558\,
            I => \N__21552\
        );

    \I__5022\ : LocalMux
    port map (
            O => \N__21555\,
            I => \N__21549\
        );

    \I__5021\ : LocalMux
    port map (
            O => \N__21552\,
            I => \N__21546\
        );

    \I__5020\ : IoSpan4Mux
    port map (
            O => \N__21549\,
            I => \N__21542\
        );

    \I__5019\ : Span4Mux_s1_h
    port map (
            O => \N__21546\,
            I => \N__21539\
        );

    \I__5018\ : IoInMux
    port map (
            O => \N__21545\,
            I => \N__21536\
        );

    \I__5017\ : Span4Mux_s3_v
    port map (
            O => \N__21542\,
            I => \N__21533\
        );

    \I__5016\ : Span4Mux_h
    port map (
            O => \N__21539\,
            I => \N__21530\
        );

    \I__5015\ : LocalMux
    port map (
            O => \N__21536\,
            I => \N__21527\
        );

    \I__5014\ : Sp12to4
    port map (
            O => \N__21533\,
            I => \N__21522\
        );

    \I__5013\ : Sp12to4
    port map (
            O => \N__21530\,
            I => \N__21522\
        );

    \I__5012\ : Span4Mux_s0_v
    port map (
            O => \N__21527\,
            I => \N__21519\
        );

    \I__5011\ : Span12Mux_s11_v
    port map (
            O => \N__21522\,
            I => \N__21516\
        );

    \I__5010\ : Span4Mux_v
    port map (
            O => \N__21519\,
            I => \N__21513\
        );

    \I__5009\ : Span12Mux_h
    port map (
            O => \N__21516\,
            I => \N__21510\
        );

    \I__5008\ : Span4Mux_v
    port map (
            O => \N__21513\,
            I => \N__21507\
        );

    \I__5007\ : Odrv12
    port map (
            O => \N__21510\,
            I => n1797
        );

    \I__5006\ : Odrv4
    port map (
            O => \N__21507\,
            I => n1797
        );

    \I__5005\ : InMux
    port map (
            O => \N__21502\,
            I => \N__21499\
        );

    \I__5004\ : LocalMux
    port map (
            O => \N__21499\,
            I => \transmit_module.Y_DELTA_PATTERN_21\
        );

    \I__5003\ : InMux
    port map (
            O => \N__21496\,
            I => \N__21493\
        );

    \I__5002\ : LocalMux
    port map (
            O => \N__21493\,
            I => \transmit_module.Y_DELTA_PATTERN_20\
        );

    \I__5001\ : CEMux
    port map (
            O => \N__21490\,
            I => \N__21485\
        );

    \I__5000\ : CEMux
    port map (
            O => \N__21489\,
            I => \N__21479\
        );

    \I__4999\ : SRMux
    port map (
            O => \N__21488\,
            I => \N__21475\
        );

    \I__4998\ : LocalMux
    port map (
            O => \N__21485\,
            I => \N__21471\
        );

    \I__4997\ : CEMux
    port map (
            O => \N__21484\,
            I => \N__21468\
        );

    \I__4996\ : CEMux
    port map (
            O => \N__21483\,
            I => \N__21465\
        );

    \I__4995\ : CEMux
    port map (
            O => \N__21482\,
            I => \N__21462\
        );

    \I__4994\ : LocalMux
    port map (
            O => \N__21479\,
            I => \N__21454\
        );

    \I__4993\ : CEMux
    port map (
            O => \N__21478\,
            I => \N__21450\
        );

    \I__4992\ : LocalMux
    port map (
            O => \N__21475\,
            I => \N__21446\
        );

    \I__4991\ : SRMux
    port map (
            O => \N__21474\,
            I => \N__21443\
        );

    \I__4990\ : Span4Mux_v
    port map (
            O => \N__21471\,
            I => \N__21438\
        );

    \I__4989\ : LocalMux
    port map (
            O => \N__21468\,
            I => \N__21438\
        );

    \I__4988\ : LocalMux
    port map (
            O => \N__21465\,
            I => \N__21433\
        );

    \I__4987\ : LocalMux
    port map (
            O => \N__21462\,
            I => \N__21433\
        );

    \I__4986\ : CEMux
    port map (
            O => \N__21461\,
            I => \N__21430\
        );

    \I__4985\ : CEMux
    port map (
            O => \N__21460\,
            I => \N__21427\
        );

    \I__4984\ : CEMux
    port map (
            O => \N__21459\,
            I => \N__21424\
        );

    \I__4983\ : SRMux
    port map (
            O => \N__21458\,
            I => \N__21421\
        );

    \I__4982\ : SRMux
    port map (
            O => \N__21457\,
            I => \N__21418\
        );

    \I__4981\ : Span4Mux_v
    port map (
            O => \N__21454\,
            I => \N__21415\
        );

    \I__4980\ : CEMux
    port map (
            O => \N__21453\,
            I => \N__21412\
        );

    \I__4979\ : LocalMux
    port map (
            O => \N__21450\,
            I => \N__21409\
        );

    \I__4978\ : CEMux
    port map (
            O => \N__21449\,
            I => \N__21406\
        );

    \I__4977\ : Span4Mux_h
    port map (
            O => \N__21446\,
            I => \N__21403\
        );

    \I__4976\ : LocalMux
    port map (
            O => \N__21443\,
            I => \N__21400\
        );

    \I__4975\ : Span4Mux_v
    port map (
            O => \N__21438\,
            I => \N__21393\
        );

    \I__4974\ : Span4Mux_v
    port map (
            O => \N__21433\,
            I => \N__21393\
        );

    \I__4973\ : LocalMux
    port map (
            O => \N__21430\,
            I => \N__21393\
        );

    \I__4972\ : LocalMux
    port map (
            O => \N__21427\,
            I => \N__21390\
        );

    \I__4971\ : LocalMux
    port map (
            O => \N__21424\,
            I => \N__21387\
        );

    \I__4970\ : LocalMux
    port map (
            O => \N__21421\,
            I => \N__21382\
        );

    \I__4969\ : LocalMux
    port map (
            O => \N__21418\,
            I => \N__21382\
        );

    \I__4968\ : Sp12to4
    port map (
            O => \N__21415\,
            I => \N__21377\
        );

    \I__4967\ : LocalMux
    port map (
            O => \N__21412\,
            I => \N__21377\
        );

    \I__4966\ : Span4Mux_h
    port map (
            O => \N__21409\,
            I => \N__21368\
        );

    \I__4965\ : LocalMux
    port map (
            O => \N__21406\,
            I => \N__21368\
        );

    \I__4964\ : Span4Mux_h
    port map (
            O => \N__21403\,
            I => \N__21368\
        );

    \I__4963\ : Span4Mux_h
    port map (
            O => \N__21400\,
            I => \N__21368\
        );

    \I__4962\ : Span4Mux_h
    port map (
            O => \N__21393\,
            I => \N__21359\
        );

    \I__4961\ : Span4Mux_v
    port map (
            O => \N__21390\,
            I => \N__21359\
        );

    \I__4960\ : Span4Mux_v
    port map (
            O => \N__21387\,
            I => \N__21359\
        );

    \I__4959\ : Span4Mux_h
    port map (
            O => \N__21382\,
            I => \N__21359\
        );

    \I__4958\ : Odrv12
    port map (
            O => \N__21377\,
            I => \transmit_module.n3797\
        );

    \I__4957\ : Odrv4
    port map (
            O => \N__21368\,
            I => \transmit_module.n3797\
        );

    \I__4956\ : Odrv4
    port map (
            O => \N__21359\,
            I => \transmit_module.n3797\
        );

    \I__4955\ : IoInMux
    port map (
            O => \N__21352\,
            I => \N__21344\
        );

    \I__4954\ : SRMux
    port map (
            O => \N__21351\,
            I => \N__21341\
        );

    \I__4953\ : SRMux
    port map (
            O => \N__21350\,
            I => \N__21338\
        );

    \I__4952\ : SRMux
    port map (
            O => \N__21349\,
            I => \N__21335\
        );

    \I__4951\ : SRMux
    port map (
            O => \N__21348\,
            I => \N__21332\
        );

    \I__4950\ : SRMux
    port map (
            O => \N__21347\,
            I => \N__21326\
        );

    \I__4949\ : LocalMux
    port map (
            O => \N__21344\,
            I => \N__21321\
        );

    \I__4948\ : LocalMux
    port map (
            O => \N__21341\,
            I => \N__21315\
        );

    \I__4947\ : LocalMux
    port map (
            O => \N__21338\,
            I => \N__21308\
        );

    \I__4946\ : LocalMux
    port map (
            O => \N__21335\,
            I => \N__21308\
        );

    \I__4945\ : LocalMux
    port map (
            O => \N__21332\,
            I => \N__21308\
        );

    \I__4944\ : SRMux
    port map (
            O => \N__21331\,
            I => \N__21305\
        );

    \I__4943\ : SRMux
    port map (
            O => \N__21330\,
            I => \N__21297\
        );

    \I__4942\ : SRMux
    port map (
            O => \N__21329\,
            I => \N__21294\
        );

    \I__4941\ : LocalMux
    port map (
            O => \N__21326\,
            I => \N__21291\
        );

    \I__4940\ : SRMux
    port map (
            O => \N__21325\,
            I => \N__21288\
        );

    \I__4939\ : SRMux
    port map (
            O => \N__21324\,
            I => \N__21285\
        );

    \I__4938\ : IoSpan4Mux
    port map (
            O => \N__21321\,
            I => \N__21277\
        );

    \I__4937\ : SRMux
    port map (
            O => \N__21320\,
            I => \N__21272\
        );

    \I__4936\ : SRMux
    port map (
            O => \N__21319\,
            I => \N__21269\
        );

    \I__4935\ : CascadeMux
    port map (
            O => \N__21318\,
            I => \N__21262\
        );

    \I__4934\ : Span4Mux_h
    port map (
            O => \N__21315\,
            I => \N__21251\
        );

    \I__4933\ : Span4Mux_v
    port map (
            O => \N__21308\,
            I => \N__21251\
        );

    \I__4932\ : LocalMux
    port map (
            O => \N__21305\,
            I => \N__21251\
        );

    \I__4931\ : SRMux
    port map (
            O => \N__21304\,
            I => \N__21248\
        );

    \I__4930\ : SRMux
    port map (
            O => \N__21303\,
            I => \N__21245\
        );

    \I__4929\ : SRMux
    port map (
            O => \N__21302\,
            I => \N__21242\
        );

    \I__4928\ : SRMux
    port map (
            O => \N__21301\,
            I => \N__21239\
        );

    \I__4927\ : SRMux
    port map (
            O => \N__21300\,
            I => \N__21236\
        );

    \I__4926\ : LocalMux
    port map (
            O => \N__21297\,
            I => \N__21230\
        );

    \I__4925\ : LocalMux
    port map (
            O => \N__21294\,
            I => \N__21221\
        );

    \I__4924\ : Span4Mux_v
    port map (
            O => \N__21291\,
            I => \N__21221\
        );

    \I__4923\ : LocalMux
    port map (
            O => \N__21288\,
            I => \N__21221\
        );

    \I__4922\ : LocalMux
    port map (
            O => \N__21285\,
            I => \N__21221\
        );

    \I__4921\ : SRMux
    port map (
            O => \N__21284\,
            I => \N__21218\
        );

    \I__4920\ : SRMux
    port map (
            O => \N__21283\,
            I => \N__21215\
        );

    \I__4919\ : CascadeMux
    port map (
            O => \N__21282\,
            I => \N__21212\
        );

    \I__4918\ : CascadeMux
    port map (
            O => \N__21281\,
            I => \N__21209\
        );

    \I__4917\ : CascadeMux
    port map (
            O => \N__21280\,
            I => \N__21206\
        );

    \I__4916\ : Span4Mux_s3_h
    port map (
            O => \N__21277\,
            I => \N__21202\
        );

    \I__4915\ : SRMux
    port map (
            O => \N__21276\,
            I => \N__21199\
        );

    \I__4914\ : SRMux
    port map (
            O => \N__21275\,
            I => \N__21196\
        );

    \I__4913\ : LocalMux
    port map (
            O => \N__21272\,
            I => \N__21192\
        );

    \I__4912\ : LocalMux
    port map (
            O => \N__21269\,
            I => \N__21189\
        );

    \I__4911\ : CascadeMux
    port map (
            O => \N__21268\,
            I => \N__21186\
        );

    \I__4910\ : SRMux
    port map (
            O => \N__21267\,
            I => \N__21182\
        );

    \I__4909\ : SRMux
    port map (
            O => \N__21266\,
            I => \N__21179\
        );

    \I__4908\ : CascadeMux
    port map (
            O => \N__21265\,
            I => \N__21175\
        );

    \I__4907\ : InMux
    port map (
            O => \N__21262\,
            I => \N__21172\
        );

    \I__4906\ : SRMux
    port map (
            O => \N__21261\,
            I => \N__21168\
        );

    \I__4905\ : SRMux
    port map (
            O => \N__21260\,
            I => \N__21163\
        );

    \I__4904\ : CascadeMux
    port map (
            O => \N__21259\,
            I => \N__21160\
        );

    \I__4903\ : CascadeMux
    port map (
            O => \N__21258\,
            I => \N__21157\
        );

    \I__4902\ : Span4Mux_h
    port map (
            O => \N__21251\,
            I => \N__21152\
        );

    \I__4901\ : LocalMux
    port map (
            O => \N__21248\,
            I => \N__21152\
        );

    \I__4900\ : LocalMux
    port map (
            O => \N__21245\,
            I => \N__21145\
        );

    \I__4899\ : LocalMux
    port map (
            O => \N__21242\,
            I => \N__21145\
        );

    \I__4898\ : LocalMux
    port map (
            O => \N__21239\,
            I => \N__21145\
        );

    \I__4897\ : LocalMux
    port map (
            O => \N__21236\,
            I => \N__21142\
        );

    \I__4896\ : SRMux
    port map (
            O => \N__21235\,
            I => \N__21139\
        );

    \I__4895\ : CascadeMux
    port map (
            O => \N__21234\,
            I => \N__21135\
        );

    \I__4894\ : CascadeMux
    port map (
            O => \N__21233\,
            I => \N__21132\
        );

    \I__4893\ : Span4Mux_v
    port map (
            O => \N__21230\,
            I => \N__21124\
        );

    \I__4892\ : Span4Mux_v
    port map (
            O => \N__21221\,
            I => \N__21124\
        );

    \I__4891\ : LocalMux
    port map (
            O => \N__21218\,
            I => \N__21124\
        );

    \I__4890\ : LocalMux
    port map (
            O => \N__21215\,
            I => \N__21121\
        );

    \I__4889\ : InMux
    port map (
            O => \N__21212\,
            I => \N__21114\
        );

    \I__4888\ : InMux
    port map (
            O => \N__21209\,
            I => \N__21111\
        );

    \I__4887\ : InMux
    port map (
            O => \N__21206\,
            I => \N__21108\
        );

    \I__4886\ : CascadeMux
    port map (
            O => \N__21205\,
            I => \N__21105\
        );

    \I__4885\ : Span4Mux_h
    port map (
            O => \N__21202\,
            I => \N__21102\
        );

    \I__4884\ : LocalMux
    port map (
            O => \N__21199\,
            I => \N__21097\
        );

    \I__4883\ : LocalMux
    port map (
            O => \N__21196\,
            I => \N__21097\
        );

    \I__4882\ : SRMux
    port map (
            O => \N__21195\,
            I => \N__21094\
        );

    \I__4881\ : Span4Mux_h
    port map (
            O => \N__21192\,
            I => \N__21089\
        );

    \I__4880\ : Span4Mux_v
    port map (
            O => \N__21189\,
            I => \N__21089\
        );

    \I__4879\ : InMux
    port map (
            O => \N__21186\,
            I => \N__21086\
        );

    \I__4878\ : SRMux
    port map (
            O => \N__21185\,
            I => \N__21083\
        );

    \I__4877\ : LocalMux
    port map (
            O => \N__21182\,
            I => \N__21080\
        );

    \I__4876\ : LocalMux
    port map (
            O => \N__21179\,
            I => \N__21077\
        );

    \I__4875\ : InMux
    port map (
            O => \N__21178\,
            I => \N__21072\
        );

    \I__4874\ : InMux
    port map (
            O => \N__21175\,
            I => \N__21072\
        );

    \I__4873\ : LocalMux
    port map (
            O => \N__21172\,
            I => \N__21069\
        );

    \I__4872\ : SRMux
    port map (
            O => \N__21171\,
            I => \N__21066\
        );

    \I__4871\ : LocalMux
    port map (
            O => \N__21168\,
            I => \N__21063\
        );

    \I__4870\ : CascadeMux
    port map (
            O => \N__21167\,
            I => \N__21060\
        );

    \I__4869\ : CascadeMux
    port map (
            O => \N__21166\,
            I => \N__21056\
        );

    \I__4868\ : LocalMux
    port map (
            O => \N__21163\,
            I => \N__21045\
        );

    \I__4867\ : InMux
    port map (
            O => \N__21160\,
            I => \N__21040\
        );

    \I__4866\ : InMux
    port map (
            O => \N__21157\,
            I => \N__21040\
        );

    \I__4865\ : Span4Mux_v
    port map (
            O => \N__21152\,
            I => \N__21037\
        );

    \I__4864\ : Span4Mux_v
    port map (
            O => \N__21145\,
            I => \N__21030\
        );

    \I__4863\ : Span4Mux_h
    port map (
            O => \N__21142\,
            I => \N__21030\
        );

    \I__4862\ : LocalMux
    port map (
            O => \N__21139\,
            I => \N__21030\
        );

    \I__4861\ : CascadeMux
    port map (
            O => \N__21138\,
            I => \N__21027\
        );

    \I__4860\ : InMux
    port map (
            O => \N__21135\,
            I => \N__21020\
        );

    \I__4859\ : InMux
    port map (
            O => \N__21132\,
            I => \N__21020\
        );

    \I__4858\ : InMux
    port map (
            O => \N__21131\,
            I => \N__21020\
        );

    \I__4857\ : Span4Mux_h
    port map (
            O => \N__21124\,
            I => \N__21017\
        );

    \I__4856\ : Span4Mux_h
    port map (
            O => \N__21121\,
            I => \N__21014\
        );

    \I__4855\ : InMux
    port map (
            O => \N__21120\,
            I => \N__21009\
        );

    \I__4854\ : InMux
    port map (
            O => \N__21119\,
            I => \N__21009\
        );

    \I__4853\ : InMux
    port map (
            O => \N__21118\,
            I => \N__21006\
        );

    \I__4852\ : SRMux
    port map (
            O => \N__21117\,
            I => \N__20999\
        );

    \I__4851\ : LocalMux
    port map (
            O => \N__21114\,
            I => \N__20992\
        );

    \I__4850\ : LocalMux
    port map (
            O => \N__21111\,
            I => \N__20992\
        );

    \I__4849\ : LocalMux
    port map (
            O => \N__21108\,
            I => \N__20992\
        );

    \I__4848\ : InMux
    port map (
            O => \N__21105\,
            I => \N__20989\
        );

    \I__4847\ : Span4Mux_h
    port map (
            O => \N__21102\,
            I => \N__20982\
        );

    \I__4846\ : Span4Mux_v
    port map (
            O => \N__21097\,
            I => \N__20982\
        );

    \I__4845\ : LocalMux
    port map (
            O => \N__21094\,
            I => \N__20982\
        );

    \I__4844\ : Span4Mux_h
    port map (
            O => \N__21089\,
            I => \N__20977\
        );

    \I__4843\ : LocalMux
    port map (
            O => \N__21086\,
            I => \N__20977\
        );

    \I__4842\ : LocalMux
    port map (
            O => \N__21083\,
            I => \N__20974\
        );

    \I__4841\ : Span4Mux_v
    port map (
            O => \N__21080\,
            I => \N__20969\
        );

    \I__4840\ : Span4Mux_v
    port map (
            O => \N__21077\,
            I => \N__20969\
        );

    \I__4839\ : LocalMux
    port map (
            O => \N__21072\,
            I => \N__20966\
        );

    \I__4838\ : Span4Mux_v
    port map (
            O => \N__21069\,
            I => \N__20963\
        );

    \I__4837\ : LocalMux
    port map (
            O => \N__21066\,
            I => \N__20960\
        );

    \I__4836\ : Span4Mux_v
    port map (
            O => \N__21063\,
            I => \N__20957\
        );

    \I__4835\ : InMux
    port map (
            O => \N__21060\,
            I => \N__20952\
        );

    \I__4834\ : InMux
    port map (
            O => \N__21059\,
            I => \N__20952\
        );

    \I__4833\ : InMux
    port map (
            O => \N__21056\,
            I => \N__20945\
        );

    \I__4832\ : InMux
    port map (
            O => \N__21055\,
            I => \N__20945\
        );

    \I__4831\ : InMux
    port map (
            O => \N__21054\,
            I => \N__20945\
        );

    \I__4830\ : SRMux
    port map (
            O => \N__21053\,
            I => \N__20942\
        );

    \I__4829\ : InMux
    port map (
            O => \N__21052\,
            I => \N__20937\
        );

    \I__4828\ : InMux
    port map (
            O => \N__21051\,
            I => \N__20937\
        );

    \I__4827\ : SRMux
    port map (
            O => \N__21050\,
            I => \N__20934\
        );

    \I__4826\ : SRMux
    port map (
            O => \N__21049\,
            I => \N__20931\
        );

    \I__4825\ : SRMux
    port map (
            O => \N__21048\,
            I => \N__20928\
        );

    \I__4824\ : Span4Mux_v
    port map (
            O => \N__21045\,
            I => \N__20925\
        );

    \I__4823\ : LocalMux
    port map (
            O => \N__21040\,
            I => \N__20918\
        );

    \I__4822\ : Span4Mux_h
    port map (
            O => \N__21037\,
            I => \N__20918\
        );

    \I__4821\ : Span4Mux_h
    port map (
            O => \N__21030\,
            I => \N__20918\
        );

    \I__4820\ : InMux
    port map (
            O => \N__21027\,
            I => \N__20915\
        );

    \I__4819\ : LocalMux
    port map (
            O => \N__21020\,
            I => \N__20908\
        );

    \I__4818\ : Span4Mux_h
    port map (
            O => \N__21017\,
            I => \N__20908\
        );

    \I__4817\ : Span4Mux_v
    port map (
            O => \N__21014\,
            I => \N__20908\
        );

    \I__4816\ : LocalMux
    port map (
            O => \N__21009\,
            I => \N__20903\
        );

    \I__4815\ : LocalMux
    port map (
            O => \N__21006\,
            I => \N__20903\
        );

    \I__4814\ : InMux
    port map (
            O => \N__21005\,
            I => \N__20898\
        );

    \I__4813\ : InMux
    port map (
            O => \N__21004\,
            I => \N__20898\
        );

    \I__4812\ : InMux
    port map (
            O => \N__21003\,
            I => \N__20893\
        );

    \I__4811\ : InMux
    port map (
            O => \N__21002\,
            I => \N__20893\
        );

    \I__4810\ : LocalMux
    port map (
            O => \N__20999\,
            I => \N__20886\
        );

    \I__4809\ : Span12Mux_v
    port map (
            O => \N__20992\,
            I => \N__20886\
        );

    \I__4808\ : LocalMux
    port map (
            O => \N__20989\,
            I => \N__20886\
        );

    \I__4807\ : Span4Mux_v
    port map (
            O => \N__20982\,
            I => \N__20873\
        );

    \I__4806\ : Span4Mux_v
    port map (
            O => \N__20977\,
            I => \N__20873\
        );

    \I__4805\ : Span4Mux_h
    port map (
            O => \N__20974\,
            I => \N__20873\
        );

    \I__4804\ : Span4Mux_h
    port map (
            O => \N__20969\,
            I => \N__20873\
        );

    \I__4803\ : Span4Mux_v
    port map (
            O => \N__20966\,
            I => \N__20873\
        );

    \I__4802\ : Span4Mux_v
    port map (
            O => \N__20963\,
            I => \N__20873\
        );

    \I__4801\ : Sp12to4
    port map (
            O => \N__20960\,
            I => \N__20864\
        );

    \I__4800\ : Sp12to4
    port map (
            O => \N__20957\,
            I => \N__20864\
        );

    \I__4799\ : LocalMux
    port map (
            O => \N__20952\,
            I => \N__20864\
        );

    \I__4798\ : LocalMux
    port map (
            O => \N__20945\,
            I => \N__20864\
        );

    \I__4797\ : LocalMux
    port map (
            O => \N__20942\,
            I => \ADV_VSYNC_c\
        );

    \I__4796\ : LocalMux
    port map (
            O => \N__20937\,
            I => \ADV_VSYNC_c\
        );

    \I__4795\ : LocalMux
    port map (
            O => \N__20934\,
            I => \ADV_VSYNC_c\
        );

    \I__4794\ : LocalMux
    port map (
            O => \N__20931\,
            I => \ADV_VSYNC_c\
        );

    \I__4793\ : LocalMux
    port map (
            O => \N__20928\,
            I => \ADV_VSYNC_c\
        );

    \I__4792\ : Odrv4
    port map (
            O => \N__20925\,
            I => \ADV_VSYNC_c\
        );

    \I__4791\ : Odrv4
    port map (
            O => \N__20918\,
            I => \ADV_VSYNC_c\
        );

    \I__4790\ : LocalMux
    port map (
            O => \N__20915\,
            I => \ADV_VSYNC_c\
        );

    \I__4789\ : Odrv4
    port map (
            O => \N__20908\,
            I => \ADV_VSYNC_c\
        );

    \I__4788\ : Odrv12
    port map (
            O => \N__20903\,
            I => \ADV_VSYNC_c\
        );

    \I__4787\ : LocalMux
    port map (
            O => \N__20898\,
            I => \ADV_VSYNC_c\
        );

    \I__4786\ : LocalMux
    port map (
            O => \N__20893\,
            I => \ADV_VSYNC_c\
        );

    \I__4785\ : Odrv12
    port map (
            O => \N__20886\,
            I => \ADV_VSYNC_c\
        );

    \I__4784\ : Odrv4
    port map (
            O => \N__20873\,
            I => \ADV_VSYNC_c\
        );

    \I__4783\ : Odrv12
    port map (
            O => \N__20864\,
            I => \ADV_VSYNC_c\
        );

    \I__4782\ : InMux
    port map (
            O => \N__20833\,
            I => \N__20830\
        );

    \I__4781\ : LocalMux
    port map (
            O => \N__20830\,
            I => \N__20827\
        );

    \I__4780\ : Sp12to4
    port map (
            O => \N__20827\,
            I => \N__20824\
        );

    \I__4779\ : Span12Mux_v
    port map (
            O => \N__20824\,
            I => \N__20821\
        );

    \I__4778\ : Odrv12
    port map (
            O => \N__20821\,
            I => \line_buffer.n544\
        );

    \I__4777\ : InMux
    port map (
            O => \N__20818\,
            I => \N__20815\
        );

    \I__4776\ : LocalMux
    port map (
            O => \N__20815\,
            I => \N__20812\
        );

    \I__4775\ : Span4Mux_h
    port map (
            O => \N__20812\,
            I => \N__20809\
        );

    \I__4774\ : Span4Mux_h
    port map (
            O => \N__20809\,
            I => \N__20806\
        );

    \I__4773\ : Odrv4
    port map (
            O => \N__20806\,
            I => \line_buffer.n536\
        );

    \I__4772\ : InMux
    port map (
            O => \N__20803\,
            I => \N__20800\
        );

    \I__4771\ : LocalMux
    port map (
            O => \N__20800\,
            I => \N__20797\
        );

    \I__4770\ : Span4Mux_v
    port map (
            O => \N__20797\,
            I => \N__20794\
        );

    \I__4769\ : Odrv4
    port map (
            O => \N__20794\,
            I => \line_buffer.n3698\
        );

    \I__4768\ : InMux
    port map (
            O => \N__20791\,
            I => \N__20788\
        );

    \I__4767\ : LocalMux
    port map (
            O => \N__20788\,
            I => \N__20785\
        );

    \I__4766\ : Sp12to4
    port map (
            O => \N__20785\,
            I => \N__20782\
        );

    \I__4765\ : Span12Mux_v
    port map (
            O => \N__20782\,
            I => \N__20779\
        );

    \I__4764\ : Odrv12
    port map (
            O => \N__20779\,
            I => \line_buffer.n508\
        );

    \I__4763\ : CascadeMux
    port map (
            O => \N__20776\,
            I => \N__20773\
        );

    \I__4762\ : InMux
    port map (
            O => \N__20773\,
            I => \N__20770\
        );

    \I__4761\ : LocalMux
    port map (
            O => \N__20770\,
            I => \N__20767\
        );

    \I__4760\ : Span4Mux_h
    port map (
            O => \N__20767\,
            I => \N__20764\
        );

    \I__4759\ : Span4Mux_h
    port map (
            O => \N__20764\,
            I => \N__20761\
        );

    \I__4758\ : Span4Mux_v
    port map (
            O => \N__20761\,
            I => \N__20758\
        );

    \I__4757\ : Odrv4
    port map (
            O => \N__20758\,
            I => \line_buffer.n500\
        );

    \I__4756\ : CascadeMux
    port map (
            O => \N__20755\,
            I => \line_buffer.n3695_cascade_\
        );

    \I__4755\ : InMux
    port map (
            O => \N__20752\,
            I => \N__20749\
        );

    \I__4754\ : LocalMux
    port map (
            O => \N__20749\,
            I => \N__20746\
        );

    \I__4753\ : Span4Mux_v
    port map (
            O => \N__20746\,
            I => \N__20743\
        );

    \I__4752\ : Odrv4
    port map (
            O => \N__20743\,
            I => \TX_DATA_1\
        );

    \I__4751\ : InMux
    port map (
            O => \N__20740\,
            I => \N__20737\
        );

    \I__4750\ : LocalMux
    port map (
            O => \N__20737\,
            I => \N__20734\
        );

    \I__4749\ : Span4Mux_v
    port map (
            O => \N__20734\,
            I => \N__20731\
        );

    \I__4748\ : Sp12to4
    port map (
            O => \N__20731\,
            I => \N__20728\
        );

    \I__4747\ : Odrv12
    port map (
            O => \N__20728\,
            I => \line_buffer.n572\
        );

    \I__4746\ : InMux
    port map (
            O => \N__20725\,
            I => \N__20722\
        );

    \I__4745\ : LocalMux
    port map (
            O => \N__20722\,
            I => \N__20719\
        );

    \I__4744\ : Span4Mux_v
    port map (
            O => \N__20719\,
            I => \N__20716\
        );

    \I__4743\ : Sp12to4
    port map (
            O => \N__20716\,
            I => \N__20713\
        );

    \I__4742\ : Span12Mux_h
    port map (
            O => \N__20713\,
            I => \N__20710\
        );

    \I__4741\ : Span12Mux_v
    port map (
            O => \N__20710\,
            I => \N__20707\
        );

    \I__4740\ : Odrv12
    port map (
            O => \N__20707\,
            I => \line_buffer.n564\
        );

    \I__4739\ : InMux
    port map (
            O => \N__20704\,
            I => \N__20701\
        );

    \I__4738\ : LocalMux
    port map (
            O => \N__20701\,
            I => \line_buffer.n3692\
        );

    \I__4737\ : InMux
    port map (
            O => \N__20698\,
            I => \N__20680\
        );

    \I__4736\ : InMux
    port map (
            O => \N__20697\,
            I => \N__20680\
        );

    \I__4735\ : InMux
    port map (
            O => \N__20696\,
            I => \N__20680\
        );

    \I__4734\ : InMux
    port map (
            O => \N__20695\,
            I => \N__20680\
        );

    \I__4733\ : InMux
    port map (
            O => \N__20694\,
            I => \N__20680\
        );

    \I__4732\ : InMux
    port map (
            O => \N__20693\,
            I => \N__20680\
        );

    \I__4731\ : LocalMux
    port map (
            O => \N__20680\,
            I => \N__20675\
        );

    \I__4730\ : InMux
    port map (
            O => \N__20679\,
            I => \N__20669\
        );

    \I__4729\ : InMux
    port map (
            O => \N__20678\,
            I => \N__20666\
        );

    \I__4728\ : Span4Mux_v
    port map (
            O => \N__20675\,
            I => \N__20663\
        );

    \I__4727\ : InMux
    port map (
            O => \N__20674\,
            I => \N__20658\
        );

    \I__4726\ : InMux
    port map (
            O => \N__20673\,
            I => \N__20658\
        );

    \I__4725\ : InMux
    port map (
            O => \N__20672\,
            I => \N__20655\
        );

    \I__4724\ : LocalMux
    port map (
            O => \N__20669\,
            I => \N__20652\
        );

    \I__4723\ : LocalMux
    port map (
            O => \N__20666\,
            I => \N__20647\
        );

    \I__4722\ : Span4Mux_v
    port map (
            O => \N__20663\,
            I => \N__20647\
        );

    \I__4721\ : LocalMux
    port map (
            O => \N__20658\,
            I => \N__20644\
        );

    \I__4720\ : LocalMux
    port map (
            O => \N__20655\,
            I => \N__20637\
        );

    \I__4719\ : Span4Mux_h
    port map (
            O => \N__20652\,
            I => \N__20637\
        );

    \I__4718\ : Span4Mux_v
    port map (
            O => \N__20647\,
            I => \N__20637\
        );

    \I__4717\ : Span4Mux_v
    port map (
            O => \N__20644\,
            I => \N__20625\
        );

    \I__4716\ : Span4Mux_v
    port map (
            O => \N__20637\,
            I => \N__20622\
        );

    \I__4715\ : InMux
    port map (
            O => \N__20636\,
            I => \N__20617\
        );

    \I__4714\ : InMux
    port map (
            O => \N__20635\,
            I => \N__20617\
        );

    \I__4713\ : InMux
    port map (
            O => \N__20634\,
            I => \N__20614\
        );

    \I__4712\ : InMux
    port map (
            O => \N__20633\,
            I => \N__20611\
        );

    \I__4711\ : InMux
    port map (
            O => \N__20632\,
            I => \N__20608\
        );

    \I__4710\ : InMux
    port map (
            O => \N__20631\,
            I => \N__20599\
        );

    \I__4709\ : InMux
    port map (
            O => \N__20630\,
            I => \N__20599\
        );

    \I__4708\ : InMux
    port map (
            O => \N__20629\,
            I => \N__20599\
        );

    \I__4707\ : InMux
    port map (
            O => \N__20628\,
            I => \N__20599\
        );

    \I__4706\ : Odrv4
    port map (
            O => \N__20625\,
            I => \RX_WE\
        );

    \I__4705\ : Odrv4
    port map (
            O => \N__20622\,
            I => \RX_WE\
        );

    \I__4704\ : LocalMux
    port map (
            O => \N__20617\,
            I => \RX_WE\
        );

    \I__4703\ : LocalMux
    port map (
            O => \N__20614\,
            I => \RX_WE\
        );

    \I__4702\ : LocalMux
    port map (
            O => \N__20611\,
            I => \RX_WE\
        );

    \I__4701\ : LocalMux
    port map (
            O => \N__20608\,
            I => \RX_WE\
        );

    \I__4700\ : LocalMux
    port map (
            O => \N__20599\,
            I => \RX_WE\
        );

    \I__4699\ : InMux
    port map (
            O => \N__20584\,
            I => \N__20581\
        );

    \I__4698\ : LocalMux
    port map (
            O => \N__20581\,
            I => \N__20578\
        );

    \I__4697\ : Span4Mux_v
    port map (
            O => \N__20578\,
            I => \N__20575\
        );

    \I__4696\ : Span4Mux_v
    port map (
            O => \N__20575\,
            I => \N__20572\
        );

    \I__4695\ : Odrv4
    port map (
            O => \N__20572\,
            I => \receive_module.n133\
        );

    \I__4694\ : CascadeMux
    port map (
            O => \N__20569\,
            I => \N__20561\
        );

    \I__4693\ : CascadeMux
    port map (
            O => \N__20568\,
            I => \N__20558\
        );

    \I__4692\ : CascadeMux
    port map (
            O => \N__20567\,
            I => \N__20554\
        );

    \I__4691\ : CascadeMux
    port map (
            O => \N__20566\,
            I => \N__20551\
        );

    \I__4690\ : InMux
    port map (
            O => \N__20565\,
            I => \N__20546\
        );

    \I__4689\ : InMux
    port map (
            O => \N__20564\,
            I => \N__20546\
        );

    \I__4688\ : InMux
    port map (
            O => \N__20561\,
            I => \N__20537\
        );

    \I__4687\ : InMux
    port map (
            O => \N__20558\,
            I => \N__20537\
        );

    \I__4686\ : InMux
    port map (
            O => \N__20557\,
            I => \N__20537\
        );

    \I__4685\ : InMux
    port map (
            O => \N__20554\,
            I => \N__20537\
        );

    \I__4684\ : InMux
    port map (
            O => \N__20551\,
            I => \N__20531\
        );

    \I__4683\ : LocalMux
    port map (
            O => \N__20546\,
            I => \N__20528\
        );

    \I__4682\ : LocalMux
    port map (
            O => \N__20537\,
            I => \N__20525\
        );

    \I__4681\ : CascadeMux
    port map (
            O => \N__20536\,
            I => \N__20522\
        );

    \I__4680\ : CascadeMux
    port map (
            O => \N__20535\,
            I => \N__20518\
        );

    \I__4679\ : InMux
    port map (
            O => \N__20534\,
            I => \N__20515\
        );

    \I__4678\ : LocalMux
    port map (
            O => \N__20531\,
            I => \N__20512\
        );

    \I__4677\ : Span4Mux_v
    port map (
            O => \N__20528\,
            I => \N__20507\
        );

    \I__4676\ : Span4Mux_v
    port map (
            O => \N__20525\,
            I => \N__20507\
        );

    \I__4675\ : InMux
    port map (
            O => \N__20522\,
            I => \N__20504\
        );

    \I__4674\ : InMux
    port map (
            O => \N__20521\,
            I => \N__20498\
        );

    \I__4673\ : InMux
    port map (
            O => \N__20518\,
            I => \N__20498\
        );

    \I__4672\ : LocalMux
    port map (
            O => \N__20515\,
            I => \N__20495\
        );

    \I__4671\ : Span4Mux_v
    port map (
            O => \N__20512\,
            I => \N__20492\
        );

    \I__4670\ : Span4Mux_v
    port map (
            O => \N__20507\,
            I => \N__20487\
        );

    \I__4669\ : LocalMux
    port map (
            O => \N__20504\,
            I => \N__20487\
        );

    \I__4668\ : CascadeMux
    port map (
            O => \N__20503\,
            I => \N__20484\
        );

    \I__4667\ : LocalMux
    port map (
            O => \N__20498\,
            I => \N__20480\
        );

    \I__4666\ : Span4Mux_v
    port map (
            O => \N__20495\,
            I => \N__20477\
        );

    \I__4665\ : Span4Mux_h
    port map (
            O => \N__20492\,
            I => \N__20472\
        );

    \I__4664\ : Span4Mux_v
    port map (
            O => \N__20487\,
            I => \N__20472\
        );

    \I__4663\ : InMux
    port map (
            O => \N__20484\,
            I => \N__20469\
        );

    \I__4662\ : InMux
    port map (
            O => \N__20483\,
            I => \N__20466\
        );

    \I__4661\ : Span4Mux_h
    port map (
            O => \N__20480\,
            I => \N__20459\
        );

    \I__4660\ : Sp12to4
    port map (
            O => \N__20477\,
            I => \N__20456\
        );

    \I__4659\ : Sp12to4
    port map (
            O => \N__20472\,
            I => \N__20449\
        );

    \I__4658\ : LocalMux
    port map (
            O => \N__20469\,
            I => \N__20449\
        );

    \I__4657\ : LocalMux
    port map (
            O => \N__20466\,
            I => \N__20449\
        );

    \I__4656\ : InMux
    port map (
            O => \N__20465\,
            I => \N__20446\
        );

    \I__4655\ : InMux
    port map (
            O => \N__20464\,
            I => \N__20439\
        );

    \I__4654\ : InMux
    port map (
            O => \N__20463\,
            I => \N__20439\
        );

    \I__4653\ : InMux
    port map (
            O => \N__20462\,
            I => \N__20439\
        );

    \I__4652\ : Span4Mux_v
    port map (
            O => \N__20459\,
            I => \N__20436\
        );

    \I__4651\ : Span12Mux_h
    port map (
            O => \N__20456\,
            I => \N__20427\
        );

    \I__4650\ : Span12Mux_v
    port map (
            O => \N__20449\,
            I => \N__20427\
        );

    \I__4649\ : LocalMux
    port map (
            O => \N__20446\,
            I => \N__20427\
        );

    \I__4648\ : LocalMux
    port map (
            O => \N__20439\,
            I => \N__20427\
        );

    \I__4647\ : Odrv4
    port map (
            O => \N__20436\,
            I => \TVP_VSYNC_c\
        );

    \I__4646\ : Odrv12
    port map (
            O => \N__20427\,
            I => \TVP_VSYNC_c\
        );

    \I__4645\ : CascadeMux
    port map (
            O => \N__20422\,
            I => \N__20418\
        );

    \I__4644\ : CascadeMux
    port map (
            O => \N__20421\,
            I => \N__20415\
        );

    \I__4643\ : CascadeBuf
    port map (
            O => \N__20418\,
            I => \N__20412\
        );

    \I__4642\ : CascadeBuf
    port map (
            O => \N__20415\,
            I => \N__20409\
        );

    \I__4641\ : CascadeMux
    port map (
            O => \N__20412\,
            I => \N__20406\
        );

    \I__4640\ : CascadeMux
    port map (
            O => \N__20409\,
            I => \N__20403\
        );

    \I__4639\ : CascadeBuf
    port map (
            O => \N__20406\,
            I => \N__20400\
        );

    \I__4638\ : CascadeBuf
    port map (
            O => \N__20403\,
            I => \N__20397\
        );

    \I__4637\ : CascadeMux
    port map (
            O => \N__20400\,
            I => \N__20394\
        );

    \I__4636\ : CascadeMux
    port map (
            O => \N__20397\,
            I => \N__20391\
        );

    \I__4635\ : CascadeBuf
    port map (
            O => \N__20394\,
            I => \N__20388\
        );

    \I__4634\ : CascadeBuf
    port map (
            O => \N__20391\,
            I => \N__20385\
        );

    \I__4633\ : CascadeMux
    port map (
            O => \N__20388\,
            I => \N__20382\
        );

    \I__4632\ : CascadeMux
    port map (
            O => \N__20385\,
            I => \N__20379\
        );

    \I__4631\ : CascadeBuf
    port map (
            O => \N__20382\,
            I => \N__20376\
        );

    \I__4630\ : CascadeBuf
    port map (
            O => \N__20379\,
            I => \N__20373\
        );

    \I__4629\ : CascadeMux
    port map (
            O => \N__20376\,
            I => \N__20370\
        );

    \I__4628\ : CascadeMux
    port map (
            O => \N__20373\,
            I => \N__20367\
        );

    \I__4627\ : CascadeBuf
    port map (
            O => \N__20370\,
            I => \N__20364\
        );

    \I__4626\ : CascadeBuf
    port map (
            O => \N__20367\,
            I => \N__20361\
        );

    \I__4625\ : CascadeMux
    port map (
            O => \N__20364\,
            I => \N__20358\
        );

    \I__4624\ : CascadeMux
    port map (
            O => \N__20361\,
            I => \N__20355\
        );

    \I__4623\ : CascadeBuf
    port map (
            O => \N__20358\,
            I => \N__20352\
        );

    \I__4622\ : CascadeBuf
    port map (
            O => \N__20355\,
            I => \N__20349\
        );

    \I__4621\ : CascadeMux
    port map (
            O => \N__20352\,
            I => \N__20346\
        );

    \I__4620\ : CascadeMux
    port map (
            O => \N__20349\,
            I => \N__20343\
        );

    \I__4619\ : CascadeBuf
    port map (
            O => \N__20346\,
            I => \N__20340\
        );

    \I__4618\ : CascadeBuf
    port map (
            O => \N__20343\,
            I => \N__20337\
        );

    \I__4617\ : CascadeMux
    port map (
            O => \N__20340\,
            I => \N__20334\
        );

    \I__4616\ : CascadeMux
    port map (
            O => \N__20337\,
            I => \N__20331\
        );

    \I__4615\ : CascadeBuf
    port map (
            O => \N__20334\,
            I => \N__20328\
        );

    \I__4614\ : CascadeBuf
    port map (
            O => \N__20331\,
            I => \N__20325\
        );

    \I__4613\ : CascadeMux
    port map (
            O => \N__20328\,
            I => \N__20322\
        );

    \I__4612\ : CascadeMux
    port map (
            O => \N__20325\,
            I => \N__20319\
        );

    \I__4611\ : CascadeBuf
    port map (
            O => \N__20322\,
            I => \N__20316\
        );

    \I__4610\ : CascadeBuf
    port map (
            O => \N__20319\,
            I => \N__20313\
        );

    \I__4609\ : CascadeMux
    port map (
            O => \N__20316\,
            I => \N__20310\
        );

    \I__4608\ : CascadeMux
    port map (
            O => \N__20313\,
            I => \N__20307\
        );

    \I__4607\ : CascadeBuf
    port map (
            O => \N__20310\,
            I => \N__20304\
        );

    \I__4606\ : CascadeBuf
    port map (
            O => \N__20307\,
            I => \N__20301\
        );

    \I__4605\ : CascadeMux
    port map (
            O => \N__20304\,
            I => \N__20298\
        );

    \I__4604\ : CascadeMux
    port map (
            O => \N__20301\,
            I => \N__20295\
        );

    \I__4603\ : CascadeBuf
    port map (
            O => \N__20298\,
            I => \N__20292\
        );

    \I__4602\ : CascadeBuf
    port map (
            O => \N__20295\,
            I => \N__20289\
        );

    \I__4601\ : CascadeMux
    port map (
            O => \N__20292\,
            I => \N__20286\
        );

    \I__4600\ : CascadeMux
    port map (
            O => \N__20289\,
            I => \N__20283\
        );

    \I__4599\ : CascadeBuf
    port map (
            O => \N__20286\,
            I => \N__20280\
        );

    \I__4598\ : CascadeBuf
    port map (
            O => \N__20283\,
            I => \N__20277\
        );

    \I__4597\ : CascadeMux
    port map (
            O => \N__20280\,
            I => \N__20274\
        );

    \I__4596\ : CascadeMux
    port map (
            O => \N__20277\,
            I => \N__20271\
        );

    \I__4595\ : CascadeBuf
    port map (
            O => \N__20274\,
            I => \N__20268\
        );

    \I__4594\ : CascadeBuf
    port map (
            O => \N__20271\,
            I => \N__20265\
        );

    \I__4593\ : CascadeMux
    port map (
            O => \N__20268\,
            I => \N__20262\
        );

    \I__4592\ : CascadeMux
    port map (
            O => \N__20265\,
            I => \N__20259\
        );

    \I__4591\ : CascadeBuf
    port map (
            O => \N__20262\,
            I => \N__20256\
        );

    \I__4590\ : CascadeBuf
    port map (
            O => \N__20259\,
            I => \N__20253\
        );

    \I__4589\ : CascadeMux
    port map (
            O => \N__20256\,
            I => \N__20250\
        );

    \I__4588\ : CascadeMux
    port map (
            O => \N__20253\,
            I => \N__20247\
        );

    \I__4587\ : CascadeBuf
    port map (
            O => \N__20250\,
            I => \N__20244\
        );

    \I__4586\ : CascadeBuf
    port map (
            O => \N__20247\,
            I => \N__20241\
        );

    \I__4585\ : CascadeMux
    port map (
            O => \N__20244\,
            I => \N__20237\
        );

    \I__4584\ : CascadeMux
    port map (
            O => \N__20241\,
            I => \N__20234\
        );

    \I__4583\ : CascadeMux
    port map (
            O => \N__20240\,
            I => \N__20231\
        );

    \I__4582\ : InMux
    port map (
            O => \N__20237\,
            I => \N__20228\
        );

    \I__4581\ : InMux
    port map (
            O => \N__20234\,
            I => \N__20225\
        );

    \I__4580\ : InMux
    port map (
            O => \N__20231\,
            I => \N__20222\
        );

    \I__4579\ : LocalMux
    port map (
            O => \N__20228\,
            I => \N__20219\
        );

    \I__4578\ : LocalMux
    port map (
            O => \N__20225\,
            I => \N__20216\
        );

    \I__4577\ : LocalMux
    port map (
            O => \N__20222\,
            I => \N__20213\
        );

    \I__4576\ : Span4Mux_h
    port map (
            O => \N__20219\,
            I => \N__20210\
        );

    \I__4575\ : Span12Mux_s1_v
    port map (
            O => \N__20216\,
            I => \N__20206\
        );

    \I__4574\ : Sp12to4
    port map (
            O => \N__20213\,
            I => \N__20203\
        );

    \I__4573\ : Sp12to4
    port map (
            O => \N__20210\,
            I => \N__20200\
        );

    \I__4572\ : InMux
    port map (
            O => \N__20209\,
            I => \N__20197\
        );

    \I__4571\ : Span12Mux_v
    port map (
            O => \N__20206\,
            I => \N__20194\
        );

    \I__4570\ : Span12Mux_v
    port map (
            O => \N__20203\,
            I => \N__20189\
        );

    \I__4569\ : Span12Mux_v
    port map (
            O => \N__20200\,
            I => \N__20189\
        );

    \I__4568\ : LocalMux
    port map (
            O => \N__20197\,
            I => \RX_ADDR_3\
        );

    \I__4567\ : Odrv12
    port map (
            O => \N__20194\,
            I => \RX_ADDR_3\
        );

    \I__4566\ : Odrv12
    port map (
            O => \N__20189\,
            I => \RX_ADDR_3\
        );

    \I__4565\ : InMux
    port map (
            O => \N__20182\,
            I => \N__20179\
        );

    \I__4564\ : LocalMux
    port map (
            O => \N__20179\,
            I => \N__20167\
        );

    \I__4563\ : ClkMux
    port map (
            O => \N__20178\,
            I => \N__20029\
        );

    \I__4562\ : ClkMux
    port map (
            O => \N__20177\,
            I => \N__20029\
        );

    \I__4561\ : ClkMux
    port map (
            O => \N__20176\,
            I => \N__20029\
        );

    \I__4560\ : ClkMux
    port map (
            O => \N__20175\,
            I => \N__20029\
        );

    \I__4559\ : ClkMux
    port map (
            O => \N__20174\,
            I => \N__20029\
        );

    \I__4558\ : ClkMux
    port map (
            O => \N__20173\,
            I => \N__20029\
        );

    \I__4557\ : ClkMux
    port map (
            O => \N__20172\,
            I => \N__20029\
        );

    \I__4556\ : ClkMux
    port map (
            O => \N__20171\,
            I => \N__20029\
        );

    \I__4555\ : ClkMux
    port map (
            O => \N__20170\,
            I => \N__20029\
        );

    \I__4554\ : Glb2LocalMux
    port map (
            O => \N__20167\,
            I => \N__20029\
        );

    \I__4553\ : ClkMux
    port map (
            O => \N__20166\,
            I => \N__20029\
        );

    \I__4552\ : ClkMux
    port map (
            O => \N__20165\,
            I => \N__20029\
        );

    \I__4551\ : ClkMux
    port map (
            O => \N__20164\,
            I => \N__20029\
        );

    \I__4550\ : ClkMux
    port map (
            O => \N__20163\,
            I => \N__20029\
        );

    \I__4549\ : ClkMux
    port map (
            O => \N__20162\,
            I => \N__20029\
        );

    \I__4548\ : ClkMux
    port map (
            O => \N__20161\,
            I => \N__20029\
        );

    \I__4547\ : ClkMux
    port map (
            O => \N__20160\,
            I => \N__20029\
        );

    \I__4546\ : ClkMux
    port map (
            O => \N__20159\,
            I => \N__20029\
        );

    \I__4545\ : ClkMux
    port map (
            O => \N__20158\,
            I => \N__20029\
        );

    \I__4544\ : ClkMux
    port map (
            O => \N__20157\,
            I => \N__20029\
        );

    \I__4543\ : ClkMux
    port map (
            O => \N__20156\,
            I => \N__20029\
        );

    \I__4542\ : ClkMux
    port map (
            O => \N__20155\,
            I => \N__20029\
        );

    \I__4541\ : ClkMux
    port map (
            O => \N__20154\,
            I => \N__20029\
        );

    \I__4540\ : ClkMux
    port map (
            O => \N__20153\,
            I => \N__20029\
        );

    \I__4539\ : ClkMux
    port map (
            O => \N__20152\,
            I => \N__20029\
        );

    \I__4538\ : ClkMux
    port map (
            O => \N__20151\,
            I => \N__20029\
        );

    \I__4537\ : ClkMux
    port map (
            O => \N__20150\,
            I => \N__20029\
        );

    \I__4536\ : ClkMux
    port map (
            O => \N__20149\,
            I => \N__20029\
        );

    \I__4535\ : ClkMux
    port map (
            O => \N__20148\,
            I => \N__20029\
        );

    \I__4534\ : ClkMux
    port map (
            O => \N__20147\,
            I => \N__20029\
        );

    \I__4533\ : ClkMux
    port map (
            O => \N__20146\,
            I => \N__20029\
        );

    \I__4532\ : ClkMux
    port map (
            O => \N__20145\,
            I => \N__20029\
        );

    \I__4531\ : ClkMux
    port map (
            O => \N__20144\,
            I => \N__20029\
        );

    \I__4530\ : ClkMux
    port map (
            O => \N__20143\,
            I => \N__20029\
        );

    \I__4529\ : ClkMux
    port map (
            O => \N__20142\,
            I => \N__20029\
        );

    \I__4528\ : ClkMux
    port map (
            O => \N__20141\,
            I => \N__20029\
        );

    \I__4527\ : ClkMux
    port map (
            O => \N__20140\,
            I => \N__20029\
        );

    \I__4526\ : ClkMux
    port map (
            O => \N__20139\,
            I => \N__20029\
        );

    \I__4525\ : ClkMux
    port map (
            O => \N__20138\,
            I => \N__20029\
        );

    \I__4524\ : ClkMux
    port map (
            O => \N__20137\,
            I => \N__20029\
        );

    \I__4523\ : ClkMux
    port map (
            O => \N__20136\,
            I => \N__20029\
        );

    \I__4522\ : ClkMux
    port map (
            O => \N__20135\,
            I => \N__20029\
        );

    \I__4521\ : ClkMux
    port map (
            O => \N__20134\,
            I => \N__20029\
        );

    \I__4520\ : ClkMux
    port map (
            O => \N__20133\,
            I => \N__20029\
        );

    \I__4519\ : ClkMux
    port map (
            O => \N__20132\,
            I => \N__20029\
        );

    \I__4518\ : ClkMux
    port map (
            O => \N__20131\,
            I => \N__20029\
        );

    \I__4517\ : ClkMux
    port map (
            O => \N__20130\,
            I => \N__20029\
        );

    \I__4516\ : ClkMux
    port map (
            O => \N__20129\,
            I => \N__20029\
        );

    \I__4515\ : ClkMux
    port map (
            O => \N__20128\,
            I => \N__20029\
        );

    \I__4514\ : GlobalMux
    port map (
            O => \N__20029\,
            I => \N__20026\
        );

    \I__4513\ : gio2CtrlBuf
    port map (
            O => \N__20026\,
            I => \TVP_CLK_c\
        );

    \I__4512\ : InMux
    port map (
            O => \N__20023\,
            I => \N__20020\
        );

    \I__4511\ : LocalMux
    port map (
            O => \N__20020\,
            I => \transmit_module.Y_DELTA_PATTERN_32\
        );

    \I__4510\ : InMux
    port map (
            O => \N__20017\,
            I => \N__20014\
        );

    \I__4509\ : LocalMux
    port map (
            O => \N__20014\,
            I => \transmit_module.Y_DELTA_PATTERN_31\
        );

    \I__4508\ : InMux
    port map (
            O => \N__20011\,
            I => \N__20008\
        );

    \I__4507\ : LocalMux
    port map (
            O => \N__20008\,
            I => \transmit_module.Y_DELTA_PATTERN_22\
        );

    \I__4506\ : InMux
    port map (
            O => \N__20005\,
            I => \N__20002\
        );

    \I__4505\ : LocalMux
    port map (
            O => \N__20002\,
            I => \transmit_module.Y_DELTA_PATTERN_24\
        );

    \I__4504\ : InMux
    port map (
            O => \N__19999\,
            I => \N__19996\
        );

    \I__4503\ : LocalMux
    port map (
            O => \N__19996\,
            I => \transmit_module.Y_DELTA_PATTERN_23\
        );

    \I__4502\ : InMux
    port map (
            O => \N__19993\,
            I => \N__19990\
        );

    \I__4501\ : LocalMux
    port map (
            O => \N__19990\,
            I => \transmit_module.Y_DELTA_PATTERN_16\
        );

    \I__4500\ : InMux
    port map (
            O => \N__19987\,
            I => \N__19984\
        );

    \I__4499\ : LocalMux
    port map (
            O => \N__19984\,
            I => \transmit_module.Y_DELTA_PATTERN_17\
        );

    \I__4498\ : InMux
    port map (
            O => \N__19981\,
            I => \N__19978\
        );

    \I__4497\ : LocalMux
    port map (
            O => \N__19978\,
            I => \transmit_module.Y_DELTA_PATTERN_19\
        );

    \I__4496\ : InMux
    port map (
            O => \N__19975\,
            I => \N__19972\
        );

    \I__4495\ : LocalMux
    port map (
            O => \N__19972\,
            I => \transmit_module.Y_DELTA_PATTERN_18\
        );

    \I__4494\ : InMux
    port map (
            O => \N__19969\,
            I => \N__19966\
        );

    \I__4493\ : LocalMux
    port map (
            O => \N__19966\,
            I => \N__19963\
        );

    \I__4492\ : Odrv12
    port map (
            O => \N__19963\,
            I => \line_buffer.n3737\
        );

    \I__4491\ : InMux
    port map (
            O => \N__19960\,
            I => \N__19957\
        );

    \I__4490\ : LocalMux
    port map (
            O => \N__19957\,
            I => \N__19954\
        );

    \I__4489\ : Span4Mux_h
    port map (
            O => \N__19954\,
            I => \N__19951\
        );

    \I__4488\ : Span4Mux_h
    port map (
            O => \N__19951\,
            I => \N__19948\
        );

    \I__4487\ : Odrv4
    port map (
            O => \N__19948\,
            I => \line_buffer.n447\
        );

    \I__4486\ : CascadeMux
    port map (
            O => \N__19945\,
            I => \N__19942\
        );

    \I__4485\ : InMux
    port map (
            O => \N__19942\,
            I => \N__19939\
        );

    \I__4484\ : LocalMux
    port map (
            O => \N__19939\,
            I => \N__19936\
        );

    \I__4483\ : Span4Mux_v
    port map (
            O => \N__19936\,
            I => \N__19933\
        );

    \I__4482\ : Sp12to4
    port map (
            O => \N__19933\,
            I => \N__19930\
        );

    \I__4481\ : Span12Mux_h
    port map (
            O => \N__19930\,
            I => \N__19927\
        );

    \I__4480\ : Odrv12
    port map (
            O => \N__19927\,
            I => \line_buffer.n439\
        );

    \I__4479\ : InMux
    port map (
            O => \N__19924\,
            I => \N__19921\
        );

    \I__4478\ : LocalMux
    port map (
            O => \N__19921\,
            I => \line_buffer.n3701\
        );

    \I__4477\ : InMux
    port map (
            O => \N__19918\,
            I => \N__19915\
        );

    \I__4476\ : LocalMux
    port map (
            O => \N__19915\,
            I => \N__19912\
        );

    \I__4475\ : Odrv12
    port map (
            O => \N__19912\,
            I => \TX_DATA_5\
        );

    \I__4474\ : IoInMux
    port map (
            O => \N__19909\,
            I => \N__19906\
        );

    \I__4473\ : LocalMux
    port map (
            O => \N__19906\,
            I => \N__19902\
        );

    \I__4472\ : IoInMux
    port map (
            O => \N__19905\,
            I => \N__19899\
        );

    \I__4471\ : IoSpan4Mux
    port map (
            O => \N__19902\,
            I => \N__19895\
        );

    \I__4470\ : LocalMux
    port map (
            O => \N__19899\,
            I => \N__19892\
        );

    \I__4469\ : IoInMux
    port map (
            O => \N__19898\,
            I => \N__19889\
        );

    \I__4468\ : Span4Mux_s3_v
    port map (
            O => \N__19895\,
            I => \N__19886\
        );

    \I__4467\ : Span4Mux_s3_v
    port map (
            O => \N__19892\,
            I => \N__19883\
        );

    \I__4466\ : LocalMux
    port map (
            O => \N__19889\,
            I => \N__19880\
        );

    \I__4465\ : Span4Mux_h
    port map (
            O => \N__19886\,
            I => \N__19877\
        );

    \I__4464\ : Span4Mux_h
    port map (
            O => \N__19883\,
            I => \N__19874\
        );

    \I__4463\ : Span12Mux_s4_h
    port map (
            O => \N__19880\,
            I => \N__19871\
        );

    \I__4462\ : Span4Mux_h
    port map (
            O => \N__19877\,
            I => \N__19866\
        );

    \I__4461\ : Span4Mux_h
    port map (
            O => \N__19874\,
            I => \N__19866\
        );

    \I__4460\ : Span12Mux_h
    port map (
            O => \N__19871\,
            I => \N__19863\
        );

    \I__4459\ : Span4Mux_v
    port map (
            O => \N__19866\,
            I => \N__19860\
        );

    \I__4458\ : Odrv12
    port map (
            O => \N__19863\,
            I => n1793
        );

    \I__4457\ : Odrv4
    port map (
            O => \N__19860\,
            I => n1793
        );

    \I__4456\ : SRMux
    port map (
            O => \N__19855\,
            I => \N__19852\
        );

    \I__4455\ : LocalMux
    port map (
            O => \N__19852\,
            I => \N__19847\
        );

    \I__4454\ : SRMux
    port map (
            O => \N__19851\,
            I => \N__19844\
        );

    \I__4453\ : SRMux
    port map (
            O => \N__19850\,
            I => \N__19840\
        );

    \I__4452\ : Span4Mux_v
    port map (
            O => \N__19847\,
            I => \N__19833\
        );

    \I__4451\ : LocalMux
    port map (
            O => \N__19844\,
            I => \N__19833\
        );

    \I__4450\ : SRMux
    port map (
            O => \N__19843\,
            I => \N__19830\
        );

    \I__4449\ : LocalMux
    port map (
            O => \N__19840\,
            I => \N__19826\
        );

    \I__4448\ : SRMux
    port map (
            O => \N__19839\,
            I => \N__19823\
        );

    \I__4447\ : SRMux
    port map (
            O => \N__19838\,
            I => \N__19820\
        );

    \I__4446\ : Span4Mux_h
    port map (
            O => \N__19833\,
            I => \N__19813\
        );

    \I__4445\ : LocalMux
    port map (
            O => \N__19830\,
            I => \N__19813\
        );

    \I__4444\ : SRMux
    port map (
            O => \N__19829\,
            I => \N__19810\
        );

    \I__4443\ : Span4Mux_s0_v
    port map (
            O => \N__19826\,
            I => \N__19802\
        );

    \I__4442\ : LocalMux
    port map (
            O => \N__19823\,
            I => \N__19802\
        );

    \I__4441\ : LocalMux
    port map (
            O => \N__19820\,
            I => \N__19799\
        );

    \I__4440\ : SRMux
    port map (
            O => \N__19819\,
            I => \N__19796\
        );

    \I__4439\ : SRMux
    port map (
            O => \N__19818\,
            I => \N__19793\
        );

    \I__4438\ : Span4Mux_v
    port map (
            O => \N__19813\,
            I => \N__19786\
        );

    \I__4437\ : LocalMux
    port map (
            O => \N__19810\,
            I => \N__19786\
        );

    \I__4436\ : SRMux
    port map (
            O => \N__19809\,
            I => \N__19783\
        );

    \I__4435\ : SRMux
    port map (
            O => \N__19808\,
            I => \N__19780\
        );

    \I__4434\ : SRMux
    port map (
            O => \N__19807\,
            I => \N__19777\
        );

    \I__4433\ : Span4Mux_v
    port map (
            O => \N__19802\,
            I => \N__19769\
        );

    \I__4432\ : Span4Mux_h
    port map (
            O => \N__19799\,
            I => \N__19769\
        );

    \I__4431\ : LocalMux
    port map (
            O => \N__19796\,
            I => \N__19769\
        );

    \I__4430\ : LocalMux
    port map (
            O => \N__19793\,
            I => \N__19766\
        );

    \I__4429\ : SRMux
    port map (
            O => \N__19792\,
            I => \N__19763\
        );

    \I__4428\ : SRMux
    port map (
            O => \N__19791\,
            I => \N__19760\
        );

    \I__4427\ : Span4Mux_h
    port map (
            O => \N__19786\,
            I => \N__19752\
        );

    \I__4426\ : LocalMux
    port map (
            O => \N__19783\,
            I => \N__19752\
        );

    \I__4425\ : LocalMux
    port map (
            O => \N__19780\,
            I => \N__19747\
        );

    \I__4424\ : LocalMux
    port map (
            O => \N__19777\,
            I => \N__19747\
        );

    \I__4423\ : SRMux
    port map (
            O => \N__19776\,
            I => \N__19744\
        );

    \I__4422\ : Span4Mux_v
    port map (
            O => \N__19769\,
            I => \N__19739\
        );

    \I__4421\ : Span4Mux_h
    port map (
            O => \N__19766\,
            I => \N__19734\
        );

    \I__4420\ : LocalMux
    port map (
            O => \N__19763\,
            I => \N__19734\
        );

    \I__4419\ : LocalMux
    port map (
            O => \N__19760\,
            I => \N__19731\
        );

    \I__4418\ : SRMux
    port map (
            O => \N__19759\,
            I => \N__19728\
        );

    \I__4417\ : SRMux
    port map (
            O => \N__19758\,
            I => \N__19725\
        );

    \I__4416\ : SRMux
    port map (
            O => \N__19757\,
            I => \N__19720\
        );

    \I__4415\ : Span4Mux_v
    port map (
            O => \N__19752\,
            I => \N__19715\
        );

    \I__4414\ : Span4Mux_v
    port map (
            O => \N__19747\,
            I => \N__19712\
        );

    \I__4413\ : LocalMux
    port map (
            O => \N__19744\,
            I => \N__19709\
        );

    \I__4412\ : SRMux
    port map (
            O => \N__19743\,
            I => \N__19706\
        );

    \I__4411\ : SRMux
    port map (
            O => \N__19742\,
            I => \N__19701\
        );

    \I__4410\ : Span4Mux_v
    port map (
            O => \N__19739\,
            I => \N__19690\
        );

    \I__4409\ : Span4Mux_v
    port map (
            O => \N__19734\,
            I => \N__19690\
        );

    \I__4408\ : Span4Mux_h
    port map (
            O => \N__19731\,
            I => \N__19690\
        );

    \I__4407\ : LocalMux
    port map (
            O => \N__19728\,
            I => \N__19690\
        );

    \I__4406\ : LocalMux
    port map (
            O => \N__19725\,
            I => \N__19687\
        );

    \I__4405\ : SRMux
    port map (
            O => \N__19724\,
            I => \N__19684\
        );

    \I__4404\ : SRMux
    port map (
            O => \N__19723\,
            I => \N__19681\
        );

    \I__4403\ : LocalMux
    port map (
            O => \N__19720\,
            I => \N__19677\
        );

    \I__4402\ : SRMux
    port map (
            O => \N__19719\,
            I => \N__19674\
        );

    \I__4401\ : SRMux
    port map (
            O => \N__19718\,
            I => \N__19671\
        );

    \I__4400\ : Span4Mux_v
    port map (
            O => \N__19715\,
            I => \N__19668\
        );

    \I__4399\ : Span4Mux_v
    port map (
            O => \N__19712\,
            I => \N__19661\
        );

    \I__4398\ : Span4Mux_v
    port map (
            O => \N__19709\,
            I => \N__19661\
        );

    \I__4397\ : LocalMux
    port map (
            O => \N__19706\,
            I => \N__19661\
        );

    \I__4396\ : SRMux
    port map (
            O => \N__19705\,
            I => \N__19658\
        );

    \I__4395\ : SRMux
    port map (
            O => \N__19704\,
            I => \N__19653\
        );

    \I__4394\ : LocalMux
    port map (
            O => \N__19701\,
            I => \N__19649\
        );

    \I__4393\ : SRMux
    port map (
            O => \N__19700\,
            I => \N__19646\
        );

    \I__4392\ : SRMux
    port map (
            O => \N__19699\,
            I => \N__19643\
        );

    \I__4391\ : Span4Mux_v
    port map (
            O => \N__19690\,
            I => \N__19636\
        );

    \I__4390\ : Span4Mux_h
    port map (
            O => \N__19687\,
            I => \N__19636\
        );

    \I__4389\ : LocalMux
    port map (
            O => \N__19684\,
            I => \N__19636\
        );

    \I__4388\ : LocalMux
    port map (
            O => \N__19681\,
            I => \N__19633\
        );

    \I__4387\ : SRMux
    port map (
            O => \N__19680\,
            I => \N__19630\
        );

    \I__4386\ : Span4Mux_s3_v
    port map (
            O => \N__19677\,
            I => \N__19622\
        );

    \I__4385\ : LocalMux
    port map (
            O => \N__19674\,
            I => \N__19622\
        );

    \I__4384\ : LocalMux
    port map (
            O => \N__19671\,
            I => \N__19622\
        );

    \I__4383\ : Span4Mux_v
    port map (
            O => \N__19668\,
            I => \N__19615\
        );

    \I__4382\ : Span4Mux_h
    port map (
            O => \N__19661\,
            I => \N__19615\
        );

    \I__4381\ : LocalMux
    port map (
            O => \N__19658\,
            I => \N__19615\
        );

    \I__4380\ : IoInMux
    port map (
            O => \N__19657\,
            I => \N__19612\
        );

    \I__4379\ : IoInMux
    port map (
            O => \N__19656\,
            I => \N__19609\
        );

    \I__4378\ : LocalMux
    port map (
            O => \N__19653\,
            I => \N__19606\
        );

    \I__4377\ : SRMux
    port map (
            O => \N__19652\,
            I => \N__19603\
        );

    \I__4376\ : Span4Mux_s3_v
    port map (
            O => \N__19649\,
            I => \N__19595\
        );

    \I__4375\ : LocalMux
    port map (
            O => \N__19646\,
            I => \N__19595\
        );

    \I__4374\ : LocalMux
    port map (
            O => \N__19643\,
            I => \N__19595\
        );

    \I__4373\ : Span4Mux_v
    port map (
            O => \N__19636\,
            I => \N__19588\
        );

    \I__4372\ : Span4Mux_h
    port map (
            O => \N__19633\,
            I => \N__19588\
        );

    \I__4371\ : LocalMux
    port map (
            O => \N__19630\,
            I => \N__19588\
        );

    \I__4370\ : SRMux
    port map (
            O => \N__19629\,
            I => \N__19585\
        );

    \I__4369\ : Span4Mux_v
    port map (
            O => \N__19622\,
            I => \N__19580\
        );

    \I__4368\ : Span4Mux_v
    port map (
            O => \N__19615\,
            I => \N__19580\
        );

    \I__4367\ : LocalMux
    port map (
            O => \N__19612\,
            I => \N__19575\
        );

    \I__4366\ : LocalMux
    port map (
            O => \N__19609\,
            I => \N__19575\
        );

    \I__4365\ : Span12Mux_s9_h
    port map (
            O => \N__19606\,
            I => \N__19572\
        );

    \I__4364\ : LocalMux
    port map (
            O => \N__19603\,
            I => \N__19569\
        );

    \I__4363\ : SRMux
    port map (
            O => \N__19602\,
            I => \N__19566\
        );

    \I__4362\ : Span4Mux_v
    port map (
            O => \N__19595\,
            I => \N__19563\
        );

    \I__4361\ : Span4Mux_v
    port map (
            O => \N__19588\,
            I => \N__19558\
        );

    \I__4360\ : LocalMux
    port map (
            O => \N__19585\,
            I => \N__19558\
        );

    \I__4359\ : Span4Mux_h
    port map (
            O => \N__19580\,
            I => \N__19555\
        );

    \I__4358\ : Span4Mux_s3_v
    port map (
            O => \N__19575\,
            I => \N__19552\
        );

    \I__4357\ : Span12Mux_v
    port map (
            O => \N__19572\,
            I => \N__19547\
        );

    \I__4356\ : Span12Mux_s9_h
    port map (
            O => \N__19569\,
            I => \N__19547\
        );

    \I__4355\ : LocalMux
    port map (
            O => \N__19566\,
            I => \N__19544\
        );

    \I__4354\ : Span4Mux_h
    port map (
            O => \N__19563\,
            I => \N__19539\
        );

    \I__4353\ : Span4Mux_h
    port map (
            O => \N__19558\,
            I => \N__19539\
        );

    \I__4352\ : Span4Mux_h
    port map (
            O => \N__19555\,
            I => \N__19534\
        );

    \I__4351\ : Span4Mux_v
    port map (
            O => \N__19552\,
            I => \N__19534\
        );

    \I__4350\ : Span12Mux_v
    port map (
            O => \N__19547\,
            I => \N__19529\
        );

    \I__4349\ : Span12Mux_s9_h
    port map (
            O => \N__19544\,
            I => \N__19529\
        );

    \I__4348\ : Span4Mux_h
    port map (
            O => \N__19539\,
            I => \N__19526\
        );

    \I__4347\ : Odrv4
    port map (
            O => \N__19534\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4346\ : Odrv12
    port map (
            O => \N__19529\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4345\ : Odrv4
    port map (
            O => \N__19526\,
            I => \CONSTANT_ONE_NET\
        );

    \I__4344\ : InMux
    port map (
            O => \N__19519\,
            I => \N__19516\
        );

    \I__4343\ : LocalMux
    port map (
            O => \N__19516\,
            I => \N__19513\
        );

    \I__4342\ : Span4Mux_h
    port map (
            O => \N__19513\,
            I => \N__19510\
        );

    \I__4341\ : Span4Mux_h
    port map (
            O => \N__19510\,
            I => \N__19507\
        );

    \I__4340\ : Odrv4
    port map (
            O => \N__19507\,
            I => \transmit_module.Y_DELTA_PATTERN_33\
        );

    \I__4339\ : InMux
    port map (
            O => \N__19504\,
            I => \N__19501\
        );

    \I__4338\ : LocalMux
    port map (
            O => \N__19501\,
            I => \N__19498\
        );

    \I__4337\ : Odrv4
    port map (
            O => \N__19498\,
            I => \transmit_module.Y_DELTA_PATTERN_27\
        );

    \I__4336\ : InMux
    port map (
            O => \N__19495\,
            I => \N__19492\
        );

    \I__4335\ : LocalMux
    port map (
            O => \N__19492\,
            I => \transmit_module.Y_DELTA_PATTERN_28\
        );

    \I__4334\ : InMux
    port map (
            O => \N__19489\,
            I => \N__19486\
        );

    \I__4333\ : LocalMux
    port map (
            O => \N__19486\,
            I => \transmit_module.Y_DELTA_PATTERN_29\
        );

    \I__4332\ : InMux
    port map (
            O => \N__19483\,
            I => \N__19480\
        );

    \I__4331\ : LocalMux
    port map (
            O => \N__19480\,
            I => \transmit_module.Y_DELTA_PATTERN_30\
        );

    \I__4330\ : InMux
    port map (
            O => \N__19477\,
            I => \N__19474\
        );

    \I__4329\ : LocalMux
    port map (
            O => \N__19474\,
            I => \transmit_module.Y_DELTA_PATTERN_12\
        );

    \I__4328\ : InMux
    port map (
            O => \N__19471\,
            I => \N__19468\
        );

    \I__4327\ : LocalMux
    port map (
            O => \N__19468\,
            I => \N__19465\
        );

    \I__4326\ : Span4Mux_h
    port map (
            O => \N__19465\,
            I => \N__19462\
        );

    \I__4325\ : Odrv4
    port map (
            O => \N__19462\,
            I => \transmit_module.Y_DELTA_PATTERN_11\
        );

    \I__4324\ : InMux
    port map (
            O => \N__19459\,
            I => \N__19456\
        );

    \I__4323\ : LocalMux
    port map (
            O => \N__19456\,
            I => \transmit_module.Y_DELTA_PATTERN_25\
        );

    \I__4322\ : InMux
    port map (
            O => \N__19453\,
            I => \N__19450\
        );

    \I__4321\ : LocalMux
    port map (
            O => \N__19450\,
            I => \transmit_module.Y_DELTA_PATTERN_26\
        );

    \I__4320\ : InMux
    port map (
            O => \N__19447\,
            I => \N__19444\
        );

    \I__4319\ : LocalMux
    port map (
            O => \N__19444\,
            I => \transmit_module.Y_DELTA_PATTERN_13\
        );

    \I__4318\ : InMux
    port map (
            O => \N__19441\,
            I => \N__19438\
        );

    \I__4317\ : LocalMux
    port map (
            O => \N__19438\,
            I => \N__19435\
        );

    \I__4316\ : Span12Mux_h
    port map (
            O => \N__19435\,
            I => \N__19432\
        );

    \I__4315\ : Odrv12
    port map (
            O => \N__19432\,
            I => \line_buffer.n539\
        );

    \I__4314\ : InMux
    port map (
            O => \N__19429\,
            I => \N__19426\
        );

    \I__4313\ : LocalMux
    port map (
            O => \N__19426\,
            I => \N__19423\
        );

    \I__4312\ : Span4Mux_h
    port map (
            O => \N__19423\,
            I => \N__19420\
        );

    \I__4311\ : Span4Mux_h
    port map (
            O => \N__19420\,
            I => \N__19417\
        );

    \I__4310\ : Odrv4
    port map (
            O => \N__19417\,
            I => \line_buffer.n531\
        );

    \I__4309\ : InMux
    port map (
            O => \N__19414\,
            I => \N__19411\
        );

    \I__4308\ : LocalMux
    port map (
            O => \N__19411\,
            I => \line_buffer.n3746\
        );

    \I__4307\ : InMux
    port map (
            O => \N__19408\,
            I => \N__19405\
        );

    \I__4306\ : LocalMux
    port map (
            O => \N__19405\,
            I => \N__19402\
        );

    \I__4305\ : Span4Mux_v
    port map (
            O => \N__19402\,
            I => \N__19399\
        );

    \I__4304\ : Sp12to4
    port map (
            O => \N__19399\,
            I => \N__19396\
        );

    \I__4303\ : Odrv12
    port map (
            O => \N__19396\,
            I => \line_buffer.n573\
        );

    \I__4302\ : InMux
    port map (
            O => \N__19393\,
            I => \N__19390\
        );

    \I__4301\ : LocalMux
    port map (
            O => \N__19390\,
            I => \N__19387\
        );

    \I__4300\ : Sp12to4
    port map (
            O => \N__19387\,
            I => \N__19384\
        );

    \I__4299\ : Span12Mux_v
    port map (
            O => \N__19384\,
            I => \N__19381\
        );

    \I__4298\ : Odrv12
    port map (
            O => \N__19381\,
            I => \line_buffer.n565\
        );

    \I__4297\ : InMux
    port map (
            O => \N__19378\,
            I => \N__19375\
        );

    \I__4296\ : LocalMux
    port map (
            O => \N__19375\,
            I => \line_buffer.n3677\
        );

    \I__4295\ : InMux
    port map (
            O => \N__19372\,
            I => \N__19369\
        );

    \I__4294\ : LocalMux
    port map (
            O => \N__19369\,
            I => \N__19366\
        );

    \I__4293\ : Span12Mux_v
    port map (
            O => \N__19366\,
            I => \N__19363\
        );

    \I__4292\ : Odrv12
    port map (
            O => \N__19363\,
            I => \line_buffer.n567\
        );

    \I__4291\ : InMux
    port map (
            O => \N__19360\,
            I => \N__19357\
        );

    \I__4290\ : LocalMux
    port map (
            O => \N__19357\,
            I => \N__19354\
        );

    \I__4289\ : Span4Mux_v
    port map (
            O => \N__19354\,
            I => \N__19351\
        );

    \I__4288\ : Sp12to4
    port map (
            O => \N__19351\,
            I => \N__19348\
        );

    \I__4287\ : Odrv12
    port map (
            O => \N__19348\,
            I => \line_buffer.n575\
        );

    \I__4286\ : InMux
    port map (
            O => \N__19345\,
            I => \N__19342\
        );

    \I__4285\ : LocalMux
    port map (
            O => \N__19342\,
            I => \line_buffer.n3635\
        );

    \I__4284\ : InMux
    port map (
            O => \N__19339\,
            I => \N__19334\
        );

    \I__4283\ : InMux
    port map (
            O => \N__19338\,
            I => \N__19329\
        );

    \I__4282\ : InMux
    port map (
            O => \N__19337\,
            I => \N__19329\
        );

    \I__4281\ : LocalMux
    port map (
            O => \N__19334\,
            I => \receive_module.rx_counter.X_4\
        );

    \I__4280\ : LocalMux
    port map (
            O => \N__19329\,
            I => \receive_module.rx_counter.X_4\
        );

    \I__4279\ : InMux
    port map (
            O => \N__19324\,
            I => \receive_module.rx_counter.n3304\
        );

    \I__4278\ : InMux
    port map (
            O => \N__19321\,
            I => \N__19316\
        );

    \I__4277\ : InMux
    port map (
            O => \N__19320\,
            I => \N__19311\
        );

    \I__4276\ : InMux
    port map (
            O => \N__19319\,
            I => \N__19311\
        );

    \I__4275\ : LocalMux
    port map (
            O => \N__19316\,
            I => \receive_module.rx_counter.X_5\
        );

    \I__4274\ : LocalMux
    port map (
            O => \N__19311\,
            I => \receive_module.rx_counter.X_5\
        );

    \I__4273\ : InMux
    port map (
            O => \N__19306\,
            I => \receive_module.rx_counter.n3305\
        );

    \I__4272\ : InMux
    port map (
            O => \N__19303\,
            I => \N__19298\
        );

    \I__4271\ : InMux
    port map (
            O => \N__19302\,
            I => \N__19293\
        );

    \I__4270\ : InMux
    port map (
            O => \N__19301\,
            I => \N__19293\
        );

    \I__4269\ : LocalMux
    port map (
            O => \N__19298\,
            I => \receive_module.rx_counter.X_6\
        );

    \I__4268\ : LocalMux
    port map (
            O => \N__19293\,
            I => \receive_module.rx_counter.X_6\
        );

    \I__4267\ : InMux
    port map (
            O => \N__19288\,
            I => \receive_module.rx_counter.n3306\
        );

    \I__4266\ : InMux
    port map (
            O => \N__19285\,
            I => \N__19280\
        );

    \I__4265\ : InMux
    port map (
            O => \N__19284\,
            I => \N__19275\
        );

    \I__4264\ : InMux
    port map (
            O => \N__19283\,
            I => \N__19275\
        );

    \I__4263\ : LocalMux
    port map (
            O => \N__19280\,
            I => \receive_module.rx_counter.X_7\
        );

    \I__4262\ : LocalMux
    port map (
            O => \N__19275\,
            I => \receive_module.rx_counter.X_7\
        );

    \I__4261\ : InMux
    port map (
            O => \N__19270\,
            I => \receive_module.rx_counter.n3307\
        );

    \I__4260\ : InMux
    port map (
            O => \N__19267\,
            I => \N__19263\
        );

    \I__4259\ : InMux
    port map (
            O => \N__19266\,
            I => \N__19260\
        );

    \I__4258\ : LocalMux
    port map (
            O => \N__19263\,
            I => \receive_module.rx_counter.X_8\
        );

    \I__4257\ : LocalMux
    port map (
            O => \N__19260\,
            I => \receive_module.rx_counter.X_8\
        );

    \I__4256\ : InMux
    port map (
            O => \N__19255\,
            I => \bfn_17_11_0_\
        );

    \I__4255\ : InMux
    port map (
            O => \N__19252\,
            I => \receive_module.rx_counter.n3309\
        );

    \I__4254\ : CascadeMux
    port map (
            O => \N__19249\,
            I => \N__19245\
        );

    \I__4253\ : InMux
    port map (
            O => \N__19248\,
            I => \N__19242\
        );

    \I__4252\ : InMux
    port map (
            O => \N__19245\,
            I => \N__19239\
        );

    \I__4251\ : LocalMux
    port map (
            O => \N__19242\,
            I => \receive_module.rx_counter.X_9\
        );

    \I__4250\ : LocalMux
    port map (
            O => \N__19239\,
            I => \receive_module.rx_counter.X_9\
        );

    \I__4249\ : SRMux
    port map (
            O => \N__19234\,
            I => \N__19230\
        );

    \I__4248\ : SRMux
    port map (
            O => \N__19233\,
            I => \N__19227\
        );

    \I__4247\ : LocalMux
    port map (
            O => \N__19230\,
            I => \N__19224\
        );

    \I__4246\ : LocalMux
    port map (
            O => \N__19227\,
            I => \N__19221\
        );

    \I__4245\ : Span4Mux_h
    port map (
            O => \N__19224\,
            I => \N__19218\
        );

    \I__4244\ : Odrv4
    port map (
            O => \N__19221\,
            I => \receive_module.rx_counter.n3790\
        );

    \I__4243\ : Odrv4
    port map (
            O => \N__19218\,
            I => \receive_module.rx_counter.n3790\
        );

    \I__4242\ : InMux
    port map (
            O => \N__19213\,
            I => \N__19210\
        );

    \I__4241\ : LocalMux
    port map (
            O => \N__19210\,
            I => \N__19207\
        );

    \I__4240\ : Odrv12
    port map (
            O => \N__19207\,
            I => \line_buffer.n576\
        );

    \I__4239\ : InMux
    port map (
            O => \N__19204\,
            I => \N__19201\
        );

    \I__4238\ : LocalMux
    port map (
            O => \N__19201\,
            I => \N__19198\
        );

    \I__4237\ : Span12Mux_v
    port map (
            O => \N__19198\,
            I => \N__19195\
        );

    \I__4236\ : Span12Mux_v
    port map (
            O => \N__19195\,
            I => \N__19192\
        );

    \I__4235\ : Odrv12
    port map (
            O => \N__19192\,
            I => \line_buffer.n568\
        );

    \I__4234\ : InMux
    port map (
            O => \N__19189\,
            I => \N__19186\
        );

    \I__4233\ : LocalMux
    port map (
            O => \N__19186\,
            I => \N__19183\
        );

    \I__4232\ : Sp12to4
    port map (
            O => \N__19183\,
            I => \N__19180\
        );

    \I__4231\ : Span12Mux_v
    port map (
            O => \N__19180\,
            I => \N__19177\
        );

    \I__4230\ : Odrv12
    port map (
            O => \N__19177\,
            I => \line_buffer.n504\
        );

    \I__4229\ : InMux
    port map (
            O => \N__19174\,
            I => \N__19171\
        );

    \I__4228\ : LocalMux
    port map (
            O => \N__19171\,
            I => \N__19168\
        );

    \I__4227\ : Span12Mux_h
    port map (
            O => \N__19168\,
            I => \N__19165\
        );

    \I__4226\ : Span12Mux_v
    port map (
            O => \N__19165\,
            I => \N__19162\
        );

    \I__4225\ : Odrv12
    port map (
            O => \N__19162\,
            I => \line_buffer.n512\
        );

    \I__4224\ : CascadeMux
    port map (
            O => \N__19159\,
            I => \line_buffer.n3734_cascade_\
        );

    \I__4223\ : InMux
    port map (
            O => \N__19156\,
            I => \N__19153\
        );

    \I__4222\ : LocalMux
    port map (
            O => \N__19153\,
            I => \N__19150\
        );

    \I__4221\ : Span4Mux_v
    port map (
            O => \N__19150\,
            I => \N__19147\
        );

    \I__4220\ : Sp12to4
    port map (
            O => \N__19147\,
            I => \N__19144\
        );

    \I__4219\ : Odrv12
    port map (
            O => \N__19144\,
            I => \line_buffer.n444\
        );

    \I__4218\ : InMux
    port map (
            O => \N__19141\,
            I => \N__19138\
        );

    \I__4217\ : LocalMux
    port map (
            O => \N__19138\,
            I => \N__19135\
        );

    \I__4216\ : Span4Mux_v
    port map (
            O => \N__19135\,
            I => \N__19132\
        );

    \I__4215\ : Sp12to4
    port map (
            O => \N__19132\,
            I => \N__19129\
        );

    \I__4214\ : Span12Mux_h
    port map (
            O => \N__19129\,
            I => \N__19126\
        );

    \I__4213\ : Odrv12
    port map (
            O => \N__19126\,
            I => \line_buffer.n436\
        );

    \I__4212\ : InMux
    port map (
            O => \N__19123\,
            I => \N__19120\
        );

    \I__4211\ : LocalMux
    port map (
            O => \N__19120\,
            I => \N__19117\
        );

    \I__4210\ : Odrv12
    port map (
            O => \N__19117\,
            I => \line_buffer.n3673\
        );

    \I__4209\ : InMux
    port map (
            O => \N__19114\,
            I => \N__19110\
        );

    \I__4208\ : InMux
    port map (
            O => \N__19113\,
            I => \N__19106\
        );

    \I__4207\ : LocalMux
    port map (
            O => \N__19110\,
            I => \N__19103\
        );

    \I__4206\ : InMux
    port map (
            O => \N__19109\,
            I => \N__19100\
        );

    \I__4205\ : LocalMux
    port map (
            O => \N__19106\,
            I => \N__19094\
        );

    \I__4204\ : Span4Mux_h
    port map (
            O => \N__19103\,
            I => \N__19090\
        );

    \I__4203\ : LocalMux
    port map (
            O => \N__19100\,
            I => \N__19087\
        );

    \I__4202\ : CascadeMux
    port map (
            O => \N__19099\,
            I => \N__19083\
        );

    \I__4201\ : InMux
    port map (
            O => \N__19098\,
            I => \N__19072\
        );

    \I__4200\ : InMux
    port map (
            O => \N__19097\,
            I => \N__19072\
        );

    \I__4199\ : Span4Mux_h
    port map (
            O => \N__19094\,
            I => \N__19069\
        );

    \I__4198\ : InMux
    port map (
            O => \N__19093\,
            I => \N__19061\
        );

    \I__4197\ : Span4Mux_v
    port map (
            O => \N__19090\,
            I => \N__19054\
        );

    \I__4196\ : Span4Mux_h
    port map (
            O => \N__19087\,
            I => \N__19054\
        );

    \I__4195\ : InMux
    port map (
            O => \N__19086\,
            I => \N__19051\
        );

    \I__4194\ : InMux
    port map (
            O => \N__19083\,
            I => \N__19048\
        );

    \I__4193\ : InMux
    port map (
            O => \N__19082\,
            I => \N__19043\
        );

    \I__4192\ : InMux
    port map (
            O => \N__19081\,
            I => \N__19043\
        );

    \I__4191\ : InMux
    port map (
            O => \N__19080\,
            I => \N__19034\
        );

    \I__4190\ : InMux
    port map (
            O => \N__19079\,
            I => \N__19034\
        );

    \I__4189\ : InMux
    port map (
            O => \N__19078\,
            I => \N__19034\
        );

    \I__4188\ : InMux
    port map (
            O => \N__19077\,
            I => \N__19034\
        );

    \I__4187\ : LocalMux
    port map (
            O => \N__19072\,
            I => \N__19031\
        );

    \I__4186\ : Span4Mux_v
    port map (
            O => \N__19069\,
            I => \N__19028\
        );

    \I__4185\ : InMux
    port map (
            O => \N__19068\,
            I => \N__19025\
        );

    \I__4184\ : InMux
    port map (
            O => \N__19067\,
            I => \N__19019\
        );

    \I__4183\ : InMux
    port map (
            O => \N__19066\,
            I => \N__19014\
        );

    \I__4182\ : InMux
    port map (
            O => \N__19065\,
            I => \N__19014\
        );

    \I__4181\ : InMux
    port map (
            O => \N__19064\,
            I => \N__19011\
        );

    \I__4180\ : LocalMux
    port map (
            O => \N__19061\,
            I => \N__19008\
        );

    \I__4179\ : InMux
    port map (
            O => \N__19060\,
            I => \N__19003\
        );

    \I__4178\ : InMux
    port map (
            O => \N__19059\,
            I => \N__19003\
        );

    \I__4177\ : Span4Mux_v
    port map (
            O => \N__19054\,
            I => \N__18998\
        );

    \I__4176\ : LocalMux
    port map (
            O => \N__19051\,
            I => \N__18998\
        );

    \I__4175\ : LocalMux
    port map (
            O => \N__19048\,
            I => \N__18993\
        );

    \I__4174\ : LocalMux
    port map (
            O => \N__19043\,
            I => \N__18993\
        );

    \I__4173\ : LocalMux
    port map (
            O => \N__19034\,
            I => \N__18990\
        );

    \I__4172\ : Span4Mux_h
    port map (
            O => \N__19031\,
            I => \N__18982\
        );

    \I__4171\ : Span4Mux_v
    port map (
            O => \N__19028\,
            I => \N__18982\
        );

    \I__4170\ : LocalMux
    port map (
            O => \N__19025\,
            I => \N__18979\
        );

    \I__4169\ : InMux
    port map (
            O => \N__19024\,
            I => \N__18976\
        );

    \I__4168\ : InMux
    port map (
            O => \N__19023\,
            I => \N__18971\
        );

    \I__4167\ : InMux
    port map (
            O => \N__19022\,
            I => \N__18971\
        );

    \I__4166\ : LocalMux
    port map (
            O => \N__19019\,
            I => \N__18966\
        );

    \I__4165\ : LocalMux
    port map (
            O => \N__19014\,
            I => \N__18966\
        );

    \I__4164\ : LocalMux
    port map (
            O => \N__19011\,
            I => \N__18957\
        );

    \I__4163\ : Span4Mux_h
    port map (
            O => \N__19008\,
            I => \N__18957\
        );

    \I__4162\ : LocalMux
    port map (
            O => \N__19003\,
            I => \N__18957\
        );

    \I__4161\ : Span4Mux_v
    port map (
            O => \N__18998\,
            I => \N__18957\
        );

    \I__4160\ : Span4Mux_v
    port map (
            O => \N__18993\,
            I => \N__18954\
        );

    \I__4159\ : Span4Mux_h
    port map (
            O => \N__18990\,
            I => \N__18951\
        );

    \I__4158\ : InMux
    port map (
            O => \N__18989\,
            I => \N__18948\
        );

    \I__4157\ : InMux
    port map (
            O => \N__18988\,
            I => \N__18943\
        );

    \I__4156\ : InMux
    port map (
            O => \N__18987\,
            I => \N__18943\
        );

    \I__4155\ : Span4Mux_v
    port map (
            O => \N__18982\,
            I => \N__18940\
        );

    \I__4154\ : Span4Mux_v
    port map (
            O => \N__18979\,
            I => \N__18929\
        );

    \I__4153\ : LocalMux
    port map (
            O => \N__18976\,
            I => \N__18929\
        );

    \I__4152\ : LocalMux
    port map (
            O => \N__18971\,
            I => \N__18929\
        );

    \I__4151\ : Span4Mux_h
    port map (
            O => \N__18966\,
            I => \N__18929\
        );

    \I__4150\ : Span4Mux_v
    port map (
            O => \N__18957\,
            I => \N__18929\
        );

    \I__4149\ : Odrv4
    port map (
            O => \N__18954\,
            I => \transmit_module.n3787\
        );

    \I__4148\ : Odrv4
    port map (
            O => \N__18951\,
            I => \transmit_module.n3787\
        );

    \I__4147\ : LocalMux
    port map (
            O => \N__18948\,
            I => \transmit_module.n3787\
        );

    \I__4146\ : LocalMux
    port map (
            O => \N__18943\,
            I => \transmit_module.n3787\
        );

    \I__4145\ : Odrv4
    port map (
            O => \N__18940\,
            I => \transmit_module.n3787\
        );

    \I__4144\ : Odrv4
    port map (
            O => \N__18929\,
            I => \transmit_module.n3787\
        );

    \I__4143\ : InMux
    port map (
            O => \N__18916\,
            I => \N__18913\
        );

    \I__4142\ : LocalMux
    port map (
            O => \N__18913\,
            I => \N__18909\
        );

    \I__4141\ : InMux
    port map (
            O => \N__18912\,
            I => \N__18906\
        );

    \I__4140\ : Span12Mux_v
    port map (
            O => \N__18909\,
            I => \N__18903\
        );

    \I__4139\ : LocalMux
    port map (
            O => \N__18906\,
            I => \transmit_module.n108\
        );

    \I__4138\ : Odrv12
    port map (
            O => \N__18903\,
            I => \transmit_module.n108\
        );

    \I__4137\ : InMux
    port map (
            O => \N__18898\,
            I => \N__18895\
        );

    \I__4136\ : LocalMux
    port map (
            O => \N__18895\,
            I => \N__18892\
        );

    \I__4135\ : Odrv12
    port map (
            O => \N__18892\,
            I => \transmit_module.n139\
        );

    \I__4134\ : CascadeMux
    port map (
            O => \N__18889\,
            I => \N__18886\
        );

    \I__4133\ : CascadeBuf
    port map (
            O => \N__18886\,
            I => \N__18882\
        );

    \I__4132\ : CascadeMux
    port map (
            O => \N__18885\,
            I => \N__18879\
        );

    \I__4131\ : CascadeMux
    port map (
            O => \N__18882\,
            I => \N__18876\
        );

    \I__4130\ : CascadeBuf
    port map (
            O => \N__18879\,
            I => \N__18873\
        );

    \I__4129\ : CascadeBuf
    port map (
            O => \N__18876\,
            I => \N__18870\
        );

    \I__4128\ : CascadeMux
    port map (
            O => \N__18873\,
            I => \N__18867\
        );

    \I__4127\ : CascadeMux
    port map (
            O => \N__18870\,
            I => \N__18864\
        );

    \I__4126\ : CascadeBuf
    port map (
            O => \N__18867\,
            I => \N__18861\
        );

    \I__4125\ : CascadeBuf
    port map (
            O => \N__18864\,
            I => \N__18858\
        );

    \I__4124\ : CascadeMux
    port map (
            O => \N__18861\,
            I => \N__18855\
        );

    \I__4123\ : CascadeMux
    port map (
            O => \N__18858\,
            I => \N__18852\
        );

    \I__4122\ : CascadeBuf
    port map (
            O => \N__18855\,
            I => \N__18849\
        );

    \I__4121\ : CascadeBuf
    port map (
            O => \N__18852\,
            I => \N__18846\
        );

    \I__4120\ : CascadeMux
    port map (
            O => \N__18849\,
            I => \N__18843\
        );

    \I__4119\ : CascadeMux
    port map (
            O => \N__18846\,
            I => \N__18840\
        );

    \I__4118\ : CascadeBuf
    port map (
            O => \N__18843\,
            I => \N__18837\
        );

    \I__4117\ : CascadeBuf
    port map (
            O => \N__18840\,
            I => \N__18834\
        );

    \I__4116\ : CascadeMux
    port map (
            O => \N__18837\,
            I => \N__18831\
        );

    \I__4115\ : CascadeMux
    port map (
            O => \N__18834\,
            I => \N__18828\
        );

    \I__4114\ : CascadeBuf
    port map (
            O => \N__18831\,
            I => \N__18825\
        );

    \I__4113\ : CascadeBuf
    port map (
            O => \N__18828\,
            I => \N__18822\
        );

    \I__4112\ : CascadeMux
    port map (
            O => \N__18825\,
            I => \N__18819\
        );

    \I__4111\ : CascadeMux
    port map (
            O => \N__18822\,
            I => \N__18816\
        );

    \I__4110\ : CascadeBuf
    port map (
            O => \N__18819\,
            I => \N__18813\
        );

    \I__4109\ : CascadeBuf
    port map (
            O => \N__18816\,
            I => \N__18810\
        );

    \I__4108\ : CascadeMux
    port map (
            O => \N__18813\,
            I => \N__18807\
        );

    \I__4107\ : CascadeMux
    port map (
            O => \N__18810\,
            I => \N__18804\
        );

    \I__4106\ : CascadeBuf
    port map (
            O => \N__18807\,
            I => \N__18801\
        );

    \I__4105\ : CascadeBuf
    port map (
            O => \N__18804\,
            I => \N__18798\
        );

    \I__4104\ : CascadeMux
    port map (
            O => \N__18801\,
            I => \N__18795\
        );

    \I__4103\ : CascadeMux
    port map (
            O => \N__18798\,
            I => \N__18792\
        );

    \I__4102\ : CascadeBuf
    port map (
            O => \N__18795\,
            I => \N__18789\
        );

    \I__4101\ : CascadeBuf
    port map (
            O => \N__18792\,
            I => \N__18786\
        );

    \I__4100\ : CascadeMux
    port map (
            O => \N__18789\,
            I => \N__18783\
        );

    \I__4099\ : CascadeMux
    port map (
            O => \N__18786\,
            I => \N__18780\
        );

    \I__4098\ : CascadeBuf
    port map (
            O => \N__18783\,
            I => \N__18777\
        );

    \I__4097\ : CascadeBuf
    port map (
            O => \N__18780\,
            I => \N__18774\
        );

    \I__4096\ : CascadeMux
    port map (
            O => \N__18777\,
            I => \N__18771\
        );

    \I__4095\ : CascadeMux
    port map (
            O => \N__18774\,
            I => \N__18768\
        );

    \I__4094\ : CascadeBuf
    port map (
            O => \N__18771\,
            I => \N__18765\
        );

    \I__4093\ : CascadeBuf
    port map (
            O => \N__18768\,
            I => \N__18762\
        );

    \I__4092\ : CascadeMux
    port map (
            O => \N__18765\,
            I => \N__18759\
        );

    \I__4091\ : CascadeMux
    port map (
            O => \N__18762\,
            I => \N__18756\
        );

    \I__4090\ : CascadeBuf
    port map (
            O => \N__18759\,
            I => \N__18753\
        );

    \I__4089\ : CascadeBuf
    port map (
            O => \N__18756\,
            I => \N__18750\
        );

    \I__4088\ : CascadeMux
    port map (
            O => \N__18753\,
            I => \N__18747\
        );

    \I__4087\ : CascadeMux
    port map (
            O => \N__18750\,
            I => \N__18744\
        );

    \I__4086\ : CascadeBuf
    port map (
            O => \N__18747\,
            I => \N__18741\
        );

    \I__4085\ : CascadeBuf
    port map (
            O => \N__18744\,
            I => \N__18738\
        );

    \I__4084\ : CascadeMux
    port map (
            O => \N__18741\,
            I => \N__18735\
        );

    \I__4083\ : CascadeMux
    port map (
            O => \N__18738\,
            I => \N__18732\
        );

    \I__4082\ : CascadeBuf
    port map (
            O => \N__18735\,
            I => \N__18729\
        );

    \I__4081\ : CascadeBuf
    port map (
            O => \N__18732\,
            I => \N__18726\
        );

    \I__4080\ : CascadeMux
    port map (
            O => \N__18729\,
            I => \N__18723\
        );

    \I__4079\ : CascadeMux
    port map (
            O => \N__18726\,
            I => \N__18720\
        );

    \I__4078\ : CascadeBuf
    port map (
            O => \N__18723\,
            I => \N__18717\
        );

    \I__4077\ : CascadeBuf
    port map (
            O => \N__18720\,
            I => \N__18714\
        );

    \I__4076\ : CascadeMux
    port map (
            O => \N__18717\,
            I => \N__18711\
        );

    \I__4075\ : CascadeMux
    port map (
            O => \N__18714\,
            I => \N__18708\
        );

    \I__4074\ : CascadeBuf
    port map (
            O => \N__18711\,
            I => \N__18705\
        );

    \I__4073\ : InMux
    port map (
            O => \N__18708\,
            I => \N__18702\
        );

    \I__4072\ : CascadeMux
    port map (
            O => \N__18705\,
            I => \N__18699\
        );

    \I__4071\ : LocalMux
    port map (
            O => \N__18702\,
            I => \N__18696\
        );

    \I__4070\ : InMux
    port map (
            O => \N__18699\,
            I => \N__18693\
        );

    \I__4069\ : Span4Mux_s3_v
    port map (
            O => \N__18696\,
            I => \N__18690\
        );

    \I__4068\ : LocalMux
    port map (
            O => \N__18693\,
            I => \N__18687\
        );

    \I__4067\ : Span4Mux_v
    port map (
            O => \N__18690\,
            I => \N__18684\
        );

    \I__4066\ : Span4Mux_h
    port map (
            O => \N__18687\,
            I => \N__18681\
        );

    \I__4065\ : Span4Mux_h
    port map (
            O => \N__18684\,
            I => \N__18678\
        );

    \I__4064\ : Span4Mux_h
    port map (
            O => \N__18681\,
            I => \N__18675\
        );

    \I__4063\ : Span4Mux_h
    port map (
            O => \N__18678\,
            I => \N__18672\
        );

    \I__4062\ : Sp12to4
    port map (
            O => \N__18675\,
            I => \N__18669\
        );

    \I__4061\ : Odrv4
    port map (
            O => \N__18672\,
            I => n20
        );

    \I__4060\ : Odrv12
    port map (
            O => \N__18669\,
            I => n20
        );

    \I__4059\ : IoInMux
    port map (
            O => \N__18664\,
            I => \N__18661\
        );

    \I__4058\ : LocalMux
    port map (
            O => \N__18661\,
            I => \N__18658\
        );

    \I__4057\ : Span4Mux_s0_v
    port map (
            O => \N__18658\,
            I => \N__18655\
        );

    \I__4056\ : Odrv4
    port map (
            O => \N__18655\,
            I => \GB_BUFFER_TVP_CLK_c_THRU_CO\
        );

    \I__4055\ : InMux
    port map (
            O => \N__18652\,
            I => \N__18646\
        );

    \I__4054\ : InMux
    port map (
            O => \N__18651\,
            I => \N__18646\
        );

    \I__4053\ : LocalMux
    port map (
            O => \N__18646\,
            I => \N__18642\
        );

    \I__4052\ : InMux
    port map (
            O => \N__18645\,
            I => \N__18639\
        );

    \I__4051\ : Span4Mux_v
    port map (
            O => \N__18642\,
            I => \N__18636\
        );

    \I__4050\ : LocalMux
    port map (
            O => \N__18639\,
            I => \N__18633\
        );

    \I__4049\ : Span4Mux_h
    port map (
            O => \N__18636\,
            I => \N__18628\
        );

    \I__4048\ : Span4Mux_h
    port map (
            O => \N__18633\,
            I => \N__18628\
        );

    \I__4047\ : Sp12to4
    port map (
            O => \N__18628\,
            I => \N__18625\
        );

    \I__4046\ : Odrv12
    port map (
            O => \N__18625\,
            I => \TVP_HSYNC_c\
        );

    \I__4045\ : InMux
    port map (
            O => \N__18622\,
            I => \N__18619\
        );

    \I__4044\ : LocalMux
    port map (
            O => \N__18619\,
            I => \receive_module.rx_counter.n10\
        );

    \I__4043\ : InMux
    port map (
            O => \N__18616\,
            I => \bfn_17_10_0_\
        );

    \I__4042\ : InMux
    port map (
            O => \N__18613\,
            I => \N__18610\
        );

    \I__4041\ : LocalMux
    port map (
            O => \N__18610\,
            I => \receive_module.rx_counter.n9\
        );

    \I__4040\ : InMux
    port map (
            O => \N__18607\,
            I => \receive_module.rx_counter.n3301\
        );

    \I__4039\ : InMux
    port map (
            O => \N__18604\,
            I => \N__18601\
        );

    \I__4038\ : LocalMux
    port map (
            O => \N__18601\,
            I => \receive_module.rx_counter.n8\
        );

    \I__4037\ : InMux
    port map (
            O => \N__18598\,
            I => \receive_module.rx_counter.n3302\
        );

    \I__4036\ : InMux
    port map (
            O => \N__18595\,
            I => \N__18590\
        );

    \I__4035\ : InMux
    port map (
            O => \N__18594\,
            I => \N__18585\
        );

    \I__4034\ : InMux
    port map (
            O => \N__18593\,
            I => \N__18585\
        );

    \I__4033\ : LocalMux
    port map (
            O => \N__18590\,
            I => \receive_module.rx_counter.X_3\
        );

    \I__4032\ : LocalMux
    port map (
            O => \N__18585\,
            I => \receive_module.rx_counter.X_3\
        );

    \I__4031\ : InMux
    port map (
            O => \N__18580\,
            I => \receive_module.rx_counter.n3303\
        );

    \I__4030\ : InMux
    port map (
            O => \N__18577\,
            I => \N__18574\
        );

    \I__4029\ : LocalMux
    port map (
            O => \N__18574\,
            I => \N__18571\
        );

    \I__4028\ : Span4Mux_h
    port map (
            O => \N__18571\,
            I => \N__18568\
        );

    \I__4027\ : Span4Mux_v
    port map (
            O => \N__18568\,
            I => \N__18564\
        );

    \I__4026\ : InMux
    port map (
            O => \N__18567\,
            I => \N__18561\
        );

    \I__4025\ : Odrv4
    port map (
            O => \N__18564\,
            I => \transmit_module.n114\
        );

    \I__4024\ : LocalMux
    port map (
            O => \N__18561\,
            I => \transmit_module.n114\
        );

    \I__4023\ : InMux
    port map (
            O => \N__18556\,
            I => \N__18553\
        );

    \I__4022\ : LocalMux
    port map (
            O => \N__18553\,
            I => \N__18550\
        );

    \I__4021\ : Span4Mux_h
    port map (
            O => \N__18550\,
            I => \N__18546\
        );

    \I__4020\ : InMux
    port map (
            O => \N__18549\,
            I => \N__18543\
        );

    \I__4019\ : Odrv4
    port map (
            O => \N__18546\,
            I => \transmit_module.n145\
        );

    \I__4018\ : LocalMux
    port map (
            O => \N__18543\,
            I => \transmit_module.n145\
        );

    \I__4017\ : CascadeMux
    port map (
            O => \N__18538\,
            I => \N__18535\
        );

    \I__4016\ : CascadeBuf
    port map (
            O => \N__18535\,
            I => \N__18531\
        );

    \I__4015\ : CascadeMux
    port map (
            O => \N__18534\,
            I => \N__18528\
        );

    \I__4014\ : CascadeMux
    port map (
            O => \N__18531\,
            I => \N__18525\
        );

    \I__4013\ : CascadeBuf
    port map (
            O => \N__18528\,
            I => \N__18522\
        );

    \I__4012\ : CascadeBuf
    port map (
            O => \N__18525\,
            I => \N__18519\
        );

    \I__4011\ : CascadeMux
    port map (
            O => \N__18522\,
            I => \N__18516\
        );

    \I__4010\ : CascadeMux
    port map (
            O => \N__18519\,
            I => \N__18513\
        );

    \I__4009\ : CascadeBuf
    port map (
            O => \N__18516\,
            I => \N__18510\
        );

    \I__4008\ : CascadeBuf
    port map (
            O => \N__18513\,
            I => \N__18507\
        );

    \I__4007\ : CascadeMux
    port map (
            O => \N__18510\,
            I => \N__18504\
        );

    \I__4006\ : CascadeMux
    port map (
            O => \N__18507\,
            I => \N__18501\
        );

    \I__4005\ : CascadeBuf
    port map (
            O => \N__18504\,
            I => \N__18498\
        );

    \I__4004\ : CascadeBuf
    port map (
            O => \N__18501\,
            I => \N__18495\
        );

    \I__4003\ : CascadeMux
    port map (
            O => \N__18498\,
            I => \N__18492\
        );

    \I__4002\ : CascadeMux
    port map (
            O => \N__18495\,
            I => \N__18489\
        );

    \I__4001\ : CascadeBuf
    port map (
            O => \N__18492\,
            I => \N__18486\
        );

    \I__4000\ : CascadeBuf
    port map (
            O => \N__18489\,
            I => \N__18483\
        );

    \I__3999\ : CascadeMux
    port map (
            O => \N__18486\,
            I => \N__18480\
        );

    \I__3998\ : CascadeMux
    port map (
            O => \N__18483\,
            I => \N__18477\
        );

    \I__3997\ : CascadeBuf
    port map (
            O => \N__18480\,
            I => \N__18474\
        );

    \I__3996\ : CascadeBuf
    port map (
            O => \N__18477\,
            I => \N__18471\
        );

    \I__3995\ : CascadeMux
    port map (
            O => \N__18474\,
            I => \N__18468\
        );

    \I__3994\ : CascadeMux
    port map (
            O => \N__18471\,
            I => \N__18465\
        );

    \I__3993\ : CascadeBuf
    port map (
            O => \N__18468\,
            I => \N__18462\
        );

    \I__3992\ : CascadeBuf
    port map (
            O => \N__18465\,
            I => \N__18459\
        );

    \I__3991\ : CascadeMux
    port map (
            O => \N__18462\,
            I => \N__18456\
        );

    \I__3990\ : CascadeMux
    port map (
            O => \N__18459\,
            I => \N__18453\
        );

    \I__3989\ : CascadeBuf
    port map (
            O => \N__18456\,
            I => \N__18450\
        );

    \I__3988\ : CascadeBuf
    port map (
            O => \N__18453\,
            I => \N__18447\
        );

    \I__3987\ : CascadeMux
    port map (
            O => \N__18450\,
            I => \N__18444\
        );

    \I__3986\ : CascadeMux
    port map (
            O => \N__18447\,
            I => \N__18441\
        );

    \I__3985\ : CascadeBuf
    port map (
            O => \N__18444\,
            I => \N__18438\
        );

    \I__3984\ : CascadeBuf
    port map (
            O => \N__18441\,
            I => \N__18435\
        );

    \I__3983\ : CascadeMux
    port map (
            O => \N__18438\,
            I => \N__18432\
        );

    \I__3982\ : CascadeMux
    port map (
            O => \N__18435\,
            I => \N__18429\
        );

    \I__3981\ : CascadeBuf
    port map (
            O => \N__18432\,
            I => \N__18426\
        );

    \I__3980\ : CascadeBuf
    port map (
            O => \N__18429\,
            I => \N__18423\
        );

    \I__3979\ : CascadeMux
    port map (
            O => \N__18426\,
            I => \N__18420\
        );

    \I__3978\ : CascadeMux
    port map (
            O => \N__18423\,
            I => \N__18417\
        );

    \I__3977\ : CascadeBuf
    port map (
            O => \N__18420\,
            I => \N__18414\
        );

    \I__3976\ : CascadeBuf
    port map (
            O => \N__18417\,
            I => \N__18411\
        );

    \I__3975\ : CascadeMux
    port map (
            O => \N__18414\,
            I => \N__18408\
        );

    \I__3974\ : CascadeMux
    port map (
            O => \N__18411\,
            I => \N__18405\
        );

    \I__3973\ : CascadeBuf
    port map (
            O => \N__18408\,
            I => \N__18402\
        );

    \I__3972\ : CascadeBuf
    port map (
            O => \N__18405\,
            I => \N__18399\
        );

    \I__3971\ : CascadeMux
    port map (
            O => \N__18402\,
            I => \N__18396\
        );

    \I__3970\ : CascadeMux
    port map (
            O => \N__18399\,
            I => \N__18393\
        );

    \I__3969\ : CascadeBuf
    port map (
            O => \N__18396\,
            I => \N__18390\
        );

    \I__3968\ : CascadeBuf
    port map (
            O => \N__18393\,
            I => \N__18387\
        );

    \I__3967\ : CascadeMux
    port map (
            O => \N__18390\,
            I => \N__18384\
        );

    \I__3966\ : CascadeMux
    port map (
            O => \N__18387\,
            I => \N__18381\
        );

    \I__3965\ : CascadeBuf
    port map (
            O => \N__18384\,
            I => \N__18378\
        );

    \I__3964\ : CascadeBuf
    port map (
            O => \N__18381\,
            I => \N__18375\
        );

    \I__3963\ : CascadeMux
    port map (
            O => \N__18378\,
            I => \N__18372\
        );

    \I__3962\ : CascadeMux
    port map (
            O => \N__18375\,
            I => \N__18369\
        );

    \I__3961\ : CascadeBuf
    port map (
            O => \N__18372\,
            I => \N__18366\
        );

    \I__3960\ : CascadeBuf
    port map (
            O => \N__18369\,
            I => \N__18363\
        );

    \I__3959\ : CascadeMux
    port map (
            O => \N__18366\,
            I => \N__18360\
        );

    \I__3958\ : CascadeMux
    port map (
            O => \N__18363\,
            I => \N__18357\
        );

    \I__3957\ : CascadeBuf
    port map (
            O => \N__18360\,
            I => \N__18354\
        );

    \I__3956\ : InMux
    port map (
            O => \N__18357\,
            I => \N__18351\
        );

    \I__3955\ : CascadeMux
    port map (
            O => \N__18354\,
            I => \N__18348\
        );

    \I__3954\ : LocalMux
    port map (
            O => \N__18351\,
            I => \N__18345\
        );

    \I__3953\ : InMux
    port map (
            O => \N__18348\,
            I => \N__18342\
        );

    \I__3952\ : Span4Mux_v
    port map (
            O => \N__18345\,
            I => \N__18339\
        );

    \I__3951\ : LocalMux
    port map (
            O => \N__18342\,
            I => \N__18336\
        );

    \I__3950\ : Span4Mux_v
    port map (
            O => \N__18339\,
            I => \N__18333\
        );

    \I__3949\ : Span4Mux_h
    port map (
            O => \N__18336\,
            I => \N__18330\
        );

    \I__3948\ : Span4Mux_v
    port map (
            O => \N__18333\,
            I => \N__18327\
        );

    \I__3947\ : Sp12to4
    port map (
            O => \N__18330\,
            I => \N__18324\
        );

    \I__3946\ : Sp12to4
    port map (
            O => \N__18327\,
            I => \N__18319\
        );

    \I__3945\ : Span12Mux_v
    port map (
            O => \N__18324\,
            I => \N__18319\
        );

    \I__3944\ : Odrv12
    port map (
            O => \N__18319\,
            I => n26
        );

    \I__3943\ : InMux
    port map (
            O => \N__18316\,
            I => \N__18311\
        );

    \I__3942\ : InMux
    port map (
            O => \N__18315\,
            I => \N__18308\
        );

    \I__3941\ : InMux
    port map (
            O => \N__18314\,
            I => \N__18304\
        );

    \I__3940\ : LocalMux
    port map (
            O => \N__18311\,
            I => \N__18295\
        );

    \I__3939\ : LocalMux
    port map (
            O => \N__18308\,
            I => \N__18291\
        );

    \I__3938\ : InMux
    port map (
            O => \N__18307\,
            I => \N__18288\
        );

    \I__3937\ : LocalMux
    port map (
            O => \N__18304\,
            I => \N__18285\
        );

    \I__3936\ : InMux
    port map (
            O => \N__18303\,
            I => \N__18280\
        );

    \I__3935\ : InMux
    port map (
            O => \N__18302\,
            I => \N__18280\
        );

    \I__3934\ : InMux
    port map (
            O => \N__18301\,
            I => \N__18275\
        );

    \I__3933\ : InMux
    port map (
            O => \N__18300\,
            I => \N__18275\
        );

    \I__3932\ : CascadeMux
    port map (
            O => \N__18299\,
            I => \N__18270\
        );

    \I__3931\ : InMux
    port map (
            O => \N__18298\,
            I => \N__18266\
        );

    \I__3930\ : Span12Mux_h
    port map (
            O => \N__18295\,
            I => \N__18263\
        );

    \I__3929\ : InMux
    port map (
            O => \N__18294\,
            I => \N__18260\
        );

    \I__3928\ : Span4Mux_h
    port map (
            O => \N__18291\,
            I => \N__18257\
        );

    \I__3927\ : LocalMux
    port map (
            O => \N__18288\,
            I => \N__18250\
        );

    \I__3926\ : Span4Mux_v
    port map (
            O => \N__18285\,
            I => \N__18250\
        );

    \I__3925\ : LocalMux
    port map (
            O => \N__18280\,
            I => \N__18250\
        );

    \I__3924\ : LocalMux
    port map (
            O => \N__18275\,
            I => \N__18247\
        );

    \I__3923\ : InMux
    port map (
            O => \N__18274\,
            I => \N__18242\
        );

    \I__3922\ : InMux
    port map (
            O => \N__18273\,
            I => \N__18242\
        );

    \I__3921\ : InMux
    port map (
            O => \N__18270\,
            I => \N__18237\
        );

    \I__3920\ : InMux
    port map (
            O => \N__18269\,
            I => \N__18237\
        );

    \I__3919\ : LocalMux
    port map (
            O => \N__18266\,
            I => \transmit_module.VGA_VISIBLE\
        );

    \I__3918\ : Odrv12
    port map (
            O => \N__18263\,
            I => \transmit_module.VGA_VISIBLE\
        );

    \I__3917\ : LocalMux
    port map (
            O => \N__18260\,
            I => \transmit_module.VGA_VISIBLE\
        );

    \I__3916\ : Odrv4
    port map (
            O => \N__18257\,
            I => \transmit_module.VGA_VISIBLE\
        );

    \I__3915\ : Odrv4
    port map (
            O => \N__18250\,
            I => \transmit_module.VGA_VISIBLE\
        );

    \I__3914\ : Odrv4
    port map (
            O => \N__18247\,
            I => \transmit_module.VGA_VISIBLE\
        );

    \I__3913\ : LocalMux
    port map (
            O => \N__18242\,
            I => \transmit_module.VGA_VISIBLE\
        );

    \I__3912\ : LocalMux
    port map (
            O => \N__18237\,
            I => \transmit_module.VGA_VISIBLE\
        );

    \I__3911\ : InMux
    port map (
            O => \N__18220\,
            I => \N__18217\
        );

    \I__3910\ : LocalMux
    port map (
            O => \N__18217\,
            I => \N__18214\
        );

    \I__3909\ : Span4Mux_v
    port map (
            O => \N__18214\,
            I => \N__18211\
        );

    \I__3908\ : Odrv4
    port map (
            O => \N__18211\,
            I => \transmit_module.n129\
        );

    \I__3907\ : InMux
    port map (
            O => \N__18208\,
            I => \N__18205\
        );

    \I__3906\ : LocalMux
    port map (
            O => \N__18205\,
            I => \N__18202\
        );

    \I__3905\ : Span4Mux_v
    port map (
            O => \N__18202\,
            I => \N__18199\
        );

    \I__3904\ : Odrv4
    port map (
            O => \N__18199\,
            I => \transmit_module.n144\
        );

    \I__3903\ : CascadeMux
    port map (
            O => \N__18196\,
            I => \transmit_module.n144_cascade_\
        );

    \I__3902\ : CascadeMux
    port map (
            O => \N__18193\,
            I => \N__18189\
        );

    \I__3901\ : CascadeMux
    port map (
            O => \N__18192\,
            I => \N__18186\
        );

    \I__3900\ : CascadeBuf
    port map (
            O => \N__18189\,
            I => \N__18183\
        );

    \I__3899\ : CascadeBuf
    port map (
            O => \N__18186\,
            I => \N__18180\
        );

    \I__3898\ : CascadeMux
    port map (
            O => \N__18183\,
            I => \N__18177\
        );

    \I__3897\ : CascadeMux
    port map (
            O => \N__18180\,
            I => \N__18174\
        );

    \I__3896\ : CascadeBuf
    port map (
            O => \N__18177\,
            I => \N__18171\
        );

    \I__3895\ : CascadeBuf
    port map (
            O => \N__18174\,
            I => \N__18168\
        );

    \I__3894\ : CascadeMux
    port map (
            O => \N__18171\,
            I => \N__18165\
        );

    \I__3893\ : CascadeMux
    port map (
            O => \N__18168\,
            I => \N__18162\
        );

    \I__3892\ : CascadeBuf
    port map (
            O => \N__18165\,
            I => \N__18159\
        );

    \I__3891\ : CascadeBuf
    port map (
            O => \N__18162\,
            I => \N__18156\
        );

    \I__3890\ : CascadeMux
    port map (
            O => \N__18159\,
            I => \N__18153\
        );

    \I__3889\ : CascadeMux
    port map (
            O => \N__18156\,
            I => \N__18150\
        );

    \I__3888\ : CascadeBuf
    port map (
            O => \N__18153\,
            I => \N__18147\
        );

    \I__3887\ : CascadeBuf
    port map (
            O => \N__18150\,
            I => \N__18144\
        );

    \I__3886\ : CascadeMux
    port map (
            O => \N__18147\,
            I => \N__18141\
        );

    \I__3885\ : CascadeMux
    port map (
            O => \N__18144\,
            I => \N__18138\
        );

    \I__3884\ : CascadeBuf
    port map (
            O => \N__18141\,
            I => \N__18135\
        );

    \I__3883\ : CascadeBuf
    port map (
            O => \N__18138\,
            I => \N__18132\
        );

    \I__3882\ : CascadeMux
    port map (
            O => \N__18135\,
            I => \N__18129\
        );

    \I__3881\ : CascadeMux
    port map (
            O => \N__18132\,
            I => \N__18126\
        );

    \I__3880\ : CascadeBuf
    port map (
            O => \N__18129\,
            I => \N__18123\
        );

    \I__3879\ : CascadeBuf
    port map (
            O => \N__18126\,
            I => \N__18120\
        );

    \I__3878\ : CascadeMux
    port map (
            O => \N__18123\,
            I => \N__18117\
        );

    \I__3877\ : CascadeMux
    port map (
            O => \N__18120\,
            I => \N__18114\
        );

    \I__3876\ : CascadeBuf
    port map (
            O => \N__18117\,
            I => \N__18111\
        );

    \I__3875\ : CascadeBuf
    port map (
            O => \N__18114\,
            I => \N__18108\
        );

    \I__3874\ : CascadeMux
    port map (
            O => \N__18111\,
            I => \N__18105\
        );

    \I__3873\ : CascadeMux
    port map (
            O => \N__18108\,
            I => \N__18102\
        );

    \I__3872\ : CascadeBuf
    port map (
            O => \N__18105\,
            I => \N__18099\
        );

    \I__3871\ : CascadeBuf
    port map (
            O => \N__18102\,
            I => \N__18096\
        );

    \I__3870\ : CascadeMux
    port map (
            O => \N__18099\,
            I => \N__18093\
        );

    \I__3869\ : CascadeMux
    port map (
            O => \N__18096\,
            I => \N__18090\
        );

    \I__3868\ : CascadeBuf
    port map (
            O => \N__18093\,
            I => \N__18087\
        );

    \I__3867\ : CascadeBuf
    port map (
            O => \N__18090\,
            I => \N__18084\
        );

    \I__3866\ : CascadeMux
    port map (
            O => \N__18087\,
            I => \N__18081\
        );

    \I__3865\ : CascadeMux
    port map (
            O => \N__18084\,
            I => \N__18078\
        );

    \I__3864\ : CascadeBuf
    port map (
            O => \N__18081\,
            I => \N__18075\
        );

    \I__3863\ : CascadeBuf
    port map (
            O => \N__18078\,
            I => \N__18072\
        );

    \I__3862\ : CascadeMux
    port map (
            O => \N__18075\,
            I => \N__18069\
        );

    \I__3861\ : CascadeMux
    port map (
            O => \N__18072\,
            I => \N__18066\
        );

    \I__3860\ : CascadeBuf
    port map (
            O => \N__18069\,
            I => \N__18063\
        );

    \I__3859\ : CascadeBuf
    port map (
            O => \N__18066\,
            I => \N__18060\
        );

    \I__3858\ : CascadeMux
    port map (
            O => \N__18063\,
            I => \N__18057\
        );

    \I__3857\ : CascadeMux
    port map (
            O => \N__18060\,
            I => \N__18054\
        );

    \I__3856\ : CascadeBuf
    port map (
            O => \N__18057\,
            I => \N__18051\
        );

    \I__3855\ : CascadeBuf
    port map (
            O => \N__18054\,
            I => \N__18048\
        );

    \I__3854\ : CascadeMux
    port map (
            O => \N__18051\,
            I => \N__18045\
        );

    \I__3853\ : CascadeMux
    port map (
            O => \N__18048\,
            I => \N__18042\
        );

    \I__3852\ : CascadeBuf
    port map (
            O => \N__18045\,
            I => \N__18039\
        );

    \I__3851\ : CascadeBuf
    port map (
            O => \N__18042\,
            I => \N__18036\
        );

    \I__3850\ : CascadeMux
    port map (
            O => \N__18039\,
            I => \N__18033\
        );

    \I__3849\ : CascadeMux
    port map (
            O => \N__18036\,
            I => \N__18030\
        );

    \I__3848\ : CascadeBuf
    port map (
            O => \N__18033\,
            I => \N__18027\
        );

    \I__3847\ : CascadeBuf
    port map (
            O => \N__18030\,
            I => \N__18024\
        );

    \I__3846\ : CascadeMux
    port map (
            O => \N__18027\,
            I => \N__18021\
        );

    \I__3845\ : CascadeMux
    port map (
            O => \N__18024\,
            I => \N__18018\
        );

    \I__3844\ : CascadeBuf
    port map (
            O => \N__18021\,
            I => \N__18015\
        );

    \I__3843\ : CascadeBuf
    port map (
            O => \N__18018\,
            I => \N__18012\
        );

    \I__3842\ : CascadeMux
    port map (
            O => \N__18015\,
            I => \N__18009\
        );

    \I__3841\ : CascadeMux
    port map (
            O => \N__18012\,
            I => \N__18006\
        );

    \I__3840\ : InMux
    port map (
            O => \N__18009\,
            I => \N__18003\
        );

    \I__3839\ : InMux
    port map (
            O => \N__18006\,
            I => \N__18000\
        );

    \I__3838\ : LocalMux
    port map (
            O => \N__18003\,
            I => \N__17997\
        );

    \I__3837\ : LocalMux
    port map (
            O => \N__18000\,
            I => \N__17994\
        );

    \I__3836\ : Span12Mux_s11_h
    port map (
            O => \N__17997\,
            I => \N__17991\
        );

    \I__3835\ : Sp12to4
    port map (
            O => \N__17994\,
            I => \N__17988\
        );

    \I__3834\ : Span12Mux_v
    port map (
            O => \N__17991\,
            I => \N__17983\
        );

    \I__3833\ : Span12Mux_v
    port map (
            O => \N__17988\,
            I => \N__17983\
        );

    \I__3832\ : Odrv12
    port map (
            O => \N__17983\,
            I => n25
        );

    \I__3831\ : InMux
    port map (
            O => \N__17980\,
            I => \N__17976\
        );

    \I__3830\ : InMux
    port map (
            O => \N__17979\,
            I => \N__17973\
        );

    \I__3829\ : LocalMux
    port map (
            O => \N__17976\,
            I => \N__17969\
        );

    \I__3828\ : LocalMux
    port map (
            O => \N__17973\,
            I => \N__17966\
        );

    \I__3827\ : InMux
    port map (
            O => \N__17972\,
            I => \N__17963\
        );

    \I__3826\ : Span4Mux_v
    port map (
            O => \N__17969\,
            I => \N__17956\
        );

    \I__3825\ : Span4Mux_h
    port map (
            O => \N__17966\,
            I => \N__17956\
        );

    \I__3824\ : LocalMux
    port map (
            O => \N__17963\,
            I => \N__17956\
        );

    \I__3823\ : Span4Mux_v
    port map (
            O => \N__17956\,
            I => \N__17952\
        );

    \I__3822\ : InMux
    port map (
            O => \N__17955\,
            I => \N__17949\
        );

    \I__3821\ : Odrv4
    port map (
            O => \N__17952\,
            I => \transmit_module.TX_ADDR_2\
        );

    \I__3820\ : LocalMux
    port map (
            O => \N__17949\,
            I => \transmit_module.TX_ADDR_2\
        );

    \I__3819\ : InMux
    port map (
            O => \N__17944\,
            I => \N__17941\
        );

    \I__3818\ : LocalMux
    port map (
            O => \N__17941\,
            I => \transmit_module.ADDR_Y_COMPONENT_2\
        );

    \I__3817\ : InMux
    port map (
            O => \N__17938\,
            I => \N__17934\
        );

    \I__3816\ : InMux
    port map (
            O => \N__17937\,
            I => \N__17930\
        );

    \I__3815\ : LocalMux
    port map (
            O => \N__17934\,
            I => \N__17924\
        );

    \I__3814\ : InMux
    port map (
            O => \N__17933\,
            I => \N__17921\
        );

    \I__3813\ : LocalMux
    port map (
            O => \N__17930\,
            I => \N__17918\
        );

    \I__3812\ : InMux
    port map (
            O => \N__17929\,
            I => \N__17915\
        );

    \I__3811\ : InMux
    port map (
            O => \N__17928\,
            I => \N__17912\
        );

    \I__3810\ : InMux
    port map (
            O => \N__17927\,
            I => \N__17909\
        );

    \I__3809\ : Span4Mux_h
    port map (
            O => \N__17924\,
            I => \N__17900\
        );

    \I__3808\ : LocalMux
    port map (
            O => \N__17921\,
            I => \N__17900\
        );

    \I__3807\ : Span4Mux_v
    port map (
            O => \N__17918\,
            I => \N__17897\
        );

    \I__3806\ : LocalMux
    port map (
            O => \N__17915\,
            I => \N__17894\
        );

    \I__3805\ : LocalMux
    port map (
            O => \N__17912\,
            I => \N__17891\
        );

    \I__3804\ : LocalMux
    port map (
            O => \N__17909\,
            I => \N__17888\
        );

    \I__3803\ : InMux
    port map (
            O => \N__17908\,
            I => \N__17885\
        );

    \I__3802\ : InMux
    port map (
            O => \N__17907\,
            I => \N__17878\
        );

    \I__3801\ : InMux
    port map (
            O => \N__17906\,
            I => \N__17875\
        );

    \I__3800\ : InMux
    port map (
            O => \N__17905\,
            I => \N__17872\
        );

    \I__3799\ : Span4Mux_v
    port map (
            O => \N__17900\,
            I => \N__17863\
        );

    \I__3798\ : Span4Mux_h
    port map (
            O => \N__17897\,
            I => \N__17863\
        );

    \I__3797\ : Span4Mux_v
    port map (
            O => \N__17894\,
            I => \N__17863\
        );

    \I__3796\ : Span4Mux_v
    port map (
            O => \N__17891\,
            I => \N__17863\
        );

    \I__3795\ : Sp12to4
    port map (
            O => \N__17888\,
            I => \N__17858\
        );

    \I__3794\ : LocalMux
    port map (
            O => \N__17885\,
            I => \N__17858\
        );

    \I__3793\ : InMux
    port map (
            O => \N__17884\,
            I => \N__17855\
        );

    \I__3792\ : InMux
    port map (
            O => \N__17883\,
            I => \N__17852\
        );

    \I__3791\ : InMux
    port map (
            O => \N__17882\,
            I => \N__17849\
        );

    \I__3790\ : InMux
    port map (
            O => \N__17881\,
            I => \N__17846\
        );

    \I__3789\ : LocalMux
    port map (
            O => \N__17878\,
            I => \transmit_module.Y_DELTA_PATTERN_0\
        );

    \I__3788\ : LocalMux
    port map (
            O => \N__17875\,
            I => \transmit_module.Y_DELTA_PATTERN_0\
        );

    \I__3787\ : LocalMux
    port map (
            O => \N__17872\,
            I => \transmit_module.Y_DELTA_PATTERN_0\
        );

    \I__3786\ : Odrv4
    port map (
            O => \N__17863\,
            I => \transmit_module.Y_DELTA_PATTERN_0\
        );

    \I__3785\ : Odrv12
    port map (
            O => \N__17858\,
            I => \transmit_module.Y_DELTA_PATTERN_0\
        );

    \I__3784\ : LocalMux
    port map (
            O => \N__17855\,
            I => \transmit_module.Y_DELTA_PATTERN_0\
        );

    \I__3783\ : LocalMux
    port map (
            O => \N__17852\,
            I => \transmit_module.Y_DELTA_PATTERN_0\
        );

    \I__3782\ : LocalMux
    port map (
            O => \N__17849\,
            I => \transmit_module.Y_DELTA_PATTERN_0\
        );

    \I__3781\ : LocalMux
    port map (
            O => \N__17846\,
            I => \transmit_module.Y_DELTA_PATTERN_0\
        );

    \I__3780\ : InMux
    port map (
            O => \N__17827\,
            I => \N__17824\
        );

    \I__3779\ : LocalMux
    port map (
            O => \N__17824\,
            I => \N__17821\
        );

    \I__3778\ : Span4Mux_v
    port map (
            O => \N__17821\,
            I => \N__17817\
        );

    \I__3777\ : InMux
    port map (
            O => \N__17820\,
            I => \N__17814\
        );

    \I__3776\ : Odrv4
    port map (
            O => \N__17817\,
            I => \transmit_module.n113\
        );

    \I__3775\ : LocalMux
    port map (
            O => \N__17814\,
            I => \transmit_module.n113\
        );

    \I__3774\ : InMux
    port map (
            O => \N__17809\,
            I => \N__17800\
        );

    \I__3773\ : InMux
    port map (
            O => \N__17808\,
            I => \N__17800\
        );

    \I__3772\ : InMux
    port map (
            O => \N__17807\,
            I => \N__17800\
        );

    \I__3771\ : LocalMux
    port map (
            O => \N__17800\,
            I => \N__17797\
        );

    \I__3770\ : Span4Mux_v
    port map (
            O => \N__17797\,
            I => \N__17793\
        );

    \I__3769\ : InMux
    port map (
            O => \N__17796\,
            I => \N__17790\
        );

    \I__3768\ : Odrv4
    port map (
            O => \N__17793\,
            I => \transmit_module.TX_ADDR_3\
        );

    \I__3767\ : LocalMux
    port map (
            O => \N__17790\,
            I => \transmit_module.TX_ADDR_3\
        );

    \I__3766\ : InMux
    port map (
            O => \N__17785\,
            I => \N__17782\
        );

    \I__3765\ : LocalMux
    port map (
            O => \N__17782\,
            I => \transmit_module.ADDR_Y_COMPONENT_3\
        );

    \I__3764\ : CEMux
    port map (
            O => \N__17779\,
            I => \N__17775\
        );

    \I__3763\ : CEMux
    port map (
            O => \N__17778\,
            I => \N__17771\
        );

    \I__3762\ : LocalMux
    port map (
            O => \N__17775\,
            I => \N__17767\
        );

    \I__3761\ : CEMux
    port map (
            O => \N__17774\,
            I => \N__17763\
        );

    \I__3760\ : LocalMux
    port map (
            O => \N__17771\,
            I => \N__17759\
        );

    \I__3759\ : CEMux
    port map (
            O => \N__17770\,
            I => \N__17756\
        );

    \I__3758\ : Span4Mux_v
    port map (
            O => \N__17767\,
            I => \N__17753\
        );

    \I__3757\ : CEMux
    port map (
            O => \N__17766\,
            I => \N__17750\
        );

    \I__3756\ : LocalMux
    port map (
            O => \N__17763\,
            I => \N__17747\
        );

    \I__3755\ : CEMux
    port map (
            O => \N__17762\,
            I => \N__17744\
        );

    \I__3754\ : Span4Mux_v
    port map (
            O => \N__17759\,
            I => \N__17738\
        );

    \I__3753\ : LocalMux
    port map (
            O => \N__17756\,
            I => \N__17738\
        );

    \I__3752\ : Span4Mux_h
    port map (
            O => \N__17753\,
            I => \N__17733\
        );

    \I__3751\ : LocalMux
    port map (
            O => \N__17750\,
            I => \N__17733\
        );

    \I__3750\ : Span4Mux_v
    port map (
            O => \N__17747\,
            I => \N__17728\
        );

    \I__3749\ : LocalMux
    port map (
            O => \N__17744\,
            I => \N__17728\
        );

    \I__3748\ : CEMux
    port map (
            O => \N__17743\,
            I => \N__17725\
        );

    \I__3747\ : Span4Mux_h
    port map (
            O => \N__17738\,
            I => \N__17720\
        );

    \I__3746\ : Span4Mux_h
    port map (
            O => \N__17733\,
            I => \N__17720\
        );

    \I__3745\ : Span4Mux_v
    port map (
            O => \N__17728\,
            I => \N__17717\
        );

    \I__3744\ : LocalMux
    port map (
            O => \N__17725\,
            I => \N__17714\
        );

    \I__3743\ : Odrv4
    port map (
            O => \N__17720\,
            I => \transmit_module.n2061\
        );

    \I__3742\ : Odrv4
    port map (
            O => \N__17717\,
            I => \transmit_module.n2061\
        );

    \I__3741\ : Odrv4
    port map (
            O => \N__17714\,
            I => \transmit_module.n2061\
        );

    \I__3740\ : InMux
    port map (
            O => \N__17707\,
            I => \N__17704\
        );

    \I__3739\ : LocalMux
    port map (
            O => \N__17704\,
            I => \N__17701\
        );

    \I__3738\ : Odrv4
    port map (
            O => \N__17701\,
            I => \TX_DATA_4\
        );

    \I__3737\ : IoInMux
    port map (
            O => \N__17698\,
            I => \N__17694\
        );

    \I__3736\ : IoInMux
    port map (
            O => \N__17697\,
            I => \N__17690\
        );

    \I__3735\ : LocalMux
    port map (
            O => \N__17694\,
            I => \N__17687\
        );

    \I__3734\ : IoInMux
    port map (
            O => \N__17693\,
            I => \N__17684\
        );

    \I__3733\ : LocalMux
    port map (
            O => \N__17690\,
            I => \N__17681\
        );

    \I__3732\ : IoSpan4Mux
    port map (
            O => \N__17687\,
            I => \N__17678\
        );

    \I__3731\ : LocalMux
    port map (
            O => \N__17684\,
            I => \N__17675\
        );

    \I__3730\ : IoSpan4Mux
    port map (
            O => \N__17681\,
            I => \N__17672\
        );

    \I__3729\ : Span4Mux_s3_h
    port map (
            O => \N__17678\,
            I => \N__17669\
        );

    \I__3728\ : Span4Mux_s2_v
    port map (
            O => \N__17675\,
            I => \N__17666\
        );

    \I__3727\ : Span4Mux_s2_v
    port map (
            O => \N__17672\,
            I => \N__17663\
        );

    \I__3726\ : Span4Mux_h
    port map (
            O => \N__17669\,
            I => \N__17660\
        );

    \I__3725\ : Sp12to4
    port map (
            O => \N__17666\,
            I => \N__17657\
        );

    \I__3724\ : Sp12to4
    port map (
            O => \N__17663\,
            I => \N__17654\
        );

    \I__3723\ : Span4Mux_h
    port map (
            O => \N__17660\,
            I => \N__17651\
        );

    \I__3722\ : Span12Mux_h
    port map (
            O => \N__17657\,
            I => \N__17646\
        );

    \I__3721\ : Span12Mux_h
    port map (
            O => \N__17654\,
            I => \N__17646\
        );

    \I__3720\ : Span4Mux_h
    port map (
            O => \N__17651\,
            I => \N__17643\
        );

    \I__3719\ : Odrv12
    port map (
            O => \N__17646\,
            I => n1794
        );

    \I__3718\ : Odrv4
    port map (
            O => \N__17643\,
            I => n1794
        );

    \I__3717\ : InMux
    port map (
            O => \N__17638\,
            I => \N__17635\
        );

    \I__3716\ : LocalMux
    port map (
            O => \N__17635\,
            I => \N__17632\
        );

    \I__3715\ : Odrv4
    port map (
            O => \N__17632\,
            I => \TX_DATA_2\
        );

    \I__3714\ : IoInMux
    port map (
            O => \N__17629\,
            I => \N__17625\
        );

    \I__3713\ : IoInMux
    port map (
            O => \N__17628\,
            I => \N__17621\
        );

    \I__3712\ : LocalMux
    port map (
            O => \N__17625\,
            I => \N__17618\
        );

    \I__3711\ : IoInMux
    port map (
            O => \N__17624\,
            I => \N__17615\
        );

    \I__3710\ : LocalMux
    port map (
            O => \N__17621\,
            I => \N__17612\
        );

    \I__3709\ : Span4Mux_s3_h
    port map (
            O => \N__17618\,
            I => \N__17609\
        );

    \I__3708\ : LocalMux
    port map (
            O => \N__17615\,
            I => \N__17606\
        );

    \I__3707\ : Span12Mux_s5_v
    port map (
            O => \N__17612\,
            I => \N__17601\
        );

    \I__3706\ : Sp12to4
    port map (
            O => \N__17609\,
            I => \N__17601\
        );

    \I__3705\ : IoSpan4Mux
    port map (
            O => \N__17606\,
            I => \N__17598\
        );

    \I__3704\ : Span12Mux_v
    port map (
            O => \N__17601\,
            I => \N__17595\
        );

    \I__3703\ : Sp12to4
    port map (
            O => \N__17598\,
            I => \N__17592\
        );

    \I__3702\ : Span12Mux_h
    port map (
            O => \N__17595\,
            I => \N__17589\
        );

    \I__3701\ : Span12Mux_v
    port map (
            O => \N__17592\,
            I => \N__17586\
        );

    \I__3700\ : Odrv12
    port map (
            O => \N__17589\,
            I => n1796
        );

    \I__3699\ : Odrv12
    port map (
            O => \N__17586\,
            I => n1796
        );

    \I__3698\ : InMux
    port map (
            O => \N__17581\,
            I => \N__17578\
        );

    \I__3697\ : LocalMux
    port map (
            O => \N__17578\,
            I => \transmit_module.ADDR_Y_COMPONENT_13\
        );

    \I__3696\ : InMux
    port map (
            O => \N__17575\,
            I => \N__17572\
        );

    \I__3695\ : LocalMux
    port map (
            O => \N__17572\,
            I => \N__17569\
        );

    \I__3694\ : Span12Mux_v
    port map (
            O => \N__17569\,
            I => \N__17566\
        );

    \I__3693\ : Odrv12
    port map (
            O => \N__17566\,
            I => \line_buffer.n3634\
        );

    \I__3692\ : InMux
    port map (
            O => \N__17563\,
            I => \N__17560\
        );

    \I__3691\ : LocalMux
    port map (
            O => \N__17560\,
            I => \N__17557\
        );

    \I__3690\ : Span4Mux_v
    port map (
            O => \N__17557\,
            I => \N__17554\
        );

    \I__3689\ : Span4Mux_h
    port map (
            O => \N__17554\,
            I => \N__17551\
        );

    \I__3688\ : Span4Mux_h
    port map (
            O => \N__17551\,
            I => \N__17548\
        );

    \I__3687\ : Odrv4
    port map (
            O => \N__17548\,
            I => \line_buffer.n442\
        );

    \I__3686\ : CascadeMux
    port map (
            O => \N__17545\,
            I => \N__17542\
        );

    \I__3685\ : InMux
    port map (
            O => \N__17542\,
            I => \N__17539\
        );

    \I__3684\ : LocalMux
    port map (
            O => \N__17539\,
            I => \N__17536\
        );

    \I__3683\ : Span4Mux_v
    port map (
            O => \N__17536\,
            I => \N__17533\
        );

    \I__3682\ : Span4Mux_h
    port map (
            O => \N__17533\,
            I => \N__17530\
        );

    \I__3681\ : Span4Mux_h
    port map (
            O => \N__17530\,
            I => \N__17527\
        );

    \I__3680\ : Span4Mux_v
    port map (
            O => \N__17527\,
            I => \N__17524\
        );

    \I__3679\ : Odrv4
    port map (
            O => \N__17524\,
            I => \line_buffer.n434\
        );

    \I__3678\ : InMux
    port map (
            O => \N__17521\,
            I => \N__17518\
        );

    \I__3677\ : LocalMux
    port map (
            O => \N__17518\,
            I => \line_buffer.n3749\
        );

    \I__3676\ : InMux
    port map (
            O => \N__17515\,
            I => \N__17512\
        );

    \I__3675\ : LocalMux
    port map (
            O => \N__17512\,
            I => \N__17509\
        );

    \I__3674\ : Span4Mux_v
    port map (
            O => \N__17509\,
            I => \N__17506\
        );

    \I__3673\ : Span4Mux_h
    port map (
            O => \N__17506\,
            I => \N__17503\
        );

    \I__3672\ : Span4Mux_h
    port map (
            O => \N__17503\,
            I => \N__17500\
        );

    \I__3671\ : Odrv4
    port map (
            O => \N__17500\,
            I => \line_buffer.n541\
        );

    \I__3670\ : InMux
    port map (
            O => \N__17497\,
            I => \N__17494\
        );

    \I__3669\ : LocalMux
    port map (
            O => \N__17494\,
            I => \N__17491\
        );

    \I__3668\ : Span4Mux_v
    port map (
            O => \N__17491\,
            I => \N__17488\
        );

    \I__3667\ : Span4Mux_h
    port map (
            O => \N__17488\,
            I => \N__17485\
        );

    \I__3666\ : Span4Mux_h
    port map (
            O => \N__17485\,
            I => \N__17482\
        );

    \I__3665\ : Odrv4
    port map (
            O => \N__17482\,
            I => \line_buffer.n533\
        );

    \I__3664\ : InMux
    port map (
            O => \N__17479\,
            I => \N__17476\
        );

    \I__3663\ : LocalMux
    port map (
            O => \N__17476\,
            I => \N__17473\
        );

    \I__3662\ : Span12Mux_v
    port map (
            O => \N__17473\,
            I => \N__17470\
        );

    \I__3661\ : Odrv12
    port map (
            O => \N__17470\,
            I => \line_buffer.n3676\
        );

    \I__3660\ : InMux
    port map (
            O => \N__17467\,
            I => \N__17464\
        );

    \I__3659\ : LocalMux
    port map (
            O => \N__17464\,
            I => \line_buffer.n3674\
        );

    \I__3658\ : InMux
    port map (
            O => \N__17461\,
            I => \N__17458\
        );

    \I__3657\ : LocalMux
    port map (
            O => \N__17458\,
            I => \line_buffer.n3716\
        );

    \I__3656\ : InMux
    port map (
            O => \N__17455\,
            I => \N__17452\
        );

    \I__3655\ : LocalMux
    port map (
            O => \N__17452\,
            I => \N__17449\
        );

    \I__3654\ : Span4Mux_v
    port map (
            O => \N__17449\,
            I => \N__17446\
        );

    \I__3653\ : Sp12to4
    port map (
            O => \N__17446\,
            I => \N__17443\
        );

    \I__3652\ : Odrv12
    port map (
            O => \N__17443\,
            I => \line_buffer.n446\
        );

    \I__3651\ : InMux
    port map (
            O => \N__17440\,
            I => \N__17437\
        );

    \I__3650\ : LocalMux
    port map (
            O => \N__17437\,
            I => \N__17434\
        );

    \I__3649\ : Span12Mux_h
    port map (
            O => \N__17434\,
            I => \N__17431\
        );

    \I__3648\ : Span12Mux_v
    port map (
            O => \N__17431\,
            I => \N__17428\
        );

    \I__3647\ : Odrv12
    port map (
            O => \N__17428\,
            I => \line_buffer.n438\
        );

    \I__3646\ : InMux
    port map (
            O => \N__17425\,
            I => \N__17422\
        );

    \I__3645\ : LocalMux
    port map (
            O => \N__17422\,
            I => \line_buffer.n3728\
        );

    \I__3644\ : CascadeMux
    port map (
            O => \N__17419\,
            I => \line_buffer.n3640_cascade_\
        );

    \I__3643\ : InMux
    port map (
            O => \N__17416\,
            I => \N__17413\
        );

    \I__3642\ : LocalMux
    port map (
            O => \N__17413\,
            I => \N__17410\
        );

    \I__3641\ : Span4Mux_v
    port map (
            O => \N__17410\,
            I => \N__17407\
        );

    \I__3640\ : Span4Mux_v
    port map (
            O => \N__17407\,
            I => \N__17404\
        );

    \I__3639\ : Odrv4
    port map (
            O => \N__17404\,
            I => \line_buffer.n3641\
        );

    \I__3638\ : InMux
    port map (
            O => \N__17401\,
            I => \N__17398\
        );

    \I__3637\ : LocalMux
    port map (
            O => \N__17398\,
            I => \N__17395\
        );

    \I__3636\ : Odrv12
    port map (
            O => \N__17395\,
            I => \RX_TX_SYNC_BUFF\
        );

    \I__3635\ : InMux
    port map (
            O => \N__17392\,
            I => \N__17389\
        );

    \I__3634\ : LocalMux
    port map (
            O => \N__17389\,
            I => \N__17386\
        );

    \I__3633\ : Span4Mux_v
    port map (
            O => \N__17386\,
            I => \N__17383\
        );

    \I__3632\ : Odrv4
    port map (
            O => \N__17383\,
            I => \RX_TX_SYNC\
        );

    \I__3631\ : InMux
    port map (
            O => \N__17380\,
            I => \N__17377\
        );

    \I__3630\ : LocalMux
    port map (
            O => \N__17377\,
            I => \sync_buffer.BUFFER_0\
        );

    \I__3629\ : InMux
    port map (
            O => \N__17374\,
            I => \N__17371\
        );

    \I__3628\ : LocalMux
    port map (
            O => \N__17371\,
            I => \sync_buffer.BUFFER_1\
        );

    \I__3627\ : InMux
    port map (
            O => \N__17368\,
            I => \N__17365\
        );

    \I__3626\ : LocalMux
    port map (
            O => \N__17365\,
            I => \transmit_module.n124\
        );

    \I__3625\ : CascadeMux
    port map (
            O => \N__17362\,
            I => \transmit_module.n139_cascade_\
        );

    \I__3624\ : InMux
    port map (
            O => \N__17359\,
            I => \N__17356\
        );

    \I__3623\ : LocalMux
    port map (
            O => \N__17356\,
            I => \transmit_module.ADDR_Y_COMPONENT_8\
        );

    \I__3622\ : CascadeMux
    port map (
            O => \N__17353\,
            I => \N__17347\
        );

    \I__3621\ : InMux
    port map (
            O => \N__17352\,
            I => \N__17342\
        );

    \I__3620\ : InMux
    port map (
            O => \N__17351\,
            I => \N__17342\
        );

    \I__3619\ : InMux
    port map (
            O => \N__17350\,
            I => \N__17337\
        );

    \I__3618\ : InMux
    port map (
            O => \N__17347\,
            I => \N__17337\
        );

    \I__3617\ : LocalMux
    port map (
            O => \N__17342\,
            I => \transmit_module.TX_ADDR_8\
        );

    \I__3616\ : LocalMux
    port map (
            O => \N__17337\,
            I => \transmit_module.TX_ADDR_8\
        );

    \I__3615\ : CascadeMux
    port map (
            O => \N__17332\,
            I => \N__17326\
        );

    \I__3614\ : InMux
    port map (
            O => \N__17331\,
            I => \N__17323\
        );

    \I__3613\ : InMux
    port map (
            O => \N__17330\,
            I => \N__17320\
        );

    \I__3612\ : InMux
    port map (
            O => \N__17329\,
            I => \N__17315\
        );

    \I__3611\ : InMux
    port map (
            O => \N__17326\,
            I => \N__17315\
        );

    \I__3610\ : LocalMux
    port map (
            O => \N__17323\,
            I => \transmit_module.TX_ADDR_9\
        );

    \I__3609\ : LocalMux
    port map (
            O => \N__17320\,
            I => \transmit_module.TX_ADDR_9\
        );

    \I__3608\ : LocalMux
    port map (
            O => \N__17315\,
            I => \transmit_module.TX_ADDR_9\
        );

    \I__3607\ : InMux
    port map (
            O => \N__17308\,
            I => \N__17305\
        );

    \I__3606\ : LocalMux
    port map (
            O => \N__17305\,
            I => \transmit_module.n123\
        );

    \I__3605\ : InMux
    port map (
            O => \N__17302\,
            I => \N__17299\
        );

    \I__3604\ : LocalMux
    port map (
            O => \N__17299\,
            I => \transmit_module.n138\
        );

    \I__3603\ : CascadeMux
    port map (
            O => \N__17296\,
            I => \transmit_module.n138_cascade_\
        );

    \I__3602\ : InMux
    port map (
            O => \N__17293\,
            I => \N__17287\
        );

    \I__3601\ : InMux
    port map (
            O => \N__17292\,
            I => \N__17287\
        );

    \I__3600\ : LocalMux
    port map (
            O => \N__17287\,
            I => \transmit_module.n107\
        );

    \I__3599\ : CascadeMux
    port map (
            O => \N__17284\,
            I => \N__17280\
        );

    \I__3598\ : CascadeMux
    port map (
            O => \N__17283\,
            I => \N__17277\
        );

    \I__3597\ : CascadeBuf
    port map (
            O => \N__17280\,
            I => \N__17274\
        );

    \I__3596\ : CascadeBuf
    port map (
            O => \N__17277\,
            I => \N__17271\
        );

    \I__3595\ : CascadeMux
    port map (
            O => \N__17274\,
            I => \N__17268\
        );

    \I__3594\ : CascadeMux
    port map (
            O => \N__17271\,
            I => \N__17265\
        );

    \I__3593\ : CascadeBuf
    port map (
            O => \N__17268\,
            I => \N__17262\
        );

    \I__3592\ : CascadeBuf
    port map (
            O => \N__17265\,
            I => \N__17259\
        );

    \I__3591\ : CascadeMux
    port map (
            O => \N__17262\,
            I => \N__17256\
        );

    \I__3590\ : CascadeMux
    port map (
            O => \N__17259\,
            I => \N__17253\
        );

    \I__3589\ : CascadeBuf
    port map (
            O => \N__17256\,
            I => \N__17250\
        );

    \I__3588\ : CascadeBuf
    port map (
            O => \N__17253\,
            I => \N__17247\
        );

    \I__3587\ : CascadeMux
    port map (
            O => \N__17250\,
            I => \N__17244\
        );

    \I__3586\ : CascadeMux
    port map (
            O => \N__17247\,
            I => \N__17241\
        );

    \I__3585\ : CascadeBuf
    port map (
            O => \N__17244\,
            I => \N__17238\
        );

    \I__3584\ : CascadeBuf
    port map (
            O => \N__17241\,
            I => \N__17235\
        );

    \I__3583\ : CascadeMux
    port map (
            O => \N__17238\,
            I => \N__17232\
        );

    \I__3582\ : CascadeMux
    port map (
            O => \N__17235\,
            I => \N__17229\
        );

    \I__3581\ : CascadeBuf
    port map (
            O => \N__17232\,
            I => \N__17226\
        );

    \I__3580\ : CascadeBuf
    port map (
            O => \N__17229\,
            I => \N__17223\
        );

    \I__3579\ : CascadeMux
    port map (
            O => \N__17226\,
            I => \N__17220\
        );

    \I__3578\ : CascadeMux
    port map (
            O => \N__17223\,
            I => \N__17217\
        );

    \I__3577\ : CascadeBuf
    port map (
            O => \N__17220\,
            I => \N__17214\
        );

    \I__3576\ : CascadeBuf
    port map (
            O => \N__17217\,
            I => \N__17211\
        );

    \I__3575\ : CascadeMux
    port map (
            O => \N__17214\,
            I => \N__17208\
        );

    \I__3574\ : CascadeMux
    port map (
            O => \N__17211\,
            I => \N__17205\
        );

    \I__3573\ : CascadeBuf
    port map (
            O => \N__17208\,
            I => \N__17202\
        );

    \I__3572\ : CascadeBuf
    port map (
            O => \N__17205\,
            I => \N__17199\
        );

    \I__3571\ : CascadeMux
    port map (
            O => \N__17202\,
            I => \N__17196\
        );

    \I__3570\ : CascadeMux
    port map (
            O => \N__17199\,
            I => \N__17193\
        );

    \I__3569\ : CascadeBuf
    port map (
            O => \N__17196\,
            I => \N__17190\
        );

    \I__3568\ : CascadeBuf
    port map (
            O => \N__17193\,
            I => \N__17187\
        );

    \I__3567\ : CascadeMux
    port map (
            O => \N__17190\,
            I => \N__17184\
        );

    \I__3566\ : CascadeMux
    port map (
            O => \N__17187\,
            I => \N__17181\
        );

    \I__3565\ : CascadeBuf
    port map (
            O => \N__17184\,
            I => \N__17178\
        );

    \I__3564\ : CascadeBuf
    port map (
            O => \N__17181\,
            I => \N__17175\
        );

    \I__3563\ : CascadeMux
    port map (
            O => \N__17178\,
            I => \N__17172\
        );

    \I__3562\ : CascadeMux
    port map (
            O => \N__17175\,
            I => \N__17169\
        );

    \I__3561\ : CascadeBuf
    port map (
            O => \N__17172\,
            I => \N__17166\
        );

    \I__3560\ : CascadeBuf
    port map (
            O => \N__17169\,
            I => \N__17163\
        );

    \I__3559\ : CascadeMux
    port map (
            O => \N__17166\,
            I => \N__17160\
        );

    \I__3558\ : CascadeMux
    port map (
            O => \N__17163\,
            I => \N__17157\
        );

    \I__3557\ : CascadeBuf
    port map (
            O => \N__17160\,
            I => \N__17154\
        );

    \I__3556\ : CascadeBuf
    port map (
            O => \N__17157\,
            I => \N__17151\
        );

    \I__3555\ : CascadeMux
    port map (
            O => \N__17154\,
            I => \N__17148\
        );

    \I__3554\ : CascadeMux
    port map (
            O => \N__17151\,
            I => \N__17145\
        );

    \I__3553\ : CascadeBuf
    port map (
            O => \N__17148\,
            I => \N__17142\
        );

    \I__3552\ : CascadeBuf
    port map (
            O => \N__17145\,
            I => \N__17139\
        );

    \I__3551\ : CascadeMux
    port map (
            O => \N__17142\,
            I => \N__17136\
        );

    \I__3550\ : CascadeMux
    port map (
            O => \N__17139\,
            I => \N__17133\
        );

    \I__3549\ : CascadeBuf
    port map (
            O => \N__17136\,
            I => \N__17130\
        );

    \I__3548\ : CascadeBuf
    port map (
            O => \N__17133\,
            I => \N__17127\
        );

    \I__3547\ : CascadeMux
    port map (
            O => \N__17130\,
            I => \N__17124\
        );

    \I__3546\ : CascadeMux
    port map (
            O => \N__17127\,
            I => \N__17121\
        );

    \I__3545\ : CascadeBuf
    port map (
            O => \N__17124\,
            I => \N__17118\
        );

    \I__3544\ : CascadeBuf
    port map (
            O => \N__17121\,
            I => \N__17115\
        );

    \I__3543\ : CascadeMux
    port map (
            O => \N__17118\,
            I => \N__17112\
        );

    \I__3542\ : CascadeMux
    port map (
            O => \N__17115\,
            I => \N__17109\
        );

    \I__3541\ : CascadeBuf
    port map (
            O => \N__17112\,
            I => \N__17106\
        );

    \I__3540\ : CascadeBuf
    port map (
            O => \N__17109\,
            I => \N__17103\
        );

    \I__3539\ : CascadeMux
    port map (
            O => \N__17106\,
            I => \N__17100\
        );

    \I__3538\ : CascadeMux
    port map (
            O => \N__17103\,
            I => \N__17097\
        );

    \I__3537\ : InMux
    port map (
            O => \N__17100\,
            I => \N__17094\
        );

    \I__3536\ : InMux
    port map (
            O => \N__17097\,
            I => \N__17091\
        );

    \I__3535\ : LocalMux
    port map (
            O => \N__17094\,
            I => \N__17088\
        );

    \I__3534\ : LocalMux
    port map (
            O => \N__17091\,
            I => \N__17085\
        );

    \I__3533\ : Span4Mux_v
    port map (
            O => \N__17088\,
            I => \N__17082\
        );

    \I__3532\ : Span4Mux_v
    port map (
            O => \N__17085\,
            I => \N__17079\
        );

    \I__3531\ : Span4Mux_v
    port map (
            O => \N__17082\,
            I => \N__17076\
        );

    \I__3530\ : Span4Mux_v
    port map (
            O => \N__17079\,
            I => \N__17073\
        );

    \I__3529\ : Span4Mux_v
    port map (
            O => \N__17076\,
            I => \N__17070\
        );

    \I__3528\ : Sp12to4
    port map (
            O => \N__17073\,
            I => \N__17067\
        );

    \I__3527\ : Span4Mux_v
    port map (
            O => \N__17070\,
            I => \N__17064\
        );

    \I__3526\ : Span12Mux_v
    port map (
            O => \N__17067\,
            I => \N__17061\
        );

    \I__3525\ : Span4Mux_h
    port map (
            O => \N__17064\,
            I => \N__17058\
        );

    \I__3524\ : Odrv12
    port map (
            O => \N__17061\,
            I => n19
        );

    \I__3523\ : Odrv4
    port map (
            O => \N__17058\,
            I => n19
        );

    \I__3522\ : CEMux
    port map (
            O => \N__17053\,
            I => \N__17050\
        );

    \I__3521\ : LocalMux
    port map (
            O => \N__17050\,
            I => \N__17047\
        );

    \I__3520\ : Span4Mux_v
    port map (
            O => \N__17047\,
            I => \N__17044\
        );

    \I__3519\ : Odrv4
    port map (
            O => \N__17044\,
            I => \receive_module.n3795\
        );

    \I__3518\ : SRMux
    port map (
            O => \N__17041\,
            I => \N__17037\
        );

    \I__3517\ : SRMux
    port map (
            O => \N__17040\,
            I => \N__17034\
        );

    \I__3516\ : LocalMux
    port map (
            O => \N__17037\,
            I => \N__17028\
        );

    \I__3515\ : LocalMux
    port map (
            O => \N__17034\,
            I => \N__17028\
        );

    \I__3514\ : SRMux
    port map (
            O => \N__17033\,
            I => \N__17025\
        );

    \I__3513\ : Span4Mux_v
    port map (
            O => \N__17028\,
            I => \N__17019\
        );

    \I__3512\ : LocalMux
    port map (
            O => \N__17025\,
            I => \N__17019\
        );

    \I__3511\ : SRMux
    port map (
            O => \N__17024\,
            I => \N__17016\
        );

    \I__3510\ : Span4Mux_h
    port map (
            O => \N__17019\,
            I => \N__17013\
        );

    \I__3509\ : LocalMux
    port map (
            O => \N__17016\,
            I => \N__17010\
        );

    \I__3508\ : Span4Mux_h
    port map (
            O => \N__17013\,
            I => \N__17007\
        );

    \I__3507\ : Span4Mux_v
    port map (
            O => \N__17010\,
            I => \N__17004\
        );

    \I__3506\ : Sp12to4
    port map (
            O => \N__17007\,
            I => \N__17001\
        );

    \I__3505\ : Span4Mux_h
    port map (
            O => \N__17004\,
            I => \N__16998\
        );

    \I__3504\ : Span12Mux_s10_v
    port map (
            O => \N__17001\,
            I => \N__16995\
        );

    \I__3503\ : Span4Mux_h
    port map (
            O => \N__16998\,
            I => \N__16992\
        );

    \I__3502\ : Odrv12
    port map (
            O => \N__16995\,
            I => \line_buffer.n451\
        );

    \I__3501\ : Odrv4
    port map (
            O => \N__16992\,
            I => \line_buffer.n451\
        );

    \I__3500\ : SRMux
    port map (
            O => \N__16987\,
            I => \N__16983\
        );

    \I__3499\ : SRMux
    port map (
            O => \N__16986\,
            I => \N__16980\
        );

    \I__3498\ : LocalMux
    port map (
            O => \N__16983\,
            I => \N__16977\
        );

    \I__3497\ : LocalMux
    port map (
            O => \N__16980\,
            I => \N__16973\
        );

    \I__3496\ : Span4Mux_v
    port map (
            O => \N__16977\,
            I => \N__16969\
        );

    \I__3495\ : SRMux
    port map (
            O => \N__16976\,
            I => \N__16966\
        );

    \I__3494\ : Span4Mux_h
    port map (
            O => \N__16973\,
            I => \N__16963\
        );

    \I__3493\ : SRMux
    port map (
            O => \N__16972\,
            I => \N__16960\
        );

    \I__3492\ : Sp12to4
    port map (
            O => \N__16969\,
            I => \N__16957\
        );

    \I__3491\ : LocalMux
    port map (
            O => \N__16966\,
            I => \N__16954\
        );

    \I__3490\ : Span4Mux_v
    port map (
            O => \N__16963\,
            I => \N__16949\
        );

    \I__3489\ : LocalMux
    port map (
            O => \N__16960\,
            I => \N__16949\
        );

    \I__3488\ : Span12Mux_v
    port map (
            O => \N__16957\,
            I => \N__16942\
        );

    \I__3487\ : Span12Mux_s11_v
    port map (
            O => \N__16954\,
            I => \N__16942\
        );

    \I__3486\ : Sp12to4
    port map (
            O => \N__16949\,
            I => \N__16942\
        );

    \I__3485\ : Odrv12
    port map (
            O => \N__16942\,
            I => \line_buffer.n549\
        );

    \I__3484\ : SRMux
    port map (
            O => \N__16939\,
            I => \N__16936\
        );

    \I__3483\ : LocalMux
    port map (
            O => \N__16936\,
            I => \N__16932\
        );

    \I__3482\ : SRMux
    port map (
            O => \N__16935\,
            I => \N__16929\
        );

    \I__3481\ : Span4Mux_s3_v
    port map (
            O => \N__16932\,
            I => \N__16925\
        );

    \I__3480\ : LocalMux
    port map (
            O => \N__16929\,
            I => \N__16922\
        );

    \I__3479\ : SRMux
    port map (
            O => \N__16928\,
            I => \N__16919\
        );

    \I__3478\ : Span4Mux_v
    port map (
            O => \N__16925\,
            I => \N__16912\
        );

    \I__3477\ : Span4Mux_h
    port map (
            O => \N__16922\,
            I => \N__16912\
        );

    \I__3476\ : LocalMux
    port map (
            O => \N__16919\,
            I => \N__16912\
        );

    \I__3475\ : Span4Mux_v
    port map (
            O => \N__16912\,
            I => \N__16909\
        );

    \I__3474\ : Span4Mux_h
    port map (
            O => \N__16909\,
            I => \N__16905\
        );

    \I__3473\ : SRMux
    port map (
            O => \N__16908\,
            I => \N__16902\
        );

    \I__3472\ : Sp12to4
    port map (
            O => \N__16905\,
            I => \N__16897\
        );

    \I__3471\ : LocalMux
    port map (
            O => \N__16902\,
            I => \N__16897\
        );

    \I__3470\ : Span12Mux_h
    port map (
            O => \N__16897\,
            I => \N__16894\
        );

    \I__3469\ : Odrv12
    port map (
            O => \N__16894\,
            I => \line_buffer.n516\
        );

    \I__3468\ : InMux
    port map (
            O => \N__16891\,
            I => \N__16888\
        );

    \I__3467\ : LocalMux
    port map (
            O => \N__16888\,
            I => \N__16885\
        );

    \I__3466\ : Span4Mux_h
    port map (
            O => \N__16885\,
            I => \N__16882\
        );

    \I__3465\ : Odrv4
    port map (
            O => \N__16882\,
            I => \receive_module.rx_counter.n3575\
        );

    \I__3464\ : InMux
    port map (
            O => \N__16879\,
            I => \N__16876\
        );

    \I__3463\ : LocalMux
    port map (
            O => \N__16876\,
            I => \N__16873\
        );

    \I__3462\ : Odrv4
    port map (
            O => \N__16873\,
            I => \receive_module.rx_counter.n4_adj_606\
        );

    \I__3461\ : CascadeMux
    port map (
            O => \N__16870\,
            I => \N__16867\
        );

    \I__3460\ : InMux
    port map (
            O => \N__16867\,
            I => \N__16864\
        );

    \I__3459\ : LocalMux
    port map (
            O => \N__16864\,
            I => \N__16859\
        );

    \I__3458\ : CascadeMux
    port map (
            O => \N__16863\,
            I => \N__16855\
        );

    \I__3457\ : InMux
    port map (
            O => \N__16862\,
            I => \N__16852\
        );

    \I__3456\ : Span4Mux_h
    port map (
            O => \N__16859\,
            I => \N__16849\
        );

    \I__3455\ : InMux
    port map (
            O => \N__16858\,
            I => \N__16846\
        );

    \I__3454\ : InMux
    port map (
            O => \N__16855\,
            I => \N__16843\
        );

    \I__3453\ : LocalMux
    port map (
            O => \N__16852\,
            I => \receive_module.rx_counter.Y_8\
        );

    \I__3452\ : Odrv4
    port map (
            O => \N__16849\,
            I => \receive_module.rx_counter.Y_8\
        );

    \I__3451\ : LocalMux
    port map (
            O => \N__16846\,
            I => \receive_module.rx_counter.Y_8\
        );

    \I__3450\ : LocalMux
    port map (
            O => \N__16843\,
            I => \receive_module.rx_counter.Y_8\
        );

    \I__3449\ : InMux
    port map (
            O => \N__16834\,
            I => \N__16831\
        );

    \I__3448\ : LocalMux
    port map (
            O => \N__16831\,
            I => \receive_module.rx_counter.n55_adj_607\
        );

    \I__3447\ : SRMux
    port map (
            O => \N__16828\,
            I => \N__16825\
        );

    \I__3446\ : LocalMux
    port map (
            O => \N__16825\,
            I => \N__16821\
        );

    \I__3445\ : SRMux
    port map (
            O => \N__16824\,
            I => \N__16818\
        );

    \I__3444\ : Span4Mux_v
    port map (
            O => \N__16821\,
            I => \N__16812\
        );

    \I__3443\ : LocalMux
    port map (
            O => \N__16818\,
            I => \N__16812\
        );

    \I__3442\ : SRMux
    port map (
            O => \N__16817\,
            I => \N__16809\
        );

    \I__3441\ : Span4Mux_v
    port map (
            O => \N__16812\,
            I => \N__16803\
        );

    \I__3440\ : LocalMux
    port map (
            O => \N__16809\,
            I => \N__16803\
        );

    \I__3439\ : SRMux
    port map (
            O => \N__16808\,
            I => \N__16800\
        );

    \I__3438\ : Span4Mux_v
    port map (
            O => \N__16803\,
            I => \N__16795\
        );

    \I__3437\ : LocalMux
    port map (
            O => \N__16800\,
            I => \N__16795\
        );

    \I__3436\ : Span4Mux_h
    port map (
            O => \N__16795\,
            I => \N__16792\
        );

    \I__3435\ : Span4Mux_h
    port map (
            O => \N__16792\,
            I => \N__16789\
        );

    \I__3434\ : Odrv4
    port map (
            O => \N__16789\,
            I => \line_buffer.n581\
        );

    \I__3433\ : CascadeMux
    port map (
            O => \N__16786\,
            I => \N__16776\
        );

    \I__3432\ : CascadeMux
    port map (
            O => \N__16785\,
            I => \N__16773\
        );

    \I__3431\ : InMux
    port map (
            O => \N__16784\,
            I => \N__16769\
        );

    \I__3430\ : InMux
    port map (
            O => \N__16783\,
            I => \N__16762\
        );

    \I__3429\ : InMux
    port map (
            O => \N__16782\,
            I => \N__16762\
        );

    \I__3428\ : InMux
    port map (
            O => \N__16781\,
            I => \N__16762\
        );

    \I__3427\ : InMux
    port map (
            O => \N__16780\,
            I => \N__16757\
        );

    \I__3426\ : InMux
    port map (
            O => \N__16779\,
            I => \N__16757\
        );

    \I__3425\ : InMux
    port map (
            O => \N__16776\,
            I => \N__16750\
        );

    \I__3424\ : InMux
    port map (
            O => \N__16773\,
            I => \N__16750\
        );

    \I__3423\ : InMux
    port map (
            O => \N__16772\,
            I => \N__16750\
        );

    \I__3422\ : LocalMux
    port map (
            O => \N__16769\,
            I => \RX_ADDR_12\
        );

    \I__3421\ : LocalMux
    port map (
            O => \N__16762\,
            I => \RX_ADDR_12\
        );

    \I__3420\ : LocalMux
    port map (
            O => \N__16757\,
            I => \RX_ADDR_12\
        );

    \I__3419\ : LocalMux
    port map (
            O => \N__16750\,
            I => \RX_ADDR_12\
        );

    \I__3418\ : CascadeMux
    port map (
            O => \N__16741\,
            I => \N__16732\
        );

    \I__3417\ : CascadeMux
    port map (
            O => \N__16740\,
            I => \N__16729\
        );

    \I__3416\ : CascadeMux
    port map (
            O => \N__16739\,
            I => \N__16726\
        );

    \I__3415\ : CascadeMux
    port map (
            O => \N__16738\,
            I => \N__16721\
        );

    \I__3414\ : InMux
    port map (
            O => \N__16737\,
            I => \N__16718\
        );

    \I__3413\ : InMux
    port map (
            O => \N__16736\,
            I => \N__16711\
        );

    \I__3412\ : InMux
    port map (
            O => \N__16735\,
            I => \N__16711\
        );

    \I__3411\ : InMux
    port map (
            O => \N__16732\,
            I => \N__16711\
        );

    \I__3410\ : InMux
    port map (
            O => \N__16729\,
            I => \N__16708\
        );

    \I__3409\ : InMux
    port map (
            O => \N__16726\,
            I => \N__16705\
        );

    \I__3408\ : InMux
    port map (
            O => \N__16725\,
            I => \N__16698\
        );

    \I__3407\ : InMux
    port map (
            O => \N__16724\,
            I => \N__16698\
        );

    \I__3406\ : InMux
    port map (
            O => \N__16721\,
            I => \N__16698\
        );

    \I__3405\ : LocalMux
    port map (
            O => \N__16718\,
            I => \RX_ADDR_13\
        );

    \I__3404\ : LocalMux
    port map (
            O => \N__16711\,
            I => \RX_ADDR_13\
        );

    \I__3403\ : LocalMux
    port map (
            O => \N__16708\,
            I => \RX_ADDR_13\
        );

    \I__3402\ : LocalMux
    port map (
            O => \N__16705\,
            I => \RX_ADDR_13\
        );

    \I__3401\ : LocalMux
    port map (
            O => \N__16698\,
            I => \RX_ADDR_13\
        );

    \I__3400\ : CascadeMux
    port map (
            O => \N__16687\,
            I => \N__16682\
        );

    \I__3399\ : CascadeMux
    port map (
            O => \N__16686\,
            I => \N__16679\
        );

    \I__3398\ : InMux
    port map (
            O => \N__16685\,
            I => \N__16670\
        );

    \I__3397\ : InMux
    port map (
            O => \N__16682\,
            I => \N__16665\
        );

    \I__3396\ : InMux
    port map (
            O => \N__16679\,
            I => \N__16665\
        );

    \I__3395\ : InMux
    port map (
            O => \N__16678\,
            I => \N__16662\
        );

    \I__3394\ : InMux
    port map (
            O => \N__16677\,
            I => \N__16657\
        );

    \I__3393\ : InMux
    port map (
            O => \N__16676\,
            I => \N__16657\
        );

    \I__3392\ : InMux
    port map (
            O => \N__16675\,
            I => \N__16650\
        );

    \I__3391\ : InMux
    port map (
            O => \N__16674\,
            I => \N__16650\
        );

    \I__3390\ : InMux
    port map (
            O => \N__16673\,
            I => \N__16650\
        );

    \I__3389\ : LocalMux
    port map (
            O => \N__16670\,
            I => \RX_ADDR_11\
        );

    \I__3388\ : LocalMux
    port map (
            O => \N__16665\,
            I => \RX_ADDR_11\
        );

    \I__3387\ : LocalMux
    port map (
            O => \N__16662\,
            I => \RX_ADDR_11\
        );

    \I__3386\ : LocalMux
    port map (
            O => \N__16657\,
            I => \RX_ADDR_11\
        );

    \I__3385\ : LocalMux
    port map (
            O => \N__16650\,
            I => \RX_ADDR_11\
        );

    \I__3384\ : SRMux
    port map (
            O => \N__16639\,
            I => \N__16635\
        );

    \I__3383\ : SRMux
    port map (
            O => \N__16638\,
            I => \N__16631\
        );

    \I__3382\ : LocalMux
    port map (
            O => \N__16635\,
            I => \N__16628\
        );

    \I__3381\ : SRMux
    port map (
            O => \N__16634\,
            I => \N__16625\
        );

    \I__3380\ : LocalMux
    port map (
            O => \N__16631\,
            I => \N__16621\
        );

    \I__3379\ : Span4Mux_h
    port map (
            O => \N__16628\,
            I => \N__16618\
        );

    \I__3378\ : LocalMux
    port map (
            O => \N__16625\,
            I => \N__16615\
        );

    \I__3377\ : SRMux
    port map (
            O => \N__16624\,
            I => \N__16612\
        );

    \I__3376\ : Span4Mux_h
    port map (
            O => \N__16621\,
            I => \N__16609\
        );

    \I__3375\ : Span4Mux_v
    port map (
            O => \N__16618\,
            I => \N__16604\
        );

    \I__3374\ : Span4Mux_h
    port map (
            O => \N__16615\,
            I => \N__16604\
        );

    \I__3373\ : LocalMux
    port map (
            O => \N__16612\,
            I => \N__16601\
        );

    \I__3372\ : Span4Mux_v
    port map (
            O => \N__16609\,
            I => \N__16598\
        );

    \I__3371\ : Sp12to4
    port map (
            O => \N__16604\,
            I => \N__16595\
        );

    \I__3370\ : Span4Mux_v
    port map (
            O => \N__16601\,
            I => \N__16592\
        );

    \I__3369\ : Sp12to4
    port map (
            O => \N__16598\,
            I => \N__16587\
        );

    \I__3368\ : Span12Mux_s7_v
    port map (
            O => \N__16595\,
            I => \N__16587\
        );

    \I__3367\ : Span4Mux_h
    port map (
            O => \N__16592\,
            I => \N__16584\
        );

    \I__3366\ : Span12Mux_v
    port map (
            O => \N__16587\,
            I => \N__16581\
        );

    \I__3365\ : Span4Mux_h
    port map (
            O => \N__16584\,
            I => \N__16578\
        );

    \I__3364\ : Odrv12
    port map (
            O => \N__16581\,
            I => \line_buffer.n580\
        );

    \I__3363\ : Odrv4
    port map (
            O => \N__16578\,
            I => \line_buffer.n580\
        );

    \I__3362\ : InMux
    port map (
            O => \N__16573\,
            I => \N__16570\
        );

    \I__3361\ : LocalMux
    port map (
            O => \N__16570\,
            I => \N__16567\
        );

    \I__3360\ : Span4Mux_v
    port map (
            O => \N__16567\,
            I => \N__16564\
        );

    \I__3359\ : Span4Mux_h
    port map (
            O => \N__16564\,
            I => \N__16561\
        );

    \I__3358\ : Span4Mux_h
    port map (
            O => \N__16561\,
            I => \N__16558\
        );

    \I__3357\ : Odrv4
    port map (
            O => \N__16558\,
            I => \line_buffer.n511\
        );

    \I__3356\ : InMux
    port map (
            O => \N__16555\,
            I => \N__16552\
        );

    \I__3355\ : LocalMux
    port map (
            O => \N__16552\,
            I => \N__16549\
        );

    \I__3354\ : Span12Mux_h
    port map (
            O => \N__16549\,
            I => \N__16546\
        );

    \I__3353\ : Odrv12
    port map (
            O => \N__16546\,
            I => \line_buffer.n503\
        );

    \I__3352\ : InMux
    port map (
            O => \N__16543\,
            I => \N__16540\
        );

    \I__3351\ : LocalMux
    port map (
            O => \N__16540\,
            I => \N__16537\
        );

    \I__3350\ : Span4Mux_v
    port map (
            O => \N__16537\,
            I => \N__16534\
        );

    \I__3349\ : Span4Mux_h
    port map (
            O => \N__16534\,
            I => \N__16531\
        );

    \I__3348\ : Span4Mux_h
    port map (
            O => \N__16531\,
            I => \N__16528\
        );

    \I__3347\ : Odrv4
    port map (
            O => \N__16528\,
            I => \line_buffer.n509\
        );

    \I__3346\ : InMux
    port map (
            O => \N__16525\,
            I => \N__16522\
        );

    \I__3345\ : LocalMux
    port map (
            O => \N__16522\,
            I => \N__16519\
        );

    \I__3344\ : Span4Mux_v
    port map (
            O => \N__16519\,
            I => \N__16516\
        );

    \I__3343\ : Sp12to4
    port map (
            O => \N__16516\,
            I => \N__16513\
        );

    \I__3342\ : Odrv12
    port map (
            O => \N__16513\,
            I => \line_buffer.n501\
        );

    \I__3341\ : CascadeMux
    port map (
            O => \N__16510\,
            I => \receive_module.rx_counter.n4_cascade_\
        );

    \I__3340\ : CascadeMux
    port map (
            O => \N__16507\,
            I => \receive_module.rx_counter.n6_cascade_\
        );

    \I__3339\ : InMux
    port map (
            O => \N__16504\,
            I => \N__16501\
        );

    \I__3338\ : LocalMux
    port map (
            O => \N__16501\,
            I => \receive_module.rx_counter.n3534\
        );

    \I__3337\ : InMux
    port map (
            O => \N__16498\,
            I => \N__16495\
        );

    \I__3336\ : LocalMux
    port map (
            O => \N__16495\,
            I => \receive_module.rx_counter.n3581\
        );

    \I__3335\ : SRMux
    port map (
            O => \N__16492\,
            I => \N__16487\
        );

    \I__3334\ : SRMux
    port map (
            O => \N__16491\,
            I => \N__16484\
        );

    \I__3333\ : SRMux
    port map (
            O => \N__16490\,
            I => \N__16480\
        );

    \I__3332\ : LocalMux
    port map (
            O => \N__16487\,
            I => \N__16475\
        );

    \I__3331\ : LocalMux
    port map (
            O => \N__16484\,
            I => \N__16475\
        );

    \I__3330\ : SRMux
    port map (
            O => \N__16483\,
            I => \N__16472\
        );

    \I__3329\ : LocalMux
    port map (
            O => \N__16480\,
            I => \N__16469\
        );

    \I__3328\ : Span4Mux_s3_v
    port map (
            O => \N__16475\,
            I => \N__16464\
        );

    \I__3327\ : LocalMux
    port map (
            O => \N__16472\,
            I => \N__16464\
        );

    \I__3326\ : Sp12to4
    port map (
            O => \N__16469\,
            I => \N__16461\
        );

    \I__3325\ : Sp12to4
    port map (
            O => \N__16464\,
            I => \N__16458\
        );

    \I__3324\ : Span12Mux_h
    port map (
            O => \N__16461\,
            I => \N__16455\
        );

    \I__3323\ : Span12Mux_s10_v
    port map (
            O => \N__16458\,
            I => \N__16452\
        );

    \I__3322\ : Odrv12
    port map (
            O => \N__16455\,
            I => \line_buffer.n517\
        );

    \I__3321\ : Odrv12
    port map (
            O => \N__16452\,
            I => \line_buffer.n517\
        );

    \I__3320\ : SRMux
    port map (
            O => \N__16447\,
            I => \N__16443\
        );

    \I__3319\ : SRMux
    port map (
            O => \N__16446\,
            I => \N__16440\
        );

    \I__3318\ : LocalMux
    port map (
            O => \N__16443\,
            I => \N__16433\
        );

    \I__3317\ : LocalMux
    port map (
            O => \N__16440\,
            I => \N__16433\
        );

    \I__3316\ : SRMux
    port map (
            O => \N__16439\,
            I => \N__16430\
        );

    \I__3315\ : SRMux
    port map (
            O => \N__16438\,
            I => \N__16427\
        );

    \I__3314\ : Span4Mux_v
    port map (
            O => \N__16433\,
            I => \N__16420\
        );

    \I__3313\ : LocalMux
    port map (
            O => \N__16430\,
            I => \N__16420\
        );

    \I__3312\ : LocalMux
    port map (
            O => \N__16427\,
            I => \N__16420\
        );

    \I__3311\ : Span4Mux_v
    port map (
            O => \N__16420\,
            I => \N__16417\
        );

    \I__3310\ : Span4Mux_h
    port map (
            O => \N__16417\,
            I => \N__16414\
        );

    \I__3309\ : Span4Mux_h
    port map (
            O => \N__16414\,
            I => \N__16411\
        );

    \I__3308\ : Span4Mux_v
    port map (
            O => \N__16411\,
            I => \N__16408\
        );

    \I__3307\ : Odrv4
    port map (
            O => \N__16408\,
            I => \line_buffer.n452\
        );

    \I__3306\ : SRMux
    port map (
            O => \N__16405\,
            I => \N__16401\
        );

    \I__3305\ : SRMux
    port map (
            O => \N__16404\,
            I => \N__16398\
        );

    \I__3304\ : LocalMux
    port map (
            O => \N__16401\,
            I => \N__16391\
        );

    \I__3303\ : LocalMux
    port map (
            O => \N__16398\,
            I => \N__16391\
        );

    \I__3302\ : SRMux
    port map (
            O => \N__16397\,
            I => \N__16388\
        );

    \I__3301\ : SRMux
    port map (
            O => \N__16396\,
            I => \N__16385\
        );

    \I__3300\ : Span4Mux_v
    port map (
            O => \N__16391\,
            I => \N__16380\
        );

    \I__3299\ : LocalMux
    port map (
            O => \N__16388\,
            I => \N__16380\
        );

    \I__3298\ : LocalMux
    port map (
            O => \N__16385\,
            I => \N__16377\
        );

    \I__3297\ : Span4Mux_h
    port map (
            O => \N__16380\,
            I => \N__16374\
        );

    \I__3296\ : Sp12to4
    port map (
            O => \N__16377\,
            I => \N__16371\
        );

    \I__3295\ : Span4Mux_h
    port map (
            O => \N__16374\,
            I => \N__16368\
        );

    \I__3294\ : Span12Mux_h
    port map (
            O => \N__16371\,
            I => \N__16365\
        );

    \I__3293\ : Span4Mux_h
    port map (
            O => \N__16368\,
            I => \N__16362\
        );

    \I__3292\ : Odrv12
    port map (
            O => \N__16365\,
            I => \line_buffer.n548\
        );

    \I__3291\ : Odrv4
    port map (
            O => \N__16362\,
            I => \line_buffer.n548\
        );

    \I__3290\ : InMux
    port map (
            O => \N__16357\,
            I => \N__16353\
        );

    \I__3289\ : InMux
    port map (
            O => \N__16356\,
            I => \N__16350\
        );

    \I__3288\ : LocalMux
    port map (
            O => \N__16353\,
            I => \receive_module.rx_counter.FRAME_COUNTER_0\
        );

    \I__3287\ : LocalMux
    port map (
            O => \N__16350\,
            I => \receive_module.rx_counter.FRAME_COUNTER_0\
        );

    \I__3286\ : InMux
    port map (
            O => \N__16345\,
            I => \bfn_16_5_0_\
        );

    \I__3285\ : InMux
    port map (
            O => \N__16342\,
            I => \N__16338\
        );

    \I__3284\ : InMux
    port map (
            O => \N__16341\,
            I => \N__16335\
        );

    \I__3283\ : LocalMux
    port map (
            O => \N__16338\,
            I => \receive_module.rx_counter.FRAME_COUNTER_1\
        );

    \I__3282\ : LocalMux
    port map (
            O => \N__16335\,
            I => \receive_module.rx_counter.FRAME_COUNTER_1\
        );

    \I__3281\ : InMux
    port map (
            O => \N__16330\,
            I => \receive_module.rx_counter.n3310\
        );

    \I__3280\ : InMux
    port map (
            O => \N__16327\,
            I => \N__16323\
        );

    \I__3279\ : InMux
    port map (
            O => \N__16326\,
            I => \N__16320\
        );

    \I__3278\ : LocalMux
    port map (
            O => \N__16323\,
            I => \receive_module.rx_counter.FRAME_COUNTER_2\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__16320\,
            I => \receive_module.rx_counter.FRAME_COUNTER_2\
        );

    \I__3276\ : InMux
    port map (
            O => \N__16315\,
            I => \receive_module.rx_counter.n3311\
        );

    \I__3275\ : InMux
    port map (
            O => \N__16312\,
            I => \N__16308\
        );

    \I__3274\ : InMux
    port map (
            O => \N__16311\,
            I => \N__16305\
        );

    \I__3273\ : LocalMux
    port map (
            O => \N__16308\,
            I => \receive_module.rx_counter.FRAME_COUNTER_3\
        );

    \I__3272\ : LocalMux
    port map (
            O => \N__16305\,
            I => \receive_module.rx_counter.FRAME_COUNTER_3\
        );

    \I__3271\ : InMux
    port map (
            O => \N__16300\,
            I => \receive_module.rx_counter.n3312\
        );

    \I__3270\ : InMux
    port map (
            O => \N__16297\,
            I => \N__16293\
        );

    \I__3269\ : InMux
    port map (
            O => \N__16296\,
            I => \N__16290\
        );

    \I__3268\ : LocalMux
    port map (
            O => \N__16293\,
            I => \receive_module.rx_counter.FRAME_COUNTER_4\
        );

    \I__3267\ : LocalMux
    port map (
            O => \N__16290\,
            I => \receive_module.rx_counter.FRAME_COUNTER_4\
        );

    \I__3266\ : InMux
    port map (
            O => \N__16285\,
            I => \receive_module.rx_counter.n3313\
        );

    \I__3265\ : InMux
    port map (
            O => \N__16282\,
            I => \receive_module.rx_counter.n3314\
        );

    \I__3264\ : InMux
    port map (
            O => \N__16279\,
            I => \N__16275\
        );

    \I__3263\ : InMux
    port map (
            O => \N__16278\,
            I => \N__16272\
        );

    \I__3262\ : LocalMux
    port map (
            O => \N__16275\,
            I => \receive_module.rx_counter.FRAME_COUNTER_5\
        );

    \I__3261\ : LocalMux
    port map (
            O => \N__16272\,
            I => \receive_module.rx_counter.FRAME_COUNTER_5\
        );

    \I__3260\ : CEMux
    port map (
            O => \N__16267\,
            I => \N__16263\
        );

    \I__3259\ : CEMux
    port map (
            O => \N__16266\,
            I => \N__16260\
        );

    \I__3258\ : LocalMux
    port map (
            O => \N__16263\,
            I => \N__16257\
        );

    \I__3257\ : LocalMux
    port map (
            O => \N__16260\,
            I => \N__16254\
        );

    \I__3256\ : Span4Mux_v
    port map (
            O => \N__16257\,
            I => \N__16251\
        );

    \I__3255\ : Span4Mux_h
    port map (
            O => \N__16254\,
            I => \N__16248\
        );

    \I__3254\ : Odrv4
    port map (
            O => \N__16251\,
            I => \receive_module.rx_counter.n3792\
        );

    \I__3253\ : Odrv4
    port map (
            O => \N__16248\,
            I => \receive_module.rx_counter.n3792\
        );

    \I__3252\ : SRMux
    port map (
            O => \N__16243\,
            I => \N__16240\
        );

    \I__3251\ : LocalMux
    port map (
            O => \N__16240\,
            I => \N__16237\
        );

    \I__3250\ : Span4Mux_h
    port map (
            O => \N__16237\,
            I => \N__16234\
        );

    \I__3249\ : Odrv4
    port map (
            O => \N__16234\,
            I => \receive_module.rx_counter.n2517\
        );

    \I__3248\ : InMux
    port map (
            O => \N__16231\,
            I => \N__16228\
        );

    \I__3247\ : LocalMux
    port map (
            O => \N__16228\,
            I => \N__16225\
        );

    \I__3246\ : Span4Mux_h
    port map (
            O => \N__16225\,
            I => \N__16222\
        );

    \I__3245\ : Odrv4
    port map (
            O => \N__16222\,
            I => \receive_module.n136\
        );

    \I__3244\ : CascadeMux
    port map (
            O => \N__16219\,
            I => \N__16216\
        );

    \I__3243\ : CascadeBuf
    port map (
            O => \N__16216\,
            I => \N__16212\
        );

    \I__3242\ : CascadeMux
    port map (
            O => \N__16215\,
            I => \N__16209\
        );

    \I__3241\ : CascadeMux
    port map (
            O => \N__16212\,
            I => \N__16206\
        );

    \I__3240\ : CascadeBuf
    port map (
            O => \N__16209\,
            I => \N__16203\
        );

    \I__3239\ : CascadeBuf
    port map (
            O => \N__16206\,
            I => \N__16200\
        );

    \I__3238\ : CascadeMux
    port map (
            O => \N__16203\,
            I => \N__16197\
        );

    \I__3237\ : CascadeMux
    port map (
            O => \N__16200\,
            I => \N__16194\
        );

    \I__3236\ : CascadeBuf
    port map (
            O => \N__16197\,
            I => \N__16191\
        );

    \I__3235\ : CascadeBuf
    port map (
            O => \N__16194\,
            I => \N__16188\
        );

    \I__3234\ : CascadeMux
    port map (
            O => \N__16191\,
            I => \N__16185\
        );

    \I__3233\ : CascadeMux
    port map (
            O => \N__16188\,
            I => \N__16182\
        );

    \I__3232\ : CascadeBuf
    port map (
            O => \N__16185\,
            I => \N__16179\
        );

    \I__3231\ : CascadeBuf
    port map (
            O => \N__16182\,
            I => \N__16176\
        );

    \I__3230\ : CascadeMux
    port map (
            O => \N__16179\,
            I => \N__16173\
        );

    \I__3229\ : CascadeMux
    port map (
            O => \N__16176\,
            I => \N__16170\
        );

    \I__3228\ : CascadeBuf
    port map (
            O => \N__16173\,
            I => \N__16167\
        );

    \I__3227\ : CascadeBuf
    port map (
            O => \N__16170\,
            I => \N__16164\
        );

    \I__3226\ : CascadeMux
    port map (
            O => \N__16167\,
            I => \N__16161\
        );

    \I__3225\ : CascadeMux
    port map (
            O => \N__16164\,
            I => \N__16158\
        );

    \I__3224\ : CascadeBuf
    port map (
            O => \N__16161\,
            I => \N__16155\
        );

    \I__3223\ : CascadeBuf
    port map (
            O => \N__16158\,
            I => \N__16152\
        );

    \I__3222\ : CascadeMux
    port map (
            O => \N__16155\,
            I => \N__16149\
        );

    \I__3221\ : CascadeMux
    port map (
            O => \N__16152\,
            I => \N__16146\
        );

    \I__3220\ : CascadeBuf
    port map (
            O => \N__16149\,
            I => \N__16143\
        );

    \I__3219\ : CascadeBuf
    port map (
            O => \N__16146\,
            I => \N__16140\
        );

    \I__3218\ : CascadeMux
    port map (
            O => \N__16143\,
            I => \N__16137\
        );

    \I__3217\ : CascadeMux
    port map (
            O => \N__16140\,
            I => \N__16134\
        );

    \I__3216\ : CascadeBuf
    port map (
            O => \N__16137\,
            I => \N__16131\
        );

    \I__3215\ : CascadeBuf
    port map (
            O => \N__16134\,
            I => \N__16128\
        );

    \I__3214\ : CascadeMux
    port map (
            O => \N__16131\,
            I => \N__16125\
        );

    \I__3213\ : CascadeMux
    port map (
            O => \N__16128\,
            I => \N__16122\
        );

    \I__3212\ : CascadeBuf
    port map (
            O => \N__16125\,
            I => \N__16119\
        );

    \I__3211\ : CascadeBuf
    port map (
            O => \N__16122\,
            I => \N__16116\
        );

    \I__3210\ : CascadeMux
    port map (
            O => \N__16119\,
            I => \N__16113\
        );

    \I__3209\ : CascadeMux
    port map (
            O => \N__16116\,
            I => \N__16110\
        );

    \I__3208\ : CascadeBuf
    port map (
            O => \N__16113\,
            I => \N__16107\
        );

    \I__3207\ : CascadeBuf
    port map (
            O => \N__16110\,
            I => \N__16104\
        );

    \I__3206\ : CascadeMux
    port map (
            O => \N__16107\,
            I => \N__16101\
        );

    \I__3205\ : CascadeMux
    port map (
            O => \N__16104\,
            I => \N__16098\
        );

    \I__3204\ : CascadeBuf
    port map (
            O => \N__16101\,
            I => \N__16095\
        );

    \I__3203\ : CascadeBuf
    port map (
            O => \N__16098\,
            I => \N__16092\
        );

    \I__3202\ : CascadeMux
    port map (
            O => \N__16095\,
            I => \N__16089\
        );

    \I__3201\ : CascadeMux
    port map (
            O => \N__16092\,
            I => \N__16086\
        );

    \I__3200\ : CascadeBuf
    port map (
            O => \N__16089\,
            I => \N__16083\
        );

    \I__3199\ : CascadeBuf
    port map (
            O => \N__16086\,
            I => \N__16080\
        );

    \I__3198\ : CascadeMux
    port map (
            O => \N__16083\,
            I => \N__16077\
        );

    \I__3197\ : CascadeMux
    port map (
            O => \N__16080\,
            I => \N__16074\
        );

    \I__3196\ : CascadeBuf
    port map (
            O => \N__16077\,
            I => \N__16071\
        );

    \I__3195\ : CascadeBuf
    port map (
            O => \N__16074\,
            I => \N__16068\
        );

    \I__3194\ : CascadeMux
    port map (
            O => \N__16071\,
            I => \N__16065\
        );

    \I__3193\ : CascadeMux
    port map (
            O => \N__16068\,
            I => \N__16062\
        );

    \I__3192\ : CascadeBuf
    port map (
            O => \N__16065\,
            I => \N__16059\
        );

    \I__3191\ : CascadeBuf
    port map (
            O => \N__16062\,
            I => \N__16056\
        );

    \I__3190\ : CascadeMux
    port map (
            O => \N__16059\,
            I => \N__16053\
        );

    \I__3189\ : CascadeMux
    port map (
            O => \N__16056\,
            I => \N__16050\
        );

    \I__3188\ : CascadeBuf
    port map (
            O => \N__16053\,
            I => \N__16047\
        );

    \I__3187\ : CascadeBuf
    port map (
            O => \N__16050\,
            I => \N__16044\
        );

    \I__3186\ : CascadeMux
    port map (
            O => \N__16047\,
            I => \N__16041\
        );

    \I__3185\ : CascadeMux
    port map (
            O => \N__16044\,
            I => \N__16038\
        );

    \I__3184\ : CascadeBuf
    port map (
            O => \N__16041\,
            I => \N__16035\
        );

    \I__3183\ : InMux
    port map (
            O => \N__16038\,
            I => \N__16032\
        );

    \I__3182\ : CascadeMux
    port map (
            O => \N__16035\,
            I => \N__16029\
        );

    \I__3181\ : LocalMux
    port map (
            O => \N__16032\,
            I => \N__16026\
        );

    \I__3180\ : InMux
    port map (
            O => \N__16029\,
            I => \N__16023\
        );

    \I__3179\ : Span4Mux_s1_v
    port map (
            O => \N__16026\,
            I => \N__16020\
        );

    \I__3178\ : LocalMux
    port map (
            O => \N__16023\,
            I => \N__16017\
        );

    \I__3177\ : Span4Mux_h
    port map (
            O => \N__16020\,
            I => \N__16014\
        );

    \I__3176\ : Span4Mux_s1_v
    port map (
            O => \N__16017\,
            I => \N__16011\
        );

    \I__3175\ : Span4Mux_h
    port map (
            O => \N__16014\,
            I => \N__16007\
        );

    \I__3174\ : Span4Mux_v
    port map (
            O => \N__16011\,
            I => \N__16004\
        );

    \I__3173\ : InMux
    port map (
            O => \N__16010\,
            I => \N__16001\
        );

    \I__3172\ : Span4Mux_v
    port map (
            O => \N__16007\,
            I => \N__15998\
        );

    \I__3171\ : Sp12to4
    port map (
            O => \N__16004\,
            I => \N__15995\
        );

    \I__3170\ : LocalMux
    port map (
            O => \N__16001\,
            I => \N__15991\
        );

    \I__3169\ : Sp12to4
    port map (
            O => \N__15998\,
            I => \N__15986\
        );

    \I__3168\ : Span12Mux_h
    port map (
            O => \N__15995\,
            I => \N__15986\
        );

    \I__3167\ : InMux
    port map (
            O => \N__15994\,
            I => \N__15983\
        );

    \I__3166\ : Sp12to4
    port map (
            O => \N__15991\,
            I => \N__15978\
        );

    \I__3165\ : Span12Mux_v
    port map (
            O => \N__15986\,
            I => \N__15978\
        );

    \I__3164\ : LocalMux
    port map (
            O => \N__15983\,
            I => \RX_ADDR_0\
        );

    \I__3163\ : Odrv12
    port map (
            O => \N__15978\,
            I => \RX_ADDR_0\
        );

    \I__3162\ : CascadeMux
    port map (
            O => \N__15973\,
            I => \N__15970\
        );

    \I__3161\ : InMux
    port map (
            O => \N__15970\,
            I => \N__15967\
        );

    \I__3160\ : LocalMux
    port map (
            O => \N__15967\,
            I => \N__15964\
        );

    \I__3159\ : Span4Mux_h
    port map (
            O => \N__15964\,
            I => \N__15961\
        );

    \I__3158\ : Odrv4
    port map (
            O => \N__15961\,
            I => \receive_module.n135\
        );

    \I__3157\ : CascadeMux
    port map (
            O => \N__15958\,
            I => \N__15954\
        );

    \I__3156\ : CascadeMux
    port map (
            O => \N__15957\,
            I => \N__15951\
        );

    \I__3155\ : CascadeBuf
    port map (
            O => \N__15954\,
            I => \N__15948\
        );

    \I__3154\ : CascadeBuf
    port map (
            O => \N__15951\,
            I => \N__15945\
        );

    \I__3153\ : CascadeMux
    port map (
            O => \N__15948\,
            I => \N__15942\
        );

    \I__3152\ : CascadeMux
    port map (
            O => \N__15945\,
            I => \N__15939\
        );

    \I__3151\ : CascadeBuf
    port map (
            O => \N__15942\,
            I => \N__15936\
        );

    \I__3150\ : CascadeBuf
    port map (
            O => \N__15939\,
            I => \N__15933\
        );

    \I__3149\ : CascadeMux
    port map (
            O => \N__15936\,
            I => \N__15930\
        );

    \I__3148\ : CascadeMux
    port map (
            O => \N__15933\,
            I => \N__15927\
        );

    \I__3147\ : CascadeBuf
    port map (
            O => \N__15930\,
            I => \N__15924\
        );

    \I__3146\ : CascadeBuf
    port map (
            O => \N__15927\,
            I => \N__15921\
        );

    \I__3145\ : CascadeMux
    port map (
            O => \N__15924\,
            I => \N__15918\
        );

    \I__3144\ : CascadeMux
    port map (
            O => \N__15921\,
            I => \N__15915\
        );

    \I__3143\ : CascadeBuf
    port map (
            O => \N__15918\,
            I => \N__15912\
        );

    \I__3142\ : CascadeBuf
    port map (
            O => \N__15915\,
            I => \N__15909\
        );

    \I__3141\ : CascadeMux
    port map (
            O => \N__15912\,
            I => \N__15906\
        );

    \I__3140\ : CascadeMux
    port map (
            O => \N__15909\,
            I => \N__15903\
        );

    \I__3139\ : CascadeBuf
    port map (
            O => \N__15906\,
            I => \N__15900\
        );

    \I__3138\ : CascadeBuf
    port map (
            O => \N__15903\,
            I => \N__15897\
        );

    \I__3137\ : CascadeMux
    port map (
            O => \N__15900\,
            I => \N__15894\
        );

    \I__3136\ : CascadeMux
    port map (
            O => \N__15897\,
            I => \N__15891\
        );

    \I__3135\ : CascadeBuf
    port map (
            O => \N__15894\,
            I => \N__15888\
        );

    \I__3134\ : CascadeBuf
    port map (
            O => \N__15891\,
            I => \N__15885\
        );

    \I__3133\ : CascadeMux
    port map (
            O => \N__15888\,
            I => \N__15882\
        );

    \I__3132\ : CascadeMux
    port map (
            O => \N__15885\,
            I => \N__15879\
        );

    \I__3131\ : CascadeBuf
    port map (
            O => \N__15882\,
            I => \N__15876\
        );

    \I__3130\ : CascadeBuf
    port map (
            O => \N__15879\,
            I => \N__15873\
        );

    \I__3129\ : CascadeMux
    port map (
            O => \N__15876\,
            I => \N__15870\
        );

    \I__3128\ : CascadeMux
    port map (
            O => \N__15873\,
            I => \N__15867\
        );

    \I__3127\ : CascadeBuf
    port map (
            O => \N__15870\,
            I => \N__15864\
        );

    \I__3126\ : CascadeBuf
    port map (
            O => \N__15867\,
            I => \N__15861\
        );

    \I__3125\ : CascadeMux
    port map (
            O => \N__15864\,
            I => \N__15858\
        );

    \I__3124\ : CascadeMux
    port map (
            O => \N__15861\,
            I => \N__15855\
        );

    \I__3123\ : CascadeBuf
    port map (
            O => \N__15858\,
            I => \N__15852\
        );

    \I__3122\ : CascadeBuf
    port map (
            O => \N__15855\,
            I => \N__15849\
        );

    \I__3121\ : CascadeMux
    port map (
            O => \N__15852\,
            I => \N__15846\
        );

    \I__3120\ : CascadeMux
    port map (
            O => \N__15849\,
            I => \N__15843\
        );

    \I__3119\ : CascadeBuf
    port map (
            O => \N__15846\,
            I => \N__15840\
        );

    \I__3118\ : CascadeBuf
    port map (
            O => \N__15843\,
            I => \N__15837\
        );

    \I__3117\ : CascadeMux
    port map (
            O => \N__15840\,
            I => \N__15834\
        );

    \I__3116\ : CascadeMux
    port map (
            O => \N__15837\,
            I => \N__15831\
        );

    \I__3115\ : CascadeBuf
    port map (
            O => \N__15834\,
            I => \N__15828\
        );

    \I__3114\ : CascadeBuf
    port map (
            O => \N__15831\,
            I => \N__15825\
        );

    \I__3113\ : CascadeMux
    port map (
            O => \N__15828\,
            I => \N__15822\
        );

    \I__3112\ : CascadeMux
    port map (
            O => \N__15825\,
            I => \N__15819\
        );

    \I__3111\ : CascadeBuf
    port map (
            O => \N__15822\,
            I => \N__15816\
        );

    \I__3110\ : CascadeBuf
    port map (
            O => \N__15819\,
            I => \N__15813\
        );

    \I__3109\ : CascadeMux
    port map (
            O => \N__15816\,
            I => \N__15810\
        );

    \I__3108\ : CascadeMux
    port map (
            O => \N__15813\,
            I => \N__15807\
        );

    \I__3107\ : CascadeBuf
    port map (
            O => \N__15810\,
            I => \N__15804\
        );

    \I__3106\ : CascadeBuf
    port map (
            O => \N__15807\,
            I => \N__15801\
        );

    \I__3105\ : CascadeMux
    port map (
            O => \N__15804\,
            I => \N__15798\
        );

    \I__3104\ : CascadeMux
    port map (
            O => \N__15801\,
            I => \N__15795\
        );

    \I__3103\ : CascadeBuf
    port map (
            O => \N__15798\,
            I => \N__15792\
        );

    \I__3102\ : CascadeBuf
    port map (
            O => \N__15795\,
            I => \N__15789\
        );

    \I__3101\ : CascadeMux
    port map (
            O => \N__15792\,
            I => \N__15786\
        );

    \I__3100\ : CascadeMux
    port map (
            O => \N__15789\,
            I => \N__15783\
        );

    \I__3099\ : CascadeBuf
    port map (
            O => \N__15786\,
            I => \N__15780\
        );

    \I__3098\ : CascadeBuf
    port map (
            O => \N__15783\,
            I => \N__15777\
        );

    \I__3097\ : CascadeMux
    port map (
            O => \N__15780\,
            I => \N__15774\
        );

    \I__3096\ : CascadeMux
    port map (
            O => \N__15777\,
            I => \N__15771\
        );

    \I__3095\ : InMux
    port map (
            O => \N__15774\,
            I => \N__15768\
        );

    \I__3094\ : InMux
    port map (
            O => \N__15771\,
            I => \N__15765\
        );

    \I__3093\ : LocalMux
    port map (
            O => \N__15768\,
            I => \N__15762\
        );

    \I__3092\ : LocalMux
    port map (
            O => \N__15765\,
            I => \N__15759\
        );

    \I__3091\ : Span4Mux_h
    port map (
            O => \N__15762\,
            I => \N__15755\
        );

    \I__3090\ : Span4Mux_h
    port map (
            O => \N__15759\,
            I => \N__15752\
        );

    \I__3089\ : InMux
    port map (
            O => \N__15758\,
            I => \N__15748\
        );

    \I__3088\ : Sp12to4
    port map (
            O => \N__15755\,
            I => \N__15745\
        );

    \I__3087\ : Sp12to4
    port map (
            O => \N__15752\,
            I => \N__15742\
        );

    \I__3086\ : InMux
    port map (
            O => \N__15751\,
            I => \N__15739\
        );

    \I__3085\ : LocalMux
    port map (
            O => \N__15748\,
            I => \N__15736\
        );

    \I__3084\ : Span12Mux_v
    port map (
            O => \N__15745\,
            I => \N__15733\
        );

    \I__3083\ : Span12Mux_v
    port map (
            O => \N__15742\,
            I => \N__15730\
        );

    \I__3082\ : LocalMux
    port map (
            O => \N__15739\,
            I => \N__15725\
        );

    \I__3081\ : Span4Mux_v
    port map (
            O => \N__15736\,
            I => \N__15725\
        );

    \I__3080\ : Span12Mux_v
    port map (
            O => \N__15733\,
            I => \N__15720\
        );

    \I__3079\ : Span12Mux_v
    port map (
            O => \N__15730\,
            I => \N__15720\
        );

    \I__3078\ : Odrv4
    port map (
            O => \N__15725\,
            I => \RX_ADDR_1\
        );

    \I__3077\ : Odrv12
    port map (
            O => \N__15720\,
            I => \RX_ADDR_1\
        );

    \I__3076\ : InMux
    port map (
            O => \N__15715\,
            I => \N__15712\
        );

    \I__3075\ : LocalMux
    port map (
            O => \N__15712\,
            I => \N__15709\
        );

    \I__3074\ : Span4Mux_v
    port map (
            O => \N__15709\,
            I => \N__15706\
        );

    \I__3073\ : Span4Mux_h
    port map (
            O => \N__15706\,
            I => \N__15703\
        );

    \I__3072\ : Odrv4
    port map (
            O => \N__15703\,
            I => \line_buffer.n545\
        );

    \I__3071\ : InMux
    port map (
            O => \N__15700\,
            I => \N__15697\
        );

    \I__3070\ : LocalMux
    port map (
            O => \N__15697\,
            I => \N__15694\
        );

    \I__3069\ : Span4Mux_v
    port map (
            O => \N__15694\,
            I => \N__15691\
        );

    \I__3068\ : Sp12to4
    port map (
            O => \N__15691\,
            I => \N__15688\
        );

    \I__3067\ : Span12Mux_h
    port map (
            O => \N__15688\,
            I => \N__15685\
        );

    \I__3066\ : Span12Mux_v
    port map (
            O => \N__15685\,
            I => \N__15682\
        );

    \I__3065\ : Odrv12
    port map (
            O => \N__15682\,
            I => \line_buffer.n537\
        );

    \I__3064\ : InMux
    port map (
            O => \N__15679\,
            I => \N__15676\
        );

    \I__3063\ : LocalMux
    port map (
            O => \N__15676\,
            I => \line_buffer.n3680\
        );

    \I__3062\ : InMux
    port map (
            O => \N__15673\,
            I => \N__15670\
        );

    \I__3061\ : LocalMux
    port map (
            O => \N__15670\,
            I => \N__15667\
        );

    \I__3060\ : Span12Mux_s10_v
    port map (
            O => \N__15667\,
            I => \N__15664\
        );

    \I__3059\ : Odrv12
    port map (
            O => \N__15664\,
            I => \receive_module.n126\
        );

    \I__3058\ : CascadeMux
    port map (
            O => \N__15661\,
            I => \N__15658\
        );

    \I__3057\ : CascadeBuf
    port map (
            O => \N__15658\,
            I => \N__15654\
        );

    \I__3056\ : CascadeMux
    port map (
            O => \N__15657\,
            I => \N__15651\
        );

    \I__3055\ : CascadeMux
    port map (
            O => \N__15654\,
            I => \N__15648\
        );

    \I__3054\ : CascadeBuf
    port map (
            O => \N__15651\,
            I => \N__15645\
        );

    \I__3053\ : CascadeBuf
    port map (
            O => \N__15648\,
            I => \N__15642\
        );

    \I__3052\ : CascadeMux
    port map (
            O => \N__15645\,
            I => \N__15639\
        );

    \I__3051\ : CascadeMux
    port map (
            O => \N__15642\,
            I => \N__15636\
        );

    \I__3050\ : CascadeBuf
    port map (
            O => \N__15639\,
            I => \N__15633\
        );

    \I__3049\ : CascadeBuf
    port map (
            O => \N__15636\,
            I => \N__15630\
        );

    \I__3048\ : CascadeMux
    port map (
            O => \N__15633\,
            I => \N__15627\
        );

    \I__3047\ : CascadeMux
    port map (
            O => \N__15630\,
            I => \N__15624\
        );

    \I__3046\ : CascadeBuf
    port map (
            O => \N__15627\,
            I => \N__15621\
        );

    \I__3045\ : CascadeBuf
    port map (
            O => \N__15624\,
            I => \N__15618\
        );

    \I__3044\ : CascadeMux
    port map (
            O => \N__15621\,
            I => \N__15615\
        );

    \I__3043\ : CascadeMux
    port map (
            O => \N__15618\,
            I => \N__15612\
        );

    \I__3042\ : CascadeBuf
    port map (
            O => \N__15615\,
            I => \N__15609\
        );

    \I__3041\ : CascadeBuf
    port map (
            O => \N__15612\,
            I => \N__15606\
        );

    \I__3040\ : CascadeMux
    port map (
            O => \N__15609\,
            I => \N__15603\
        );

    \I__3039\ : CascadeMux
    port map (
            O => \N__15606\,
            I => \N__15600\
        );

    \I__3038\ : CascadeBuf
    port map (
            O => \N__15603\,
            I => \N__15597\
        );

    \I__3037\ : CascadeBuf
    port map (
            O => \N__15600\,
            I => \N__15594\
        );

    \I__3036\ : CascadeMux
    port map (
            O => \N__15597\,
            I => \N__15591\
        );

    \I__3035\ : CascadeMux
    port map (
            O => \N__15594\,
            I => \N__15588\
        );

    \I__3034\ : CascadeBuf
    port map (
            O => \N__15591\,
            I => \N__15585\
        );

    \I__3033\ : CascadeBuf
    port map (
            O => \N__15588\,
            I => \N__15582\
        );

    \I__3032\ : CascadeMux
    port map (
            O => \N__15585\,
            I => \N__15579\
        );

    \I__3031\ : CascadeMux
    port map (
            O => \N__15582\,
            I => \N__15576\
        );

    \I__3030\ : CascadeBuf
    port map (
            O => \N__15579\,
            I => \N__15573\
        );

    \I__3029\ : CascadeBuf
    port map (
            O => \N__15576\,
            I => \N__15570\
        );

    \I__3028\ : CascadeMux
    port map (
            O => \N__15573\,
            I => \N__15567\
        );

    \I__3027\ : CascadeMux
    port map (
            O => \N__15570\,
            I => \N__15564\
        );

    \I__3026\ : CascadeBuf
    port map (
            O => \N__15567\,
            I => \N__15561\
        );

    \I__3025\ : CascadeBuf
    port map (
            O => \N__15564\,
            I => \N__15558\
        );

    \I__3024\ : CascadeMux
    port map (
            O => \N__15561\,
            I => \N__15555\
        );

    \I__3023\ : CascadeMux
    port map (
            O => \N__15558\,
            I => \N__15552\
        );

    \I__3022\ : CascadeBuf
    port map (
            O => \N__15555\,
            I => \N__15549\
        );

    \I__3021\ : CascadeBuf
    port map (
            O => \N__15552\,
            I => \N__15546\
        );

    \I__3020\ : CascadeMux
    port map (
            O => \N__15549\,
            I => \N__15543\
        );

    \I__3019\ : CascadeMux
    port map (
            O => \N__15546\,
            I => \N__15540\
        );

    \I__3018\ : CascadeBuf
    port map (
            O => \N__15543\,
            I => \N__15537\
        );

    \I__3017\ : CascadeBuf
    port map (
            O => \N__15540\,
            I => \N__15534\
        );

    \I__3016\ : CascadeMux
    port map (
            O => \N__15537\,
            I => \N__15531\
        );

    \I__3015\ : CascadeMux
    port map (
            O => \N__15534\,
            I => \N__15528\
        );

    \I__3014\ : CascadeBuf
    port map (
            O => \N__15531\,
            I => \N__15525\
        );

    \I__3013\ : CascadeBuf
    port map (
            O => \N__15528\,
            I => \N__15522\
        );

    \I__3012\ : CascadeMux
    port map (
            O => \N__15525\,
            I => \N__15519\
        );

    \I__3011\ : CascadeMux
    port map (
            O => \N__15522\,
            I => \N__15516\
        );

    \I__3010\ : CascadeBuf
    port map (
            O => \N__15519\,
            I => \N__15513\
        );

    \I__3009\ : CascadeBuf
    port map (
            O => \N__15516\,
            I => \N__15510\
        );

    \I__3008\ : CascadeMux
    port map (
            O => \N__15513\,
            I => \N__15507\
        );

    \I__3007\ : CascadeMux
    port map (
            O => \N__15510\,
            I => \N__15504\
        );

    \I__3006\ : CascadeBuf
    port map (
            O => \N__15507\,
            I => \N__15501\
        );

    \I__3005\ : CascadeBuf
    port map (
            O => \N__15504\,
            I => \N__15498\
        );

    \I__3004\ : CascadeMux
    port map (
            O => \N__15501\,
            I => \N__15495\
        );

    \I__3003\ : CascadeMux
    port map (
            O => \N__15498\,
            I => \N__15492\
        );

    \I__3002\ : CascadeBuf
    port map (
            O => \N__15495\,
            I => \N__15489\
        );

    \I__3001\ : CascadeBuf
    port map (
            O => \N__15492\,
            I => \N__15486\
        );

    \I__3000\ : CascadeMux
    port map (
            O => \N__15489\,
            I => \N__15483\
        );

    \I__2999\ : CascadeMux
    port map (
            O => \N__15486\,
            I => \N__15480\
        );

    \I__2998\ : CascadeBuf
    port map (
            O => \N__15483\,
            I => \N__15476\
        );

    \I__2997\ : InMux
    port map (
            O => \N__15480\,
            I => \N__15473\
        );

    \I__2996\ : InMux
    port map (
            O => \N__15479\,
            I => \N__15470\
        );

    \I__2995\ : CascadeMux
    port map (
            O => \N__15476\,
            I => \N__15467\
        );

    \I__2994\ : LocalMux
    port map (
            O => \N__15473\,
            I => \N__15464\
        );

    \I__2993\ : LocalMux
    port map (
            O => \N__15470\,
            I => \N__15461\
        );

    \I__2992\ : InMux
    port map (
            O => \N__15467\,
            I => \N__15458\
        );

    \I__2991\ : Span4Mux_s1_v
    port map (
            O => \N__15464\,
            I => \N__15455\
        );

    \I__2990\ : Span4Mux_h
    port map (
            O => \N__15461\,
            I => \N__15452\
        );

    \I__2989\ : LocalMux
    port map (
            O => \N__15458\,
            I => \N__15449\
        );

    \I__2988\ : Span4Mux_h
    port map (
            O => \N__15455\,
            I => \N__15446\
        );

    \I__2987\ : Span4Mux_v
    port map (
            O => \N__15452\,
            I => \N__15443\
        );

    \I__2986\ : Sp12to4
    port map (
            O => \N__15449\,
            I => \N__15439\
        );

    \I__2985\ : Span4Mux_v
    port map (
            O => \N__15446\,
            I => \N__15436\
        );

    \I__2984\ : Span4Mux_v
    port map (
            O => \N__15443\,
            I => \N__15433\
        );

    \I__2983\ : InMux
    port map (
            O => \N__15442\,
            I => \N__15430\
        );

    \I__2982\ : Span12Mux_s9_v
    port map (
            O => \N__15439\,
            I => \N__15427\
        );

    \I__2981\ : Span4Mux_v
    port map (
            O => \N__15436\,
            I => \N__15424\
        );

    \I__2980\ : Odrv4
    port map (
            O => \N__15433\,
            I => \RX_ADDR_10\
        );

    \I__2979\ : LocalMux
    port map (
            O => \N__15430\,
            I => \RX_ADDR_10\
        );

    \I__2978\ : Odrv12
    port map (
            O => \N__15427\,
            I => \RX_ADDR_10\
        );

    \I__2977\ : Odrv4
    port map (
            O => \N__15424\,
            I => \RX_ADDR_10\
        );

    \I__2976\ : InMux
    port map (
            O => \N__15415\,
            I => \N__15412\
        );

    \I__2975\ : LocalMux
    port map (
            O => \N__15412\,
            I => \N__15409\
        );

    \I__2974\ : Span12Mux_s5_v
    port map (
            O => \N__15409\,
            I => \N__15406\
        );

    \I__2973\ : Span12Mux_v
    port map (
            O => \N__15406\,
            I => \N__15403\
        );

    \I__2972\ : Odrv12
    port map (
            O => \N__15403\,
            I => \receive_module.n132\
        );

    \I__2971\ : CascadeMux
    port map (
            O => \N__15400\,
            I => \N__15396\
        );

    \I__2970\ : CascadeMux
    port map (
            O => \N__15399\,
            I => \N__15393\
        );

    \I__2969\ : CascadeBuf
    port map (
            O => \N__15396\,
            I => \N__15390\
        );

    \I__2968\ : CascadeBuf
    port map (
            O => \N__15393\,
            I => \N__15387\
        );

    \I__2967\ : CascadeMux
    port map (
            O => \N__15390\,
            I => \N__15384\
        );

    \I__2966\ : CascadeMux
    port map (
            O => \N__15387\,
            I => \N__15381\
        );

    \I__2965\ : CascadeBuf
    port map (
            O => \N__15384\,
            I => \N__15378\
        );

    \I__2964\ : CascadeBuf
    port map (
            O => \N__15381\,
            I => \N__15375\
        );

    \I__2963\ : CascadeMux
    port map (
            O => \N__15378\,
            I => \N__15372\
        );

    \I__2962\ : CascadeMux
    port map (
            O => \N__15375\,
            I => \N__15369\
        );

    \I__2961\ : CascadeBuf
    port map (
            O => \N__15372\,
            I => \N__15366\
        );

    \I__2960\ : CascadeBuf
    port map (
            O => \N__15369\,
            I => \N__15363\
        );

    \I__2959\ : CascadeMux
    port map (
            O => \N__15366\,
            I => \N__15360\
        );

    \I__2958\ : CascadeMux
    port map (
            O => \N__15363\,
            I => \N__15357\
        );

    \I__2957\ : CascadeBuf
    port map (
            O => \N__15360\,
            I => \N__15354\
        );

    \I__2956\ : CascadeBuf
    port map (
            O => \N__15357\,
            I => \N__15351\
        );

    \I__2955\ : CascadeMux
    port map (
            O => \N__15354\,
            I => \N__15348\
        );

    \I__2954\ : CascadeMux
    port map (
            O => \N__15351\,
            I => \N__15345\
        );

    \I__2953\ : CascadeBuf
    port map (
            O => \N__15348\,
            I => \N__15342\
        );

    \I__2952\ : CascadeBuf
    port map (
            O => \N__15345\,
            I => \N__15339\
        );

    \I__2951\ : CascadeMux
    port map (
            O => \N__15342\,
            I => \N__15336\
        );

    \I__2950\ : CascadeMux
    port map (
            O => \N__15339\,
            I => \N__15333\
        );

    \I__2949\ : CascadeBuf
    port map (
            O => \N__15336\,
            I => \N__15330\
        );

    \I__2948\ : CascadeBuf
    port map (
            O => \N__15333\,
            I => \N__15327\
        );

    \I__2947\ : CascadeMux
    port map (
            O => \N__15330\,
            I => \N__15324\
        );

    \I__2946\ : CascadeMux
    port map (
            O => \N__15327\,
            I => \N__15321\
        );

    \I__2945\ : CascadeBuf
    port map (
            O => \N__15324\,
            I => \N__15318\
        );

    \I__2944\ : CascadeBuf
    port map (
            O => \N__15321\,
            I => \N__15315\
        );

    \I__2943\ : CascadeMux
    port map (
            O => \N__15318\,
            I => \N__15312\
        );

    \I__2942\ : CascadeMux
    port map (
            O => \N__15315\,
            I => \N__15309\
        );

    \I__2941\ : CascadeBuf
    port map (
            O => \N__15312\,
            I => \N__15306\
        );

    \I__2940\ : CascadeBuf
    port map (
            O => \N__15309\,
            I => \N__15303\
        );

    \I__2939\ : CascadeMux
    port map (
            O => \N__15306\,
            I => \N__15300\
        );

    \I__2938\ : CascadeMux
    port map (
            O => \N__15303\,
            I => \N__15297\
        );

    \I__2937\ : CascadeBuf
    port map (
            O => \N__15300\,
            I => \N__15294\
        );

    \I__2936\ : CascadeBuf
    port map (
            O => \N__15297\,
            I => \N__15291\
        );

    \I__2935\ : CascadeMux
    port map (
            O => \N__15294\,
            I => \N__15288\
        );

    \I__2934\ : CascadeMux
    port map (
            O => \N__15291\,
            I => \N__15285\
        );

    \I__2933\ : CascadeBuf
    port map (
            O => \N__15288\,
            I => \N__15282\
        );

    \I__2932\ : CascadeBuf
    port map (
            O => \N__15285\,
            I => \N__15279\
        );

    \I__2931\ : CascadeMux
    port map (
            O => \N__15282\,
            I => \N__15276\
        );

    \I__2930\ : CascadeMux
    port map (
            O => \N__15279\,
            I => \N__15273\
        );

    \I__2929\ : CascadeBuf
    port map (
            O => \N__15276\,
            I => \N__15270\
        );

    \I__2928\ : CascadeBuf
    port map (
            O => \N__15273\,
            I => \N__15267\
        );

    \I__2927\ : CascadeMux
    port map (
            O => \N__15270\,
            I => \N__15264\
        );

    \I__2926\ : CascadeMux
    port map (
            O => \N__15267\,
            I => \N__15261\
        );

    \I__2925\ : CascadeBuf
    port map (
            O => \N__15264\,
            I => \N__15258\
        );

    \I__2924\ : CascadeBuf
    port map (
            O => \N__15261\,
            I => \N__15255\
        );

    \I__2923\ : CascadeMux
    port map (
            O => \N__15258\,
            I => \N__15252\
        );

    \I__2922\ : CascadeMux
    port map (
            O => \N__15255\,
            I => \N__15249\
        );

    \I__2921\ : CascadeBuf
    port map (
            O => \N__15252\,
            I => \N__15246\
        );

    \I__2920\ : CascadeBuf
    port map (
            O => \N__15249\,
            I => \N__15243\
        );

    \I__2919\ : CascadeMux
    port map (
            O => \N__15246\,
            I => \N__15240\
        );

    \I__2918\ : CascadeMux
    port map (
            O => \N__15243\,
            I => \N__15237\
        );

    \I__2917\ : CascadeBuf
    port map (
            O => \N__15240\,
            I => \N__15234\
        );

    \I__2916\ : CascadeBuf
    port map (
            O => \N__15237\,
            I => \N__15231\
        );

    \I__2915\ : CascadeMux
    port map (
            O => \N__15234\,
            I => \N__15228\
        );

    \I__2914\ : CascadeMux
    port map (
            O => \N__15231\,
            I => \N__15225\
        );

    \I__2913\ : CascadeBuf
    port map (
            O => \N__15228\,
            I => \N__15222\
        );

    \I__2912\ : CascadeBuf
    port map (
            O => \N__15225\,
            I => \N__15219\
        );

    \I__2911\ : CascadeMux
    port map (
            O => \N__15222\,
            I => \N__15215\
        );

    \I__2910\ : CascadeMux
    port map (
            O => \N__15219\,
            I => \N__15212\
        );

    \I__2909\ : InMux
    port map (
            O => \N__15218\,
            I => \N__15209\
        );

    \I__2908\ : InMux
    port map (
            O => \N__15215\,
            I => \N__15206\
        );

    \I__2907\ : InMux
    port map (
            O => \N__15212\,
            I => \N__15203\
        );

    \I__2906\ : LocalMux
    port map (
            O => \N__15209\,
            I => \N__15199\
        );

    \I__2905\ : LocalMux
    port map (
            O => \N__15206\,
            I => \N__15196\
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__15203\,
            I => \N__15193\
        );

    \I__2903\ : InMux
    port map (
            O => \N__15202\,
            I => \N__15190\
        );

    \I__2902\ : Span12Mux_v
    port map (
            O => \N__15199\,
            I => \N__15183\
        );

    \I__2901\ : Span12Mux_h
    port map (
            O => \N__15196\,
            I => \N__15183\
        );

    \I__2900\ : Span12Mux_h
    port map (
            O => \N__15193\,
            I => \N__15183\
        );

    \I__2899\ : LocalMux
    port map (
            O => \N__15190\,
            I => \RX_ADDR_4\
        );

    \I__2898\ : Odrv12
    port map (
            O => \N__15183\,
            I => \RX_ADDR_4\
        );

    \I__2897\ : InMux
    port map (
            O => \N__15178\,
            I => \N__15175\
        );

    \I__2896\ : LocalMux
    port map (
            O => \N__15175\,
            I => \N__15172\
        );

    \I__2895\ : Span12Mux_s4_v
    port map (
            O => \N__15172\,
            I => \N__15169\
        );

    \I__2894\ : Span12Mux_v
    port map (
            O => \N__15169\,
            I => \N__15166\
        );

    \I__2893\ : Odrv12
    port map (
            O => \N__15166\,
            I => \receive_module.n131\
        );

    \I__2892\ : CascadeMux
    port map (
            O => \N__15163\,
            I => \N__15159\
        );

    \I__2891\ : CascadeMux
    port map (
            O => \N__15162\,
            I => \N__15156\
        );

    \I__2890\ : CascadeBuf
    port map (
            O => \N__15159\,
            I => \N__15153\
        );

    \I__2889\ : CascadeBuf
    port map (
            O => \N__15156\,
            I => \N__15150\
        );

    \I__2888\ : CascadeMux
    port map (
            O => \N__15153\,
            I => \N__15147\
        );

    \I__2887\ : CascadeMux
    port map (
            O => \N__15150\,
            I => \N__15144\
        );

    \I__2886\ : CascadeBuf
    port map (
            O => \N__15147\,
            I => \N__15141\
        );

    \I__2885\ : CascadeBuf
    port map (
            O => \N__15144\,
            I => \N__15138\
        );

    \I__2884\ : CascadeMux
    port map (
            O => \N__15141\,
            I => \N__15135\
        );

    \I__2883\ : CascadeMux
    port map (
            O => \N__15138\,
            I => \N__15132\
        );

    \I__2882\ : CascadeBuf
    port map (
            O => \N__15135\,
            I => \N__15129\
        );

    \I__2881\ : CascadeBuf
    port map (
            O => \N__15132\,
            I => \N__15126\
        );

    \I__2880\ : CascadeMux
    port map (
            O => \N__15129\,
            I => \N__15123\
        );

    \I__2879\ : CascadeMux
    port map (
            O => \N__15126\,
            I => \N__15120\
        );

    \I__2878\ : CascadeBuf
    port map (
            O => \N__15123\,
            I => \N__15117\
        );

    \I__2877\ : CascadeBuf
    port map (
            O => \N__15120\,
            I => \N__15114\
        );

    \I__2876\ : CascadeMux
    port map (
            O => \N__15117\,
            I => \N__15111\
        );

    \I__2875\ : CascadeMux
    port map (
            O => \N__15114\,
            I => \N__15108\
        );

    \I__2874\ : CascadeBuf
    port map (
            O => \N__15111\,
            I => \N__15105\
        );

    \I__2873\ : CascadeBuf
    port map (
            O => \N__15108\,
            I => \N__15102\
        );

    \I__2872\ : CascadeMux
    port map (
            O => \N__15105\,
            I => \N__15099\
        );

    \I__2871\ : CascadeMux
    port map (
            O => \N__15102\,
            I => \N__15096\
        );

    \I__2870\ : CascadeBuf
    port map (
            O => \N__15099\,
            I => \N__15093\
        );

    \I__2869\ : CascadeBuf
    port map (
            O => \N__15096\,
            I => \N__15090\
        );

    \I__2868\ : CascadeMux
    port map (
            O => \N__15093\,
            I => \N__15087\
        );

    \I__2867\ : CascadeMux
    port map (
            O => \N__15090\,
            I => \N__15084\
        );

    \I__2866\ : CascadeBuf
    port map (
            O => \N__15087\,
            I => \N__15081\
        );

    \I__2865\ : CascadeBuf
    port map (
            O => \N__15084\,
            I => \N__15078\
        );

    \I__2864\ : CascadeMux
    port map (
            O => \N__15081\,
            I => \N__15075\
        );

    \I__2863\ : CascadeMux
    port map (
            O => \N__15078\,
            I => \N__15072\
        );

    \I__2862\ : CascadeBuf
    port map (
            O => \N__15075\,
            I => \N__15069\
        );

    \I__2861\ : CascadeBuf
    port map (
            O => \N__15072\,
            I => \N__15066\
        );

    \I__2860\ : CascadeMux
    port map (
            O => \N__15069\,
            I => \N__15063\
        );

    \I__2859\ : CascadeMux
    port map (
            O => \N__15066\,
            I => \N__15060\
        );

    \I__2858\ : CascadeBuf
    port map (
            O => \N__15063\,
            I => \N__15057\
        );

    \I__2857\ : CascadeBuf
    port map (
            O => \N__15060\,
            I => \N__15054\
        );

    \I__2856\ : CascadeMux
    port map (
            O => \N__15057\,
            I => \N__15051\
        );

    \I__2855\ : CascadeMux
    port map (
            O => \N__15054\,
            I => \N__15048\
        );

    \I__2854\ : CascadeBuf
    port map (
            O => \N__15051\,
            I => \N__15045\
        );

    \I__2853\ : CascadeBuf
    port map (
            O => \N__15048\,
            I => \N__15042\
        );

    \I__2852\ : CascadeMux
    port map (
            O => \N__15045\,
            I => \N__15039\
        );

    \I__2851\ : CascadeMux
    port map (
            O => \N__15042\,
            I => \N__15036\
        );

    \I__2850\ : CascadeBuf
    port map (
            O => \N__15039\,
            I => \N__15033\
        );

    \I__2849\ : CascadeBuf
    port map (
            O => \N__15036\,
            I => \N__15030\
        );

    \I__2848\ : CascadeMux
    port map (
            O => \N__15033\,
            I => \N__15027\
        );

    \I__2847\ : CascadeMux
    port map (
            O => \N__15030\,
            I => \N__15024\
        );

    \I__2846\ : CascadeBuf
    port map (
            O => \N__15027\,
            I => \N__15021\
        );

    \I__2845\ : CascadeBuf
    port map (
            O => \N__15024\,
            I => \N__15018\
        );

    \I__2844\ : CascadeMux
    port map (
            O => \N__15021\,
            I => \N__15015\
        );

    \I__2843\ : CascadeMux
    port map (
            O => \N__15018\,
            I => \N__15012\
        );

    \I__2842\ : CascadeBuf
    port map (
            O => \N__15015\,
            I => \N__15009\
        );

    \I__2841\ : CascadeBuf
    port map (
            O => \N__15012\,
            I => \N__15006\
        );

    \I__2840\ : CascadeMux
    port map (
            O => \N__15009\,
            I => \N__15003\
        );

    \I__2839\ : CascadeMux
    port map (
            O => \N__15006\,
            I => \N__15000\
        );

    \I__2838\ : CascadeBuf
    port map (
            O => \N__15003\,
            I => \N__14997\
        );

    \I__2837\ : CascadeBuf
    port map (
            O => \N__15000\,
            I => \N__14994\
        );

    \I__2836\ : CascadeMux
    port map (
            O => \N__14997\,
            I => \N__14991\
        );

    \I__2835\ : CascadeMux
    port map (
            O => \N__14994\,
            I => \N__14987\
        );

    \I__2834\ : CascadeBuf
    port map (
            O => \N__14991\,
            I => \N__14984\
        );

    \I__2833\ : InMux
    port map (
            O => \N__14990\,
            I => \N__14981\
        );

    \I__2832\ : CascadeBuf
    port map (
            O => \N__14987\,
            I => \N__14978\
        );

    \I__2831\ : CascadeMux
    port map (
            O => \N__14984\,
            I => \N__14975\
        );

    \I__2830\ : LocalMux
    port map (
            O => \N__14981\,
            I => \N__14972\
        );

    \I__2829\ : CascadeMux
    port map (
            O => \N__14978\,
            I => \N__14969\
        );

    \I__2828\ : InMux
    port map (
            O => \N__14975\,
            I => \N__14966\
        );

    \I__2827\ : Span4Mux_v
    port map (
            O => \N__14972\,
            I => \N__14963\
        );

    \I__2826\ : InMux
    port map (
            O => \N__14969\,
            I => \N__14960\
        );

    \I__2825\ : LocalMux
    port map (
            O => \N__14966\,
            I => \N__14957\
        );

    \I__2824\ : Span4Mux_v
    port map (
            O => \N__14963\,
            I => \N__14953\
        );

    \I__2823\ : LocalMux
    port map (
            O => \N__14960\,
            I => \N__14950\
        );

    \I__2822\ : Span4Mux_s1_v
    port map (
            O => \N__14957\,
            I => \N__14947\
        );

    \I__2821\ : CascadeMux
    port map (
            O => \N__14956\,
            I => \N__14944\
        );

    \I__2820\ : Span4Mux_v
    port map (
            O => \N__14953\,
            I => \N__14941\
        );

    \I__2819\ : Span4Mux_s1_v
    port map (
            O => \N__14950\,
            I => \N__14938\
        );

    \I__2818\ : Span4Mux_h
    port map (
            O => \N__14947\,
            I => \N__14935\
        );

    \I__2817\ : InMux
    port map (
            O => \N__14944\,
            I => \N__14932\
        );

    \I__2816\ : Sp12to4
    port map (
            O => \N__14941\,
            I => \N__14929\
        );

    \I__2815\ : Span4Mux_h
    port map (
            O => \N__14938\,
            I => \N__14926\
        );

    \I__2814\ : Span4Mux_h
    port map (
            O => \N__14935\,
            I => \N__14923\
        );

    \I__2813\ : LocalMux
    port map (
            O => \N__14932\,
            I => \RX_ADDR_5\
        );

    \I__2812\ : Odrv12
    port map (
            O => \N__14929\,
            I => \RX_ADDR_5\
        );

    \I__2811\ : Odrv4
    port map (
            O => \N__14926\,
            I => \RX_ADDR_5\
        );

    \I__2810\ : Odrv4
    port map (
            O => \N__14923\,
            I => \RX_ADDR_5\
        );

    \I__2809\ : InMux
    port map (
            O => \N__14914\,
            I => \N__14911\
        );

    \I__2808\ : LocalMux
    port map (
            O => \N__14911\,
            I => \N__14908\
        );

    \I__2807\ : Span12Mux_s3_v
    port map (
            O => \N__14908\,
            I => \N__14905\
        );

    \I__2806\ : Span12Mux_v
    port map (
            O => \N__14905\,
            I => \N__14902\
        );

    \I__2805\ : Odrv12
    port map (
            O => \N__14902\,
            I => \receive_module.n130\
        );

    \I__2804\ : CascadeMux
    port map (
            O => \N__14899\,
            I => \N__14896\
        );

    \I__2803\ : CascadeBuf
    port map (
            O => \N__14896\,
            I => \N__14892\
        );

    \I__2802\ : CascadeMux
    port map (
            O => \N__14895\,
            I => \N__14889\
        );

    \I__2801\ : CascadeMux
    port map (
            O => \N__14892\,
            I => \N__14886\
        );

    \I__2800\ : CascadeBuf
    port map (
            O => \N__14889\,
            I => \N__14883\
        );

    \I__2799\ : CascadeBuf
    port map (
            O => \N__14886\,
            I => \N__14880\
        );

    \I__2798\ : CascadeMux
    port map (
            O => \N__14883\,
            I => \N__14877\
        );

    \I__2797\ : CascadeMux
    port map (
            O => \N__14880\,
            I => \N__14874\
        );

    \I__2796\ : CascadeBuf
    port map (
            O => \N__14877\,
            I => \N__14871\
        );

    \I__2795\ : CascadeBuf
    port map (
            O => \N__14874\,
            I => \N__14868\
        );

    \I__2794\ : CascadeMux
    port map (
            O => \N__14871\,
            I => \N__14865\
        );

    \I__2793\ : CascadeMux
    port map (
            O => \N__14868\,
            I => \N__14862\
        );

    \I__2792\ : CascadeBuf
    port map (
            O => \N__14865\,
            I => \N__14859\
        );

    \I__2791\ : CascadeBuf
    port map (
            O => \N__14862\,
            I => \N__14856\
        );

    \I__2790\ : CascadeMux
    port map (
            O => \N__14859\,
            I => \N__14853\
        );

    \I__2789\ : CascadeMux
    port map (
            O => \N__14856\,
            I => \N__14850\
        );

    \I__2788\ : CascadeBuf
    port map (
            O => \N__14853\,
            I => \N__14847\
        );

    \I__2787\ : CascadeBuf
    port map (
            O => \N__14850\,
            I => \N__14844\
        );

    \I__2786\ : CascadeMux
    port map (
            O => \N__14847\,
            I => \N__14841\
        );

    \I__2785\ : CascadeMux
    port map (
            O => \N__14844\,
            I => \N__14838\
        );

    \I__2784\ : CascadeBuf
    port map (
            O => \N__14841\,
            I => \N__14835\
        );

    \I__2783\ : CascadeBuf
    port map (
            O => \N__14838\,
            I => \N__14832\
        );

    \I__2782\ : CascadeMux
    port map (
            O => \N__14835\,
            I => \N__14829\
        );

    \I__2781\ : CascadeMux
    port map (
            O => \N__14832\,
            I => \N__14826\
        );

    \I__2780\ : CascadeBuf
    port map (
            O => \N__14829\,
            I => \N__14823\
        );

    \I__2779\ : CascadeBuf
    port map (
            O => \N__14826\,
            I => \N__14820\
        );

    \I__2778\ : CascadeMux
    port map (
            O => \N__14823\,
            I => \N__14817\
        );

    \I__2777\ : CascadeMux
    port map (
            O => \N__14820\,
            I => \N__14814\
        );

    \I__2776\ : CascadeBuf
    port map (
            O => \N__14817\,
            I => \N__14811\
        );

    \I__2775\ : CascadeBuf
    port map (
            O => \N__14814\,
            I => \N__14808\
        );

    \I__2774\ : CascadeMux
    port map (
            O => \N__14811\,
            I => \N__14805\
        );

    \I__2773\ : CascadeMux
    port map (
            O => \N__14808\,
            I => \N__14802\
        );

    \I__2772\ : CascadeBuf
    port map (
            O => \N__14805\,
            I => \N__14799\
        );

    \I__2771\ : CascadeBuf
    port map (
            O => \N__14802\,
            I => \N__14796\
        );

    \I__2770\ : CascadeMux
    port map (
            O => \N__14799\,
            I => \N__14793\
        );

    \I__2769\ : CascadeMux
    port map (
            O => \N__14796\,
            I => \N__14790\
        );

    \I__2768\ : CascadeBuf
    port map (
            O => \N__14793\,
            I => \N__14787\
        );

    \I__2767\ : CascadeBuf
    port map (
            O => \N__14790\,
            I => \N__14784\
        );

    \I__2766\ : CascadeMux
    port map (
            O => \N__14787\,
            I => \N__14781\
        );

    \I__2765\ : CascadeMux
    port map (
            O => \N__14784\,
            I => \N__14778\
        );

    \I__2764\ : CascadeBuf
    port map (
            O => \N__14781\,
            I => \N__14775\
        );

    \I__2763\ : CascadeBuf
    port map (
            O => \N__14778\,
            I => \N__14772\
        );

    \I__2762\ : CascadeMux
    port map (
            O => \N__14775\,
            I => \N__14769\
        );

    \I__2761\ : CascadeMux
    port map (
            O => \N__14772\,
            I => \N__14766\
        );

    \I__2760\ : CascadeBuf
    port map (
            O => \N__14769\,
            I => \N__14763\
        );

    \I__2759\ : CascadeBuf
    port map (
            O => \N__14766\,
            I => \N__14760\
        );

    \I__2758\ : CascadeMux
    port map (
            O => \N__14763\,
            I => \N__14757\
        );

    \I__2757\ : CascadeMux
    port map (
            O => \N__14760\,
            I => \N__14754\
        );

    \I__2756\ : CascadeBuf
    port map (
            O => \N__14757\,
            I => \N__14751\
        );

    \I__2755\ : CascadeBuf
    port map (
            O => \N__14754\,
            I => \N__14748\
        );

    \I__2754\ : CascadeMux
    port map (
            O => \N__14751\,
            I => \N__14745\
        );

    \I__2753\ : CascadeMux
    port map (
            O => \N__14748\,
            I => \N__14742\
        );

    \I__2752\ : CascadeBuf
    port map (
            O => \N__14745\,
            I => \N__14739\
        );

    \I__2751\ : CascadeBuf
    port map (
            O => \N__14742\,
            I => \N__14736\
        );

    \I__2750\ : CascadeMux
    port map (
            O => \N__14739\,
            I => \N__14733\
        );

    \I__2749\ : CascadeMux
    port map (
            O => \N__14736\,
            I => \N__14730\
        );

    \I__2748\ : CascadeBuf
    port map (
            O => \N__14733\,
            I => \N__14727\
        );

    \I__2747\ : CascadeBuf
    port map (
            O => \N__14730\,
            I => \N__14724\
        );

    \I__2746\ : CascadeMux
    port map (
            O => \N__14727\,
            I => \N__14721\
        );

    \I__2745\ : CascadeMux
    port map (
            O => \N__14724\,
            I => \N__14718\
        );

    \I__2744\ : CascadeBuf
    port map (
            O => \N__14721\,
            I => \N__14715\
        );

    \I__2743\ : InMux
    port map (
            O => \N__14718\,
            I => \N__14711\
        );

    \I__2742\ : CascadeMux
    port map (
            O => \N__14715\,
            I => \N__14708\
        );

    \I__2741\ : CascadeMux
    port map (
            O => \N__14714\,
            I => \N__14705\
        );

    \I__2740\ : LocalMux
    port map (
            O => \N__14711\,
            I => \N__14702\
        );

    \I__2739\ : InMux
    port map (
            O => \N__14708\,
            I => \N__14699\
        );

    \I__2738\ : InMux
    port map (
            O => \N__14705\,
            I => \N__14696\
        );

    \I__2737\ : Span4Mux_h
    port map (
            O => \N__14702\,
            I => \N__14693\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__14699\,
            I => \N__14690\
        );

    \I__2735\ : LocalMux
    port map (
            O => \N__14696\,
            I => \N__14687\
        );

    \I__2734\ : Span4Mux_h
    port map (
            O => \N__14693\,
            I => \N__14683\
        );

    \I__2733\ : Span4Mux_h
    port map (
            O => \N__14690\,
            I => \N__14680\
        );

    \I__2732\ : Span12Mux_v
    port map (
            O => \N__14687\,
            I => \N__14677\
        );

    \I__2731\ : InMux
    port map (
            O => \N__14686\,
            I => \N__14674\
        );

    \I__2730\ : Span4Mux_h
    port map (
            O => \N__14683\,
            I => \N__14669\
        );

    \I__2729\ : Span4Mux_h
    port map (
            O => \N__14680\,
            I => \N__14669\
        );

    \I__2728\ : Odrv12
    port map (
            O => \N__14677\,
            I => \RX_ADDR_6\
        );

    \I__2727\ : LocalMux
    port map (
            O => \N__14674\,
            I => \RX_ADDR_6\
        );

    \I__2726\ : Odrv4
    port map (
            O => \N__14669\,
            I => \RX_ADDR_6\
        );

    \I__2725\ : InMux
    port map (
            O => \N__14662\,
            I => \N__14659\
        );

    \I__2724\ : LocalMux
    port map (
            O => \N__14659\,
            I => \N__14656\
        );

    \I__2723\ : Span12Mux_s2_v
    port map (
            O => \N__14656\,
            I => \N__14653\
        );

    \I__2722\ : Span12Mux_v
    port map (
            O => \N__14653\,
            I => \N__14650\
        );

    \I__2721\ : Odrv12
    port map (
            O => \N__14650\,
            I => \receive_module.n129\
        );

    \I__2720\ : CascadeMux
    port map (
            O => \N__14647\,
            I => \N__14643\
        );

    \I__2719\ : CascadeMux
    port map (
            O => \N__14646\,
            I => \N__14640\
        );

    \I__2718\ : CascadeBuf
    port map (
            O => \N__14643\,
            I => \N__14637\
        );

    \I__2717\ : CascadeBuf
    port map (
            O => \N__14640\,
            I => \N__14634\
        );

    \I__2716\ : CascadeMux
    port map (
            O => \N__14637\,
            I => \N__14631\
        );

    \I__2715\ : CascadeMux
    port map (
            O => \N__14634\,
            I => \N__14628\
        );

    \I__2714\ : CascadeBuf
    port map (
            O => \N__14631\,
            I => \N__14625\
        );

    \I__2713\ : CascadeBuf
    port map (
            O => \N__14628\,
            I => \N__14622\
        );

    \I__2712\ : CascadeMux
    port map (
            O => \N__14625\,
            I => \N__14619\
        );

    \I__2711\ : CascadeMux
    port map (
            O => \N__14622\,
            I => \N__14616\
        );

    \I__2710\ : CascadeBuf
    port map (
            O => \N__14619\,
            I => \N__14613\
        );

    \I__2709\ : CascadeBuf
    port map (
            O => \N__14616\,
            I => \N__14610\
        );

    \I__2708\ : CascadeMux
    port map (
            O => \N__14613\,
            I => \N__14607\
        );

    \I__2707\ : CascadeMux
    port map (
            O => \N__14610\,
            I => \N__14604\
        );

    \I__2706\ : CascadeBuf
    port map (
            O => \N__14607\,
            I => \N__14601\
        );

    \I__2705\ : CascadeBuf
    port map (
            O => \N__14604\,
            I => \N__14598\
        );

    \I__2704\ : CascadeMux
    port map (
            O => \N__14601\,
            I => \N__14595\
        );

    \I__2703\ : CascadeMux
    port map (
            O => \N__14598\,
            I => \N__14592\
        );

    \I__2702\ : CascadeBuf
    port map (
            O => \N__14595\,
            I => \N__14589\
        );

    \I__2701\ : CascadeBuf
    port map (
            O => \N__14592\,
            I => \N__14586\
        );

    \I__2700\ : CascadeMux
    port map (
            O => \N__14589\,
            I => \N__14583\
        );

    \I__2699\ : CascadeMux
    port map (
            O => \N__14586\,
            I => \N__14580\
        );

    \I__2698\ : CascadeBuf
    port map (
            O => \N__14583\,
            I => \N__14577\
        );

    \I__2697\ : CascadeBuf
    port map (
            O => \N__14580\,
            I => \N__14574\
        );

    \I__2696\ : CascadeMux
    port map (
            O => \N__14577\,
            I => \N__14571\
        );

    \I__2695\ : CascadeMux
    port map (
            O => \N__14574\,
            I => \N__14568\
        );

    \I__2694\ : CascadeBuf
    port map (
            O => \N__14571\,
            I => \N__14565\
        );

    \I__2693\ : CascadeBuf
    port map (
            O => \N__14568\,
            I => \N__14562\
        );

    \I__2692\ : CascadeMux
    port map (
            O => \N__14565\,
            I => \N__14559\
        );

    \I__2691\ : CascadeMux
    port map (
            O => \N__14562\,
            I => \N__14556\
        );

    \I__2690\ : CascadeBuf
    port map (
            O => \N__14559\,
            I => \N__14553\
        );

    \I__2689\ : CascadeBuf
    port map (
            O => \N__14556\,
            I => \N__14550\
        );

    \I__2688\ : CascadeMux
    port map (
            O => \N__14553\,
            I => \N__14547\
        );

    \I__2687\ : CascadeMux
    port map (
            O => \N__14550\,
            I => \N__14544\
        );

    \I__2686\ : CascadeBuf
    port map (
            O => \N__14547\,
            I => \N__14541\
        );

    \I__2685\ : CascadeBuf
    port map (
            O => \N__14544\,
            I => \N__14538\
        );

    \I__2684\ : CascadeMux
    port map (
            O => \N__14541\,
            I => \N__14535\
        );

    \I__2683\ : CascadeMux
    port map (
            O => \N__14538\,
            I => \N__14532\
        );

    \I__2682\ : CascadeBuf
    port map (
            O => \N__14535\,
            I => \N__14529\
        );

    \I__2681\ : CascadeBuf
    port map (
            O => \N__14532\,
            I => \N__14526\
        );

    \I__2680\ : CascadeMux
    port map (
            O => \N__14529\,
            I => \N__14523\
        );

    \I__2679\ : CascadeMux
    port map (
            O => \N__14526\,
            I => \N__14520\
        );

    \I__2678\ : CascadeBuf
    port map (
            O => \N__14523\,
            I => \N__14517\
        );

    \I__2677\ : CascadeBuf
    port map (
            O => \N__14520\,
            I => \N__14514\
        );

    \I__2676\ : CascadeMux
    port map (
            O => \N__14517\,
            I => \N__14511\
        );

    \I__2675\ : CascadeMux
    port map (
            O => \N__14514\,
            I => \N__14508\
        );

    \I__2674\ : CascadeBuf
    port map (
            O => \N__14511\,
            I => \N__14505\
        );

    \I__2673\ : CascadeBuf
    port map (
            O => \N__14508\,
            I => \N__14502\
        );

    \I__2672\ : CascadeMux
    port map (
            O => \N__14505\,
            I => \N__14499\
        );

    \I__2671\ : CascadeMux
    port map (
            O => \N__14502\,
            I => \N__14496\
        );

    \I__2670\ : CascadeBuf
    port map (
            O => \N__14499\,
            I => \N__14493\
        );

    \I__2669\ : CascadeBuf
    port map (
            O => \N__14496\,
            I => \N__14490\
        );

    \I__2668\ : CascadeMux
    port map (
            O => \N__14493\,
            I => \N__14487\
        );

    \I__2667\ : CascadeMux
    port map (
            O => \N__14490\,
            I => \N__14484\
        );

    \I__2666\ : CascadeBuf
    port map (
            O => \N__14487\,
            I => \N__14481\
        );

    \I__2665\ : CascadeBuf
    port map (
            O => \N__14484\,
            I => \N__14478\
        );

    \I__2664\ : CascadeMux
    port map (
            O => \N__14481\,
            I => \N__14475\
        );

    \I__2663\ : CascadeMux
    port map (
            O => \N__14478\,
            I => \N__14472\
        );

    \I__2662\ : CascadeBuf
    port map (
            O => \N__14475\,
            I => \N__14469\
        );

    \I__2661\ : CascadeBuf
    port map (
            O => \N__14472\,
            I => \N__14466\
        );

    \I__2660\ : CascadeMux
    port map (
            O => \N__14469\,
            I => \N__14463\
        );

    \I__2659\ : CascadeMux
    port map (
            O => \N__14466\,
            I => \N__14459\
        );

    \I__2658\ : InMux
    port map (
            O => \N__14463\,
            I => \N__14456\
        );

    \I__2657\ : InMux
    port map (
            O => \N__14462\,
            I => \N__14453\
        );

    \I__2656\ : InMux
    port map (
            O => \N__14459\,
            I => \N__14450\
        );

    \I__2655\ : LocalMux
    port map (
            O => \N__14456\,
            I => \N__14447\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__14453\,
            I => \N__14443\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__14450\,
            I => \N__14440\
        );

    \I__2652\ : Span4Mux_s1_v
    port map (
            O => \N__14447\,
            I => \N__14437\
        );

    \I__2651\ : CascadeMux
    port map (
            O => \N__14446\,
            I => \N__14434\
        );

    \I__2650\ : Span12Mux_v
    port map (
            O => \N__14443\,
            I => \N__14431\
        );

    \I__2649\ : Span4Mux_s1_v
    port map (
            O => \N__14440\,
            I => \N__14428\
        );

    \I__2648\ : Span4Mux_h
    port map (
            O => \N__14437\,
            I => \N__14425\
        );

    \I__2647\ : InMux
    port map (
            O => \N__14434\,
            I => \N__14422\
        );

    \I__2646\ : Span12Mux_v
    port map (
            O => \N__14431\,
            I => \N__14419\
        );

    \I__2645\ : Span4Mux_h
    port map (
            O => \N__14428\,
            I => \N__14414\
        );

    \I__2644\ : Span4Mux_h
    port map (
            O => \N__14425\,
            I => \N__14414\
        );

    \I__2643\ : LocalMux
    port map (
            O => \N__14422\,
            I => \RX_ADDR_7\
        );

    \I__2642\ : Odrv12
    port map (
            O => \N__14419\,
            I => \RX_ADDR_7\
        );

    \I__2641\ : Odrv4
    port map (
            O => \N__14414\,
            I => \RX_ADDR_7\
        );

    \I__2640\ : InMux
    port map (
            O => \N__14407\,
            I => \N__14404\
        );

    \I__2639\ : LocalMux
    port map (
            O => \N__14404\,
            I => \N__14401\
        );

    \I__2638\ : Span12Mux_v
    port map (
            O => \N__14401\,
            I => \N__14398\
        );

    \I__2637\ : Odrv12
    port map (
            O => \N__14398\,
            I => \receive_module.n128\
        );

    \I__2636\ : CascadeMux
    port map (
            O => \N__14395\,
            I => \N__14392\
        );

    \I__2635\ : CascadeBuf
    port map (
            O => \N__14392\,
            I => \N__14388\
        );

    \I__2634\ : CascadeMux
    port map (
            O => \N__14391\,
            I => \N__14385\
        );

    \I__2633\ : CascadeMux
    port map (
            O => \N__14388\,
            I => \N__14382\
        );

    \I__2632\ : CascadeBuf
    port map (
            O => \N__14385\,
            I => \N__14379\
        );

    \I__2631\ : CascadeBuf
    port map (
            O => \N__14382\,
            I => \N__14376\
        );

    \I__2630\ : CascadeMux
    port map (
            O => \N__14379\,
            I => \N__14373\
        );

    \I__2629\ : CascadeMux
    port map (
            O => \N__14376\,
            I => \N__14370\
        );

    \I__2628\ : CascadeBuf
    port map (
            O => \N__14373\,
            I => \N__14367\
        );

    \I__2627\ : CascadeBuf
    port map (
            O => \N__14370\,
            I => \N__14364\
        );

    \I__2626\ : CascadeMux
    port map (
            O => \N__14367\,
            I => \N__14361\
        );

    \I__2625\ : CascadeMux
    port map (
            O => \N__14364\,
            I => \N__14358\
        );

    \I__2624\ : CascadeBuf
    port map (
            O => \N__14361\,
            I => \N__14355\
        );

    \I__2623\ : CascadeBuf
    port map (
            O => \N__14358\,
            I => \N__14352\
        );

    \I__2622\ : CascadeMux
    port map (
            O => \N__14355\,
            I => \N__14349\
        );

    \I__2621\ : CascadeMux
    port map (
            O => \N__14352\,
            I => \N__14346\
        );

    \I__2620\ : CascadeBuf
    port map (
            O => \N__14349\,
            I => \N__14343\
        );

    \I__2619\ : CascadeBuf
    port map (
            O => \N__14346\,
            I => \N__14340\
        );

    \I__2618\ : CascadeMux
    port map (
            O => \N__14343\,
            I => \N__14337\
        );

    \I__2617\ : CascadeMux
    port map (
            O => \N__14340\,
            I => \N__14334\
        );

    \I__2616\ : CascadeBuf
    port map (
            O => \N__14337\,
            I => \N__14331\
        );

    \I__2615\ : CascadeBuf
    port map (
            O => \N__14334\,
            I => \N__14328\
        );

    \I__2614\ : CascadeMux
    port map (
            O => \N__14331\,
            I => \N__14325\
        );

    \I__2613\ : CascadeMux
    port map (
            O => \N__14328\,
            I => \N__14322\
        );

    \I__2612\ : CascadeBuf
    port map (
            O => \N__14325\,
            I => \N__14319\
        );

    \I__2611\ : CascadeBuf
    port map (
            O => \N__14322\,
            I => \N__14316\
        );

    \I__2610\ : CascadeMux
    port map (
            O => \N__14319\,
            I => \N__14313\
        );

    \I__2609\ : CascadeMux
    port map (
            O => \N__14316\,
            I => \N__14310\
        );

    \I__2608\ : CascadeBuf
    port map (
            O => \N__14313\,
            I => \N__14307\
        );

    \I__2607\ : CascadeBuf
    port map (
            O => \N__14310\,
            I => \N__14304\
        );

    \I__2606\ : CascadeMux
    port map (
            O => \N__14307\,
            I => \N__14301\
        );

    \I__2605\ : CascadeMux
    port map (
            O => \N__14304\,
            I => \N__14298\
        );

    \I__2604\ : CascadeBuf
    port map (
            O => \N__14301\,
            I => \N__14295\
        );

    \I__2603\ : CascadeBuf
    port map (
            O => \N__14298\,
            I => \N__14292\
        );

    \I__2602\ : CascadeMux
    port map (
            O => \N__14295\,
            I => \N__14289\
        );

    \I__2601\ : CascadeMux
    port map (
            O => \N__14292\,
            I => \N__14286\
        );

    \I__2600\ : CascadeBuf
    port map (
            O => \N__14289\,
            I => \N__14283\
        );

    \I__2599\ : CascadeBuf
    port map (
            O => \N__14286\,
            I => \N__14280\
        );

    \I__2598\ : CascadeMux
    port map (
            O => \N__14283\,
            I => \N__14277\
        );

    \I__2597\ : CascadeMux
    port map (
            O => \N__14280\,
            I => \N__14274\
        );

    \I__2596\ : CascadeBuf
    port map (
            O => \N__14277\,
            I => \N__14271\
        );

    \I__2595\ : CascadeBuf
    port map (
            O => \N__14274\,
            I => \N__14268\
        );

    \I__2594\ : CascadeMux
    port map (
            O => \N__14271\,
            I => \N__14265\
        );

    \I__2593\ : CascadeMux
    port map (
            O => \N__14268\,
            I => \N__14262\
        );

    \I__2592\ : CascadeBuf
    port map (
            O => \N__14265\,
            I => \N__14259\
        );

    \I__2591\ : CascadeBuf
    port map (
            O => \N__14262\,
            I => \N__14256\
        );

    \I__2590\ : CascadeMux
    port map (
            O => \N__14259\,
            I => \N__14253\
        );

    \I__2589\ : CascadeMux
    port map (
            O => \N__14256\,
            I => \N__14250\
        );

    \I__2588\ : CascadeBuf
    port map (
            O => \N__14253\,
            I => \N__14247\
        );

    \I__2587\ : CascadeBuf
    port map (
            O => \N__14250\,
            I => \N__14244\
        );

    \I__2586\ : CascadeMux
    port map (
            O => \N__14247\,
            I => \N__14241\
        );

    \I__2585\ : CascadeMux
    port map (
            O => \N__14244\,
            I => \N__14238\
        );

    \I__2584\ : CascadeBuf
    port map (
            O => \N__14241\,
            I => \N__14235\
        );

    \I__2583\ : CascadeBuf
    port map (
            O => \N__14238\,
            I => \N__14232\
        );

    \I__2582\ : CascadeMux
    port map (
            O => \N__14235\,
            I => \N__14229\
        );

    \I__2581\ : CascadeMux
    port map (
            O => \N__14232\,
            I => \N__14226\
        );

    \I__2580\ : CascadeBuf
    port map (
            O => \N__14229\,
            I => \N__14223\
        );

    \I__2579\ : CascadeBuf
    port map (
            O => \N__14226\,
            I => \N__14220\
        );

    \I__2578\ : CascadeMux
    port map (
            O => \N__14223\,
            I => \N__14217\
        );

    \I__2577\ : CascadeMux
    port map (
            O => \N__14220\,
            I => \N__14214\
        );

    \I__2576\ : CascadeBuf
    port map (
            O => \N__14217\,
            I => \N__14211\
        );

    \I__2575\ : InMux
    port map (
            O => \N__14214\,
            I => \N__14207\
        );

    \I__2574\ : CascadeMux
    port map (
            O => \N__14211\,
            I => \N__14204\
        );

    \I__2573\ : InMux
    port map (
            O => \N__14210\,
            I => \N__14201\
        );

    \I__2572\ : LocalMux
    port map (
            O => \N__14207\,
            I => \N__14198\
        );

    \I__2571\ : InMux
    port map (
            O => \N__14204\,
            I => \N__14195\
        );

    \I__2570\ : LocalMux
    port map (
            O => \N__14201\,
            I => \N__14192\
        );

    \I__2569\ : Span4Mux_s1_v
    port map (
            O => \N__14198\,
            I => \N__14189\
        );

    \I__2568\ : LocalMux
    port map (
            O => \N__14195\,
            I => \N__14186\
        );

    \I__2567\ : Span12Mux_h
    port map (
            O => \N__14192\,
            I => \N__14183\
        );

    \I__2566\ : Span4Mux_h
    port map (
            O => \N__14189\,
            I => \N__14179\
        );

    \I__2565\ : Span4Mux_s1_v
    port map (
            O => \N__14186\,
            I => \N__14176\
        );

    \I__2564\ : Span12Mux_v
    port map (
            O => \N__14183\,
            I => \N__14173\
        );

    \I__2563\ : InMux
    port map (
            O => \N__14182\,
            I => \N__14170\
        );

    \I__2562\ : Span4Mux_h
    port map (
            O => \N__14179\,
            I => \N__14165\
        );

    \I__2561\ : Span4Mux_h
    port map (
            O => \N__14176\,
            I => \N__14165\
        );

    \I__2560\ : Odrv12
    port map (
            O => \N__14173\,
            I => \RX_ADDR_8\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__14170\,
            I => \RX_ADDR_8\
        );

    \I__2558\ : Odrv4
    port map (
            O => \N__14165\,
            I => \RX_ADDR_8\
        );

    \I__2557\ : InMux
    port map (
            O => \N__14158\,
            I => \N__14155\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__14155\,
            I => \N__14152\
        );

    \I__2555\ : Span12Mux_s7_v
    port map (
            O => \N__14152\,
            I => \N__14149\
        );

    \I__2554\ : Span12Mux_v
    port map (
            O => \N__14149\,
            I => \N__14146\
        );

    \I__2553\ : Odrv12
    port map (
            O => \N__14146\,
            I => \receive_module.n127\
        );

    \I__2552\ : CascadeMux
    port map (
            O => \N__14143\,
            I => \N__14140\
        );

    \I__2551\ : CascadeBuf
    port map (
            O => \N__14140\,
            I => \N__14136\
        );

    \I__2550\ : CascadeMux
    port map (
            O => \N__14139\,
            I => \N__14133\
        );

    \I__2549\ : CascadeMux
    port map (
            O => \N__14136\,
            I => \N__14130\
        );

    \I__2548\ : CascadeBuf
    port map (
            O => \N__14133\,
            I => \N__14127\
        );

    \I__2547\ : CascadeBuf
    port map (
            O => \N__14130\,
            I => \N__14124\
        );

    \I__2546\ : CascadeMux
    port map (
            O => \N__14127\,
            I => \N__14121\
        );

    \I__2545\ : CascadeMux
    port map (
            O => \N__14124\,
            I => \N__14118\
        );

    \I__2544\ : CascadeBuf
    port map (
            O => \N__14121\,
            I => \N__14115\
        );

    \I__2543\ : CascadeBuf
    port map (
            O => \N__14118\,
            I => \N__14112\
        );

    \I__2542\ : CascadeMux
    port map (
            O => \N__14115\,
            I => \N__14109\
        );

    \I__2541\ : CascadeMux
    port map (
            O => \N__14112\,
            I => \N__14106\
        );

    \I__2540\ : CascadeBuf
    port map (
            O => \N__14109\,
            I => \N__14103\
        );

    \I__2539\ : CascadeBuf
    port map (
            O => \N__14106\,
            I => \N__14100\
        );

    \I__2538\ : CascadeMux
    port map (
            O => \N__14103\,
            I => \N__14097\
        );

    \I__2537\ : CascadeMux
    port map (
            O => \N__14100\,
            I => \N__14094\
        );

    \I__2536\ : CascadeBuf
    port map (
            O => \N__14097\,
            I => \N__14091\
        );

    \I__2535\ : CascadeBuf
    port map (
            O => \N__14094\,
            I => \N__14088\
        );

    \I__2534\ : CascadeMux
    port map (
            O => \N__14091\,
            I => \N__14085\
        );

    \I__2533\ : CascadeMux
    port map (
            O => \N__14088\,
            I => \N__14082\
        );

    \I__2532\ : CascadeBuf
    port map (
            O => \N__14085\,
            I => \N__14079\
        );

    \I__2531\ : CascadeBuf
    port map (
            O => \N__14082\,
            I => \N__14076\
        );

    \I__2530\ : CascadeMux
    port map (
            O => \N__14079\,
            I => \N__14073\
        );

    \I__2529\ : CascadeMux
    port map (
            O => \N__14076\,
            I => \N__14070\
        );

    \I__2528\ : CascadeBuf
    port map (
            O => \N__14073\,
            I => \N__14067\
        );

    \I__2527\ : CascadeBuf
    port map (
            O => \N__14070\,
            I => \N__14064\
        );

    \I__2526\ : CascadeMux
    port map (
            O => \N__14067\,
            I => \N__14061\
        );

    \I__2525\ : CascadeMux
    port map (
            O => \N__14064\,
            I => \N__14058\
        );

    \I__2524\ : CascadeBuf
    port map (
            O => \N__14061\,
            I => \N__14055\
        );

    \I__2523\ : CascadeBuf
    port map (
            O => \N__14058\,
            I => \N__14052\
        );

    \I__2522\ : CascadeMux
    port map (
            O => \N__14055\,
            I => \N__14049\
        );

    \I__2521\ : CascadeMux
    port map (
            O => \N__14052\,
            I => \N__14046\
        );

    \I__2520\ : CascadeBuf
    port map (
            O => \N__14049\,
            I => \N__14043\
        );

    \I__2519\ : CascadeBuf
    port map (
            O => \N__14046\,
            I => \N__14040\
        );

    \I__2518\ : CascadeMux
    port map (
            O => \N__14043\,
            I => \N__14037\
        );

    \I__2517\ : CascadeMux
    port map (
            O => \N__14040\,
            I => \N__14034\
        );

    \I__2516\ : CascadeBuf
    port map (
            O => \N__14037\,
            I => \N__14031\
        );

    \I__2515\ : CascadeBuf
    port map (
            O => \N__14034\,
            I => \N__14028\
        );

    \I__2514\ : CascadeMux
    port map (
            O => \N__14031\,
            I => \N__14025\
        );

    \I__2513\ : CascadeMux
    port map (
            O => \N__14028\,
            I => \N__14022\
        );

    \I__2512\ : CascadeBuf
    port map (
            O => \N__14025\,
            I => \N__14019\
        );

    \I__2511\ : CascadeBuf
    port map (
            O => \N__14022\,
            I => \N__14016\
        );

    \I__2510\ : CascadeMux
    port map (
            O => \N__14019\,
            I => \N__14013\
        );

    \I__2509\ : CascadeMux
    port map (
            O => \N__14016\,
            I => \N__14010\
        );

    \I__2508\ : CascadeBuf
    port map (
            O => \N__14013\,
            I => \N__14007\
        );

    \I__2507\ : CascadeBuf
    port map (
            O => \N__14010\,
            I => \N__14004\
        );

    \I__2506\ : CascadeMux
    port map (
            O => \N__14007\,
            I => \N__14001\
        );

    \I__2505\ : CascadeMux
    port map (
            O => \N__14004\,
            I => \N__13998\
        );

    \I__2504\ : CascadeBuf
    port map (
            O => \N__14001\,
            I => \N__13995\
        );

    \I__2503\ : CascadeBuf
    port map (
            O => \N__13998\,
            I => \N__13992\
        );

    \I__2502\ : CascadeMux
    port map (
            O => \N__13995\,
            I => \N__13989\
        );

    \I__2501\ : CascadeMux
    port map (
            O => \N__13992\,
            I => \N__13986\
        );

    \I__2500\ : CascadeBuf
    port map (
            O => \N__13989\,
            I => \N__13983\
        );

    \I__2499\ : CascadeBuf
    port map (
            O => \N__13986\,
            I => \N__13980\
        );

    \I__2498\ : CascadeMux
    port map (
            O => \N__13983\,
            I => \N__13977\
        );

    \I__2497\ : CascadeMux
    port map (
            O => \N__13980\,
            I => \N__13973\
        );

    \I__2496\ : CascadeBuf
    port map (
            O => \N__13977\,
            I => \N__13970\
        );

    \I__2495\ : InMux
    port map (
            O => \N__13976\,
            I => \N__13967\
        );

    \I__2494\ : CascadeBuf
    port map (
            O => \N__13973\,
            I => \N__13964\
        );

    \I__2493\ : CascadeMux
    port map (
            O => \N__13970\,
            I => \N__13961\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__13967\,
            I => \N__13958\
        );

    \I__2491\ : CascadeMux
    port map (
            O => \N__13964\,
            I => \N__13955\
        );

    \I__2490\ : CascadeBuf
    port map (
            O => \N__13961\,
            I => \N__13952\
        );

    \I__2489\ : Span4Mux_v
    port map (
            O => \N__13958\,
            I => \N__13949\
        );

    \I__2488\ : InMux
    port map (
            O => \N__13955\,
            I => \N__13946\
        );

    \I__2487\ : CascadeMux
    port map (
            O => \N__13952\,
            I => \N__13943\
        );

    \I__2486\ : Span4Mux_v
    port map (
            O => \N__13949\,
            I => \N__13939\
        );

    \I__2485\ : LocalMux
    port map (
            O => \N__13946\,
            I => \N__13936\
        );

    \I__2484\ : InMux
    port map (
            O => \N__13943\,
            I => \N__13933\
        );

    \I__2483\ : CascadeMux
    port map (
            O => \N__13942\,
            I => \N__13930\
        );

    \I__2482\ : Span4Mux_v
    port map (
            O => \N__13939\,
            I => \N__13927\
        );

    \I__2481\ : Span4Mux_s1_v
    port map (
            O => \N__13936\,
            I => \N__13924\
        );

    \I__2480\ : LocalMux
    port map (
            O => \N__13933\,
            I => \N__13921\
        );

    \I__2479\ : InMux
    port map (
            O => \N__13930\,
            I => \N__13918\
        );

    \I__2478\ : Sp12to4
    port map (
            O => \N__13927\,
            I => \N__13915\
        );

    \I__2477\ : Span4Mux_h
    port map (
            O => \N__13924\,
            I => \N__13912\
        );

    \I__2476\ : Span12Mux_s1_v
    port map (
            O => \N__13921\,
            I => \N__13909\
        );

    \I__2475\ : LocalMux
    port map (
            O => \N__13918\,
            I => \RX_ADDR_9\
        );

    \I__2474\ : Odrv12
    port map (
            O => \N__13915\,
            I => \RX_ADDR_9\
        );

    \I__2473\ : Odrv4
    port map (
            O => \N__13912\,
            I => \RX_ADDR_9\
        );

    \I__2472\ : Odrv12
    port map (
            O => \N__13909\,
            I => \RX_ADDR_9\
        );

    \I__2471\ : InMux
    port map (
            O => \N__13900\,
            I => \N__13897\
        );

    \I__2470\ : LocalMux
    port map (
            O => \N__13897\,
            I => \transmit_module.ADDR_Y_COMPONENT_9\
        );

    \I__2469\ : InMux
    port map (
            O => \N__13894\,
            I => \N__13891\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__13891\,
            I => \N__13888\
        );

    \I__2467\ : Odrv4
    port map (
            O => \N__13888\,
            I => \transmit_module.ADDR_Y_COMPONENT_12\
        );

    \I__2466\ : InMux
    port map (
            O => \N__13885\,
            I => \N__13882\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__13882\,
            I => \N__13879\
        );

    \I__2464\ : Odrv4
    port map (
            O => \N__13879\,
            I => \transmit_module.n120\
        );

    \I__2463\ : InMux
    port map (
            O => \N__13876\,
            I => \N__13873\
        );

    \I__2462\ : LocalMux
    port map (
            O => \N__13873\,
            I => \N__13870\
        );

    \I__2461\ : Odrv4
    port map (
            O => \N__13870\,
            I => \transmit_module.n119\
        );

    \I__2460\ : InMux
    port map (
            O => \N__13867\,
            I => \N__13864\
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__13864\,
            I => \N__13861\
        );

    \I__2458\ : Span4Mux_h
    port map (
            O => \N__13861\,
            I => \N__13858\
        );

    \I__2457\ : Odrv4
    port map (
            O => \N__13858\,
            I => \transmit_module.ADDR_Y_COMPONENT_11\
        );

    \I__2456\ : InMux
    port map (
            O => \N__13855\,
            I => \N__13852\
        );

    \I__2455\ : LocalMux
    port map (
            O => \N__13852\,
            I => \N__13849\
        );

    \I__2454\ : Odrv4
    port map (
            O => \N__13849\,
            I => \transmit_module.n121\
        );

    \I__2453\ : CEMux
    port map (
            O => \N__13846\,
            I => \N__13843\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__13843\,
            I => \N__13839\
        );

    \I__2451\ : CEMux
    port map (
            O => \N__13842\,
            I => \N__13836\
        );

    \I__2450\ : Span4Mux_v
    port map (
            O => \N__13839\,
            I => \N__13833\
        );

    \I__2449\ : LocalMux
    port map (
            O => \N__13836\,
            I => \N__13830\
        );

    \I__2448\ : Span4Mux_h
    port map (
            O => \N__13833\,
            I => \N__13827\
        );

    \I__2447\ : Odrv4
    port map (
            O => \N__13830\,
            I => \transmit_module.n2039\
        );

    \I__2446\ : Odrv4
    port map (
            O => \N__13827\,
            I => \transmit_module.n2039\
        );

    \I__2445\ : InMux
    port map (
            O => \N__13822\,
            I => \N__13819\
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__13819\,
            I => \N__13816\
        );

    \I__2443\ : Odrv12
    port map (
            O => \N__13816\,
            I => \transmit_module.n130\
        );

    \I__2442\ : InMux
    port map (
            O => \N__13813\,
            I => \N__13810\
        );

    \I__2441\ : LocalMux
    port map (
            O => \N__13810\,
            I => \line_buffer.n3755\
        );

    \I__2440\ : InMux
    port map (
            O => \N__13807\,
            I => \N__13804\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__13804\,
            I => \N__13801\
        );

    \I__2438\ : Span4Mux_v
    port map (
            O => \N__13801\,
            I => \N__13798\
        );

    \I__2437\ : Odrv4
    port map (
            O => \N__13798\,
            I => \TX_DATA_0\
        );

    \I__2436\ : InMux
    port map (
            O => \N__13795\,
            I => \N__13792\
        );

    \I__2435\ : LocalMux
    port map (
            O => \N__13792\,
            I => \N__13789\
        );

    \I__2434\ : Span12Mux_v
    port map (
            O => \N__13789\,
            I => \N__13786\
        );

    \I__2433\ : Odrv12
    port map (
            O => \N__13786\,
            I => \receive_module.n134\
        );

    \I__2432\ : CascadeMux
    port map (
            O => \N__13783\,
            I => \N__13779\
        );

    \I__2431\ : CascadeMux
    port map (
            O => \N__13782\,
            I => \N__13776\
        );

    \I__2430\ : CascadeBuf
    port map (
            O => \N__13779\,
            I => \N__13773\
        );

    \I__2429\ : CascadeBuf
    port map (
            O => \N__13776\,
            I => \N__13770\
        );

    \I__2428\ : CascadeMux
    port map (
            O => \N__13773\,
            I => \N__13767\
        );

    \I__2427\ : CascadeMux
    port map (
            O => \N__13770\,
            I => \N__13764\
        );

    \I__2426\ : CascadeBuf
    port map (
            O => \N__13767\,
            I => \N__13761\
        );

    \I__2425\ : CascadeBuf
    port map (
            O => \N__13764\,
            I => \N__13758\
        );

    \I__2424\ : CascadeMux
    port map (
            O => \N__13761\,
            I => \N__13755\
        );

    \I__2423\ : CascadeMux
    port map (
            O => \N__13758\,
            I => \N__13752\
        );

    \I__2422\ : CascadeBuf
    port map (
            O => \N__13755\,
            I => \N__13749\
        );

    \I__2421\ : CascadeBuf
    port map (
            O => \N__13752\,
            I => \N__13746\
        );

    \I__2420\ : CascadeMux
    port map (
            O => \N__13749\,
            I => \N__13743\
        );

    \I__2419\ : CascadeMux
    port map (
            O => \N__13746\,
            I => \N__13740\
        );

    \I__2418\ : CascadeBuf
    port map (
            O => \N__13743\,
            I => \N__13737\
        );

    \I__2417\ : CascadeBuf
    port map (
            O => \N__13740\,
            I => \N__13734\
        );

    \I__2416\ : CascadeMux
    port map (
            O => \N__13737\,
            I => \N__13731\
        );

    \I__2415\ : CascadeMux
    port map (
            O => \N__13734\,
            I => \N__13728\
        );

    \I__2414\ : CascadeBuf
    port map (
            O => \N__13731\,
            I => \N__13725\
        );

    \I__2413\ : CascadeBuf
    port map (
            O => \N__13728\,
            I => \N__13722\
        );

    \I__2412\ : CascadeMux
    port map (
            O => \N__13725\,
            I => \N__13719\
        );

    \I__2411\ : CascadeMux
    port map (
            O => \N__13722\,
            I => \N__13716\
        );

    \I__2410\ : CascadeBuf
    port map (
            O => \N__13719\,
            I => \N__13713\
        );

    \I__2409\ : CascadeBuf
    port map (
            O => \N__13716\,
            I => \N__13710\
        );

    \I__2408\ : CascadeMux
    port map (
            O => \N__13713\,
            I => \N__13707\
        );

    \I__2407\ : CascadeMux
    port map (
            O => \N__13710\,
            I => \N__13704\
        );

    \I__2406\ : CascadeBuf
    port map (
            O => \N__13707\,
            I => \N__13701\
        );

    \I__2405\ : CascadeBuf
    port map (
            O => \N__13704\,
            I => \N__13698\
        );

    \I__2404\ : CascadeMux
    port map (
            O => \N__13701\,
            I => \N__13695\
        );

    \I__2403\ : CascadeMux
    port map (
            O => \N__13698\,
            I => \N__13692\
        );

    \I__2402\ : CascadeBuf
    port map (
            O => \N__13695\,
            I => \N__13689\
        );

    \I__2401\ : CascadeBuf
    port map (
            O => \N__13692\,
            I => \N__13686\
        );

    \I__2400\ : CascadeMux
    port map (
            O => \N__13689\,
            I => \N__13683\
        );

    \I__2399\ : CascadeMux
    port map (
            O => \N__13686\,
            I => \N__13680\
        );

    \I__2398\ : CascadeBuf
    port map (
            O => \N__13683\,
            I => \N__13677\
        );

    \I__2397\ : CascadeBuf
    port map (
            O => \N__13680\,
            I => \N__13674\
        );

    \I__2396\ : CascadeMux
    port map (
            O => \N__13677\,
            I => \N__13671\
        );

    \I__2395\ : CascadeMux
    port map (
            O => \N__13674\,
            I => \N__13668\
        );

    \I__2394\ : CascadeBuf
    port map (
            O => \N__13671\,
            I => \N__13665\
        );

    \I__2393\ : CascadeBuf
    port map (
            O => \N__13668\,
            I => \N__13662\
        );

    \I__2392\ : CascadeMux
    port map (
            O => \N__13665\,
            I => \N__13659\
        );

    \I__2391\ : CascadeMux
    port map (
            O => \N__13662\,
            I => \N__13656\
        );

    \I__2390\ : CascadeBuf
    port map (
            O => \N__13659\,
            I => \N__13653\
        );

    \I__2389\ : CascadeBuf
    port map (
            O => \N__13656\,
            I => \N__13650\
        );

    \I__2388\ : CascadeMux
    port map (
            O => \N__13653\,
            I => \N__13647\
        );

    \I__2387\ : CascadeMux
    port map (
            O => \N__13650\,
            I => \N__13644\
        );

    \I__2386\ : CascadeBuf
    port map (
            O => \N__13647\,
            I => \N__13641\
        );

    \I__2385\ : CascadeBuf
    port map (
            O => \N__13644\,
            I => \N__13638\
        );

    \I__2384\ : CascadeMux
    port map (
            O => \N__13641\,
            I => \N__13635\
        );

    \I__2383\ : CascadeMux
    port map (
            O => \N__13638\,
            I => \N__13632\
        );

    \I__2382\ : CascadeBuf
    port map (
            O => \N__13635\,
            I => \N__13629\
        );

    \I__2381\ : CascadeBuf
    port map (
            O => \N__13632\,
            I => \N__13626\
        );

    \I__2380\ : CascadeMux
    port map (
            O => \N__13629\,
            I => \N__13623\
        );

    \I__2379\ : CascadeMux
    port map (
            O => \N__13626\,
            I => \N__13620\
        );

    \I__2378\ : CascadeBuf
    port map (
            O => \N__13623\,
            I => \N__13617\
        );

    \I__2377\ : CascadeBuf
    port map (
            O => \N__13620\,
            I => \N__13614\
        );

    \I__2376\ : CascadeMux
    port map (
            O => \N__13617\,
            I => \N__13611\
        );

    \I__2375\ : CascadeMux
    port map (
            O => \N__13614\,
            I => \N__13608\
        );

    \I__2374\ : CascadeBuf
    port map (
            O => \N__13611\,
            I => \N__13605\
        );

    \I__2373\ : CascadeBuf
    port map (
            O => \N__13608\,
            I => \N__13602\
        );

    \I__2372\ : CascadeMux
    port map (
            O => \N__13605\,
            I => \N__13599\
        );

    \I__2371\ : CascadeMux
    port map (
            O => \N__13602\,
            I => \N__13596\
        );

    \I__2370\ : InMux
    port map (
            O => \N__13599\,
            I => \N__13593\
        );

    \I__2369\ : InMux
    port map (
            O => \N__13596\,
            I => \N__13590\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__13593\,
            I => \N__13586\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__13590\,
            I => \N__13583\
        );

    \I__2366\ : InMux
    port map (
            O => \N__13589\,
            I => \N__13580\
        );

    \I__2365\ : Span4Mux_h
    port map (
            O => \N__13586\,
            I => \N__13577\
        );

    \I__2364\ : Span4Mux_h
    port map (
            O => \N__13583\,
            I => \N__13574\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__13580\,
            I => \N__13571\
        );

    \I__2362\ : Sp12to4
    port map (
            O => \N__13577\,
            I => \N__13567\
        );

    \I__2361\ : Sp12to4
    port map (
            O => \N__13574\,
            I => \N__13564\
        );

    \I__2360\ : Span12Mux_v
    port map (
            O => \N__13571\,
            I => \N__13561\
        );

    \I__2359\ : InMux
    port map (
            O => \N__13570\,
            I => \N__13558\
        );

    \I__2358\ : Span12Mux_v
    port map (
            O => \N__13567\,
            I => \N__13553\
        );

    \I__2357\ : Span12Mux_v
    port map (
            O => \N__13564\,
            I => \N__13553\
        );

    \I__2356\ : Odrv12
    port map (
            O => \N__13561\,
            I => \RX_ADDR_2\
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__13558\,
            I => \RX_ADDR_2\
        );

    \I__2354\ : Odrv12
    port map (
            O => \N__13553\,
            I => \RX_ADDR_2\
        );

    \I__2353\ : CascadeMux
    port map (
            O => \N__13546\,
            I => \N__13540\
        );

    \I__2352\ : InMux
    port map (
            O => \N__13545\,
            I => \N__13537\
        );

    \I__2351\ : CascadeMux
    port map (
            O => \N__13544\,
            I => \N__13534\
        );

    \I__2350\ : InMux
    port map (
            O => \N__13543\,
            I => \N__13531\
        );

    \I__2349\ : InMux
    port map (
            O => \N__13540\,
            I => \N__13528\
        );

    \I__2348\ : LocalMux
    port map (
            O => \N__13537\,
            I => \N__13525\
        );

    \I__2347\ : InMux
    port map (
            O => \N__13534\,
            I => \N__13522\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__13531\,
            I => \transmit_module.TX_ADDR_7\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__13528\,
            I => \transmit_module.TX_ADDR_7\
        );

    \I__2344\ : Odrv4
    port map (
            O => \N__13525\,
            I => \transmit_module.TX_ADDR_7\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__13522\,
            I => \transmit_module.TX_ADDR_7\
        );

    \I__2342\ : InMux
    port map (
            O => \N__13513\,
            I => \N__13510\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__13510\,
            I => \transmit_module.n125\
        );

    \I__2340\ : InMux
    port map (
            O => \N__13507\,
            I => \transmit_module.n3264\
        );

    \I__2339\ : InMux
    port map (
            O => \N__13504\,
            I => \bfn_15_14_0_\
        );

    \I__2338\ : InMux
    port map (
            O => \N__13501\,
            I => \transmit_module.n3266\
        );

    \I__2337\ : InMux
    port map (
            O => \N__13498\,
            I => \N__13492\
        );

    \I__2336\ : InMux
    port map (
            O => \N__13497\,
            I => \N__13487\
        );

    \I__2335\ : InMux
    port map (
            O => \N__13496\,
            I => \N__13487\
        );

    \I__2334\ : InMux
    port map (
            O => \N__13495\,
            I => \N__13484\
        );

    \I__2333\ : LocalMux
    port map (
            O => \N__13492\,
            I => \transmit_module.TX_ADDR_10\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__13487\,
            I => \transmit_module.TX_ADDR_10\
        );

    \I__2331\ : LocalMux
    port map (
            O => \N__13484\,
            I => \transmit_module.TX_ADDR_10\
        );

    \I__2330\ : InMux
    port map (
            O => \N__13477\,
            I => \N__13474\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__13474\,
            I => \transmit_module.n122\
        );

    \I__2328\ : InMux
    port map (
            O => \N__13471\,
            I => \transmit_module.n3267\
        );

    \I__2327\ : InMux
    port map (
            O => \N__13468\,
            I => \transmit_module.n3268\
        );

    \I__2326\ : InMux
    port map (
            O => \N__13465\,
            I => \transmit_module.n3269\
        );

    \I__2325\ : InMux
    port map (
            O => \N__13462\,
            I => \transmit_module.n3270\
        );

    \I__2324\ : InMux
    port map (
            O => \N__13459\,
            I => \receive_module.n3257\
        );

    \I__2323\ : InMux
    port map (
            O => \N__13456\,
            I => \N__13451\
        );

    \I__2322\ : InMux
    port map (
            O => \N__13455\,
            I => \N__13448\
        );

    \I__2321\ : InMux
    port map (
            O => \N__13454\,
            I => \N__13445\
        );

    \I__2320\ : LocalMux
    port map (
            O => \N__13451\,
            I => \N__13440\
        );

    \I__2319\ : LocalMux
    port map (
            O => \N__13448\,
            I => \N__13440\
        );

    \I__2318\ : LocalMux
    port map (
            O => \N__13445\,
            I => \N__13434\
        );

    \I__2317\ : Span4Mux_v
    port map (
            O => \N__13440\,
            I => \N__13434\
        );

    \I__2316\ : InMux
    port map (
            O => \N__13439\,
            I => \N__13431\
        );

    \I__2315\ : Odrv4
    port map (
            O => \N__13434\,
            I => \transmit_module.TX_ADDR_0\
        );

    \I__2314\ : LocalMux
    port map (
            O => \N__13431\,
            I => \transmit_module.TX_ADDR_0\
        );

    \I__2313\ : InMux
    port map (
            O => \N__13426\,
            I => \N__13423\
        );

    \I__2312\ : LocalMux
    port map (
            O => \N__13423\,
            I => \N__13419\
        );

    \I__2311\ : CascadeMux
    port map (
            O => \N__13422\,
            I => \N__13416\
        );

    \I__2310\ : Span4Mux_v
    port map (
            O => \N__13419\,
            I => \N__13413\
        );

    \I__2309\ : InMux
    port map (
            O => \N__13416\,
            I => \N__13410\
        );

    \I__2308\ : Span4Mux_h
    port map (
            O => \N__13413\,
            I => \N__13407\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__13410\,
            I => \N__13404\
        );

    \I__2306\ : Odrv4
    port map (
            O => \N__13407\,
            I => \transmit_module.X_DELTA_PATTERN_0\
        );

    \I__2305\ : Odrv4
    port map (
            O => \N__13404\,
            I => \transmit_module.X_DELTA_PATTERN_0\
        );

    \I__2304\ : InMux
    port map (
            O => \N__13399\,
            I => \N__13396\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__13396\,
            I => \N__13393\
        );

    \I__2302\ : Odrv4
    port map (
            O => \N__13393\,
            I => \transmit_module.n132\
        );

    \I__2301\ : InMux
    port map (
            O => \N__13390\,
            I => \N__13386\
        );

    \I__2300\ : CascadeMux
    port map (
            O => \N__13389\,
            I => \N__13381\
        );

    \I__2299\ : LocalMux
    port map (
            O => \N__13386\,
            I => \N__13378\
        );

    \I__2298\ : InMux
    port map (
            O => \N__13385\,
            I => \N__13373\
        );

    \I__2297\ : InMux
    port map (
            O => \N__13384\,
            I => \N__13373\
        );

    \I__2296\ : InMux
    port map (
            O => \N__13381\,
            I => \N__13370\
        );

    \I__2295\ : Odrv4
    port map (
            O => \N__13378\,
            I => \transmit_module.TX_ADDR_1\
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__13373\,
            I => \transmit_module.TX_ADDR_1\
        );

    \I__2293\ : LocalMux
    port map (
            O => \N__13370\,
            I => \transmit_module.TX_ADDR_1\
        );

    \I__2292\ : CascadeMux
    port map (
            O => \N__13363\,
            I => \N__13360\
        );

    \I__2291\ : InMux
    port map (
            O => \N__13360\,
            I => \N__13357\
        );

    \I__2290\ : LocalMux
    port map (
            O => \N__13357\,
            I => \N__13354\
        );

    \I__2289\ : Odrv4
    port map (
            O => \N__13354\,
            I => \transmit_module.n131\
        );

    \I__2288\ : InMux
    port map (
            O => \N__13351\,
            I => \transmit_module.n3258\
        );

    \I__2287\ : InMux
    port map (
            O => \N__13348\,
            I => \transmit_module.n3259\
        );

    \I__2286\ : InMux
    port map (
            O => \N__13345\,
            I => \transmit_module.n3260\
        );

    \I__2285\ : InMux
    port map (
            O => \N__13342\,
            I => \N__13339\
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__13339\,
            I => \N__13333\
        );

    \I__2283\ : InMux
    port map (
            O => \N__13338\,
            I => \N__13330\
        );

    \I__2282\ : InMux
    port map (
            O => \N__13337\,
            I => \N__13327\
        );

    \I__2281\ : InMux
    port map (
            O => \N__13336\,
            I => \N__13324\
        );

    \I__2280\ : Odrv4
    port map (
            O => \N__13333\,
            I => \transmit_module.TX_ADDR_4\
        );

    \I__2279\ : LocalMux
    port map (
            O => \N__13330\,
            I => \transmit_module.TX_ADDR_4\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__13327\,
            I => \transmit_module.TX_ADDR_4\
        );

    \I__2277\ : LocalMux
    port map (
            O => \N__13324\,
            I => \transmit_module.TX_ADDR_4\
        );

    \I__2276\ : InMux
    port map (
            O => \N__13315\,
            I => \N__13312\
        );

    \I__2275\ : LocalMux
    port map (
            O => \N__13312\,
            I => \transmit_module.n128\
        );

    \I__2274\ : InMux
    port map (
            O => \N__13309\,
            I => \transmit_module.n3261\
        );

    \I__2273\ : InMux
    port map (
            O => \N__13306\,
            I => \N__13301\
        );

    \I__2272\ : InMux
    port map (
            O => \N__13305\,
            I => \N__13298\
        );

    \I__2271\ : CascadeMux
    port map (
            O => \N__13304\,
            I => \N__13294\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__13301\,
            I => \N__13289\
        );

    \I__2269\ : LocalMux
    port map (
            O => \N__13298\,
            I => \N__13289\
        );

    \I__2268\ : InMux
    port map (
            O => \N__13297\,
            I => \N__13286\
        );

    \I__2267\ : InMux
    port map (
            O => \N__13294\,
            I => \N__13283\
        );

    \I__2266\ : Odrv4
    port map (
            O => \N__13289\,
            I => \transmit_module.TX_ADDR_5\
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__13286\,
            I => \transmit_module.TX_ADDR_5\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__13283\,
            I => \transmit_module.TX_ADDR_5\
        );

    \I__2263\ : InMux
    port map (
            O => \N__13276\,
            I => \N__13273\
        );

    \I__2262\ : LocalMux
    port map (
            O => \N__13273\,
            I => \transmit_module.n127\
        );

    \I__2261\ : InMux
    port map (
            O => \N__13270\,
            I => \transmit_module.n3262\
        );

    \I__2260\ : InMux
    port map (
            O => \N__13267\,
            I => \N__13262\
        );

    \I__2259\ : InMux
    port map (
            O => \N__13266\,
            I => \N__13259\
        );

    \I__2258\ : CascadeMux
    port map (
            O => \N__13265\,
            I => \N__13255\
        );

    \I__2257\ : LocalMux
    port map (
            O => \N__13262\,
            I => \N__13252\
        );

    \I__2256\ : LocalMux
    port map (
            O => \N__13259\,
            I => \N__13249\
        );

    \I__2255\ : InMux
    port map (
            O => \N__13258\,
            I => \N__13246\
        );

    \I__2254\ : InMux
    port map (
            O => \N__13255\,
            I => \N__13243\
        );

    \I__2253\ : Odrv12
    port map (
            O => \N__13252\,
            I => \transmit_module.TX_ADDR_6\
        );

    \I__2252\ : Odrv4
    port map (
            O => \N__13249\,
            I => \transmit_module.TX_ADDR_6\
        );

    \I__2251\ : LocalMux
    port map (
            O => \N__13246\,
            I => \transmit_module.TX_ADDR_6\
        );

    \I__2250\ : LocalMux
    port map (
            O => \N__13243\,
            I => \transmit_module.TX_ADDR_6\
        );

    \I__2249\ : InMux
    port map (
            O => \N__13234\,
            I => \N__13231\
        );

    \I__2248\ : LocalMux
    port map (
            O => \N__13231\,
            I => \transmit_module.n126\
        );

    \I__2247\ : InMux
    port map (
            O => \N__13228\,
            I => \transmit_module.n3263\
        );

    \I__2246\ : InMux
    port map (
            O => \N__13225\,
            I => \receive_module.n3248\
        );

    \I__2245\ : InMux
    port map (
            O => \N__13222\,
            I => \receive_module.n3249\
        );

    \I__2244\ : InMux
    port map (
            O => \N__13219\,
            I => \receive_module.n3250\
        );

    \I__2243\ : InMux
    port map (
            O => \N__13216\,
            I => \receive_module.n3251\
        );

    \I__2242\ : InMux
    port map (
            O => \N__13213\,
            I => \bfn_15_12_0_\
        );

    \I__2241\ : InMux
    port map (
            O => \N__13210\,
            I => \receive_module.n3253\
        );

    \I__2240\ : InMux
    port map (
            O => \N__13207\,
            I => \receive_module.n3254\
        );

    \I__2239\ : InMux
    port map (
            O => \N__13204\,
            I => \receive_module.n3255\
        );

    \I__2238\ : InMux
    port map (
            O => \N__13201\,
            I => \receive_module.n3256\
        );

    \I__2237\ : InMux
    port map (
            O => \N__13198\,
            I => \N__13195\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__13195\,
            I => \N__13192\
        );

    \I__2235\ : Span4Mux_h
    port map (
            O => \N__13192\,
            I => \N__13189\
        );

    \I__2234\ : Span4Mux_h
    port map (
            O => \N__13189\,
            I => \N__13186\
        );

    \I__2233\ : Odrv4
    port map (
            O => \N__13186\,
            I => \line_buffer.n543\
        );

    \I__2232\ : InMux
    port map (
            O => \N__13183\,
            I => \N__13180\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__13180\,
            I => \N__13177\
        );

    \I__2230\ : Span4Mux_h
    port map (
            O => \N__13177\,
            I => \N__13174\
        );

    \I__2229\ : Span4Mux_h
    port map (
            O => \N__13174\,
            I => \N__13171\
        );

    \I__2228\ : Span4Mux_h
    port map (
            O => \N__13171\,
            I => \N__13168\
        );

    \I__2227\ : Odrv4
    port map (
            O => \N__13168\,
            I => \line_buffer.n535\
        );

    \I__2226\ : InMux
    port map (
            O => \N__13165\,
            I => \N__13161\
        );

    \I__2225\ : InMux
    port map (
            O => \N__13164\,
            I => \N__13156\
        );

    \I__2224\ : LocalMux
    port map (
            O => \N__13161\,
            I => \N__13153\
        );

    \I__2223\ : InMux
    port map (
            O => \N__13160\,
            I => \N__13148\
        );

    \I__2222\ : InMux
    port map (
            O => \N__13159\,
            I => \N__13148\
        );

    \I__2221\ : LocalMux
    port map (
            O => \N__13156\,
            I => \receive_module.rx_counter.Y_7\
        );

    \I__2220\ : Odrv4
    port map (
            O => \N__13153\,
            I => \receive_module.rx_counter.Y_7\
        );

    \I__2219\ : LocalMux
    port map (
            O => \N__13148\,
            I => \receive_module.rx_counter.Y_7\
        );

    \I__2218\ : InMux
    port map (
            O => \N__13141\,
            I => \N__13137\
        );

    \I__2217\ : InMux
    port map (
            O => \N__13140\,
            I => \N__13134\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__13137\,
            I => \receive_module.rx_counter.n3791\
        );

    \I__2215\ : LocalMux
    port map (
            O => \N__13134\,
            I => \receive_module.rx_counter.n3791\
        );

    \I__2214\ : CascadeMux
    port map (
            O => \N__13129\,
            I => \N__13126\
        );

    \I__2213\ : InMux
    port map (
            O => \N__13126\,
            I => \N__13123\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__13123\,
            I => \N__13117\
        );

    \I__2211\ : InMux
    port map (
            O => \N__13122\,
            I => \N__13114\
        );

    \I__2210\ : InMux
    port map (
            O => \N__13121\,
            I => \N__13109\
        );

    \I__2209\ : InMux
    port map (
            O => \N__13120\,
            I => \N__13109\
        );

    \I__2208\ : Odrv4
    port map (
            O => \N__13117\,
            I => \receive_module.rx_counter.Y_4\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__13114\,
            I => \receive_module.rx_counter.Y_4\
        );

    \I__2206\ : LocalMux
    port map (
            O => \N__13109\,
            I => \receive_module.rx_counter.Y_4\
        );

    \I__2205\ : InMux
    port map (
            O => \N__13102\,
            I => \N__13099\
        );

    \I__2204\ : LocalMux
    port map (
            O => \N__13099\,
            I => \receive_module.rx_counter.n3551\
        );

    \I__2203\ : CEMux
    port map (
            O => \N__13096\,
            I => \N__13093\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__13093\,
            I => \N__13089\
        );

    \I__2201\ : CEMux
    port map (
            O => \N__13092\,
            I => \N__13086\
        );

    \I__2200\ : Span4Mux_h
    port map (
            O => \N__13089\,
            I => \N__13083\
        );

    \I__2199\ : LocalMux
    port map (
            O => \N__13086\,
            I => \N__13080\
        );

    \I__2198\ : Odrv4
    port map (
            O => \N__13083\,
            I => \receive_module.rx_counter.n2045\
        );

    \I__2197\ : Odrv12
    port map (
            O => \N__13080\,
            I => \receive_module.rx_counter.n2045\
        );

    \I__2196\ : InMux
    port map (
            O => \N__13075\,
            I => \N__13072\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__13072\,
            I => \receive_module.rx_counter.old_HS\
        );

    \I__2194\ : InMux
    port map (
            O => \N__13069\,
            I => \bfn_15_11_0_\
        );

    \I__2193\ : InMux
    port map (
            O => \N__13066\,
            I => \receive_module.n3245\
        );

    \I__2192\ : InMux
    port map (
            O => \N__13063\,
            I => \receive_module.n3246\
        );

    \I__2191\ : InMux
    port map (
            O => \N__13060\,
            I => \receive_module.n3247\
        );

    \I__2190\ : InMux
    port map (
            O => \N__13057\,
            I => \N__13054\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__13054\,
            I => \N__13050\
        );

    \I__2188\ : InMux
    port map (
            O => \N__13053\,
            I => \N__13047\
        );

    \I__2187\ : Span4Mux_v
    port map (
            O => \N__13050\,
            I => \N__13044\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__13047\,
            I => \N__13041\
        );

    \I__2185\ : Span4Mux_v
    port map (
            O => \N__13044\,
            I => \N__13038\
        );

    \I__2184\ : Odrv4
    port map (
            O => \N__13041\,
            I => \transmit_module.n110\
        );

    \I__2183\ : Odrv4
    port map (
            O => \N__13038\,
            I => \transmit_module.n110\
        );

    \I__2182\ : InMux
    port map (
            O => \N__13033\,
            I => \N__13030\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__13030\,
            I => \N__13027\
        );

    \I__2180\ : Span12Mux_v
    port map (
            O => \N__13027\,
            I => \N__13024\
        );

    \I__2179\ : Odrv12
    port map (
            O => \N__13024\,
            I => \transmit_module.n141\
        );

    \I__2178\ : CascadeMux
    port map (
            O => \N__13021\,
            I => \N__13018\
        );

    \I__2177\ : CascadeBuf
    port map (
            O => \N__13018\,
            I => \N__13015\
        );

    \I__2176\ : CascadeMux
    port map (
            O => \N__13015\,
            I => \N__13011\
        );

    \I__2175\ : CascadeMux
    port map (
            O => \N__13014\,
            I => \N__13008\
        );

    \I__2174\ : CascadeBuf
    port map (
            O => \N__13011\,
            I => \N__13005\
        );

    \I__2173\ : CascadeBuf
    port map (
            O => \N__13008\,
            I => \N__13002\
        );

    \I__2172\ : CascadeMux
    port map (
            O => \N__13005\,
            I => \N__12999\
        );

    \I__2171\ : CascadeMux
    port map (
            O => \N__13002\,
            I => \N__12996\
        );

    \I__2170\ : CascadeBuf
    port map (
            O => \N__12999\,
            I => \N__12993\
        );

    \I__2169\ : CascadeBuf
    port map (
            O => \N__12996\,
            I => \N__12990\
        );

    \I__2168\ : CascadeMux
    port map (
            O => \N__12993\,
            I => \N__12987\
        );

    \I__2167\ : CascadeMux
    port map (
            O => \N__12990\,
            I => \N__12984\
        );

    \I__2166\ : CascadeBuf
    port map (
            O => \N__12987\,
            I => \N__12981\
        );

    \I__2165\ : CascadeBuf
    port map (
            O => \N__12984\,
            I => \N__12978\
        );

    \I__2164\ : CascadeMux
    port map (
            O => \N__12981\,
            I => \N__12975\
        );

    \I__2163\ : CascadeMux
    port map (
            O => \N__12978\,
            I => \N__12972\
        );

    \I__2162\ : CascadeBuf
    port map (
            O => \N__12975\,
            I => \N__12969\
        );

    \I__2161\ : CascadeBuf
    port map (
            O => \N__12972\,
            I => \N__12966\
        );

    \I__2160\ : CascadeMux
    port map (
            O => \N__12969\,
            I => \N__12963\
        );

    \I__2159\ : CascadeMux
    port map (
            O => \N__12966\,
            I => \N__12960\
        );

    \I__2158\ : CascadeBuf
    port map (
            O => \N__12963\,
            I => \N__12957\
        );

    \I__2157\ : CascadeBuf
    port map (
            O => \N__12960\,
            I => \N__12954\
        );

    \I__2156\ : CascadeMux
    port map (
            O => \N__12957\,
            I => \N__12951\
        );

    \I__2155\ : CascadeMux
    port map (
            O => \N__12954\,
            I => \N__12948\
        );

    \I__2154\ : CascadeBuf
    port map (
            O => \N__12951\,
            I => \N__12945\
        );

    \I__2153\ : CascadeBuf
    port map (
            O => \N__12948\,
            I => \N__12942\
        );

    \I__2152\ : CascadeMux
    port map (
            O => \N__12945\,
            I => \N__12939\
        );

    \I__2151\ : CascadeMux
    port map (
            O => \N__12942\,
            I => \N__12936\
        );

    \I__2150\ : CascadeBuf
    port map (
            O => \N__12939\,
            I => \N__12933\
        );

    \I__2149\ : CascadeBuf
    port map (
            O => \N__12936\,
            I => \N__12930\
        );

    \I__2148\ : CascadeMux
    port map (
            O => \N__12933\,
            I => \N__12927\
        );

    \I__2147\ : CascadeMux
    port map (
            O => \N__12930\,
            I => \N__12924\
        );

    \I__2146\ : CascadeBuf
    port map (
            O => \N__12927\,
            I => \N__12921\
        );

    \I__2145\ : CascadeBuf
    port map (
            O => \N__12924\,
            I => \N__12918\
        );

    \I__2144\ : CascadeMux
    port map (
            O => \N__12921\,
            I => \N__12915\
        );

    \I__2143\ : CascadeMux
    port map (
            O => \N__12918\,
            I => \N__12912\
        );

    \I__2142\ : CascadeBuf
    port map (
            O => \N__12915\,
            I => \N__12909\
        );

    \I__2141\ : CascadeBuf
    port map (
            O => \N__12912\,
            I => \N__12906\
        );

    \I__2140\ : CascadeMux
    port map (
            O => \N__12909\,
            I => \N__12903\
        );

    \I__2139\ : CascadeMux
    port map (
            O => \N__12906\,
            I => \N__12900\
        );

    \I__2138\ : CascadeBuf
    port map (
            O => \N__12903\,
            I => \N__12897\
        );

    \I__2137\ : CascadeBuf
    port map (
            O => \N__12900\,
            I => \N__12894\
        );

    \I__2136\ : CascadeMux
    port map (
            O => \N__12897\,
            I => \N__12891\
        );

    \I__2135\ : CascadeMux
    port map (
            O => \N__12894\,
            I => \N__12888\
        );

    \I__2134\ : CascadeBuf
    port map (
            O => \N__12891\,
            I => \N__12885\
        );

    \I__2133\ : CascadeBuf
    port map (
            O => \N__12888\,
            I => \N__12882\
        );

    \I__2132\ : CascadeMux
    port map (
            O => \N__12885\,
            I => \N__12879\
        );

    \I__2131\ : CascadeMux
    port map (
            O => \N__12882\,
            I => \N__12876\
        );

    \I__2130\ : CascadeBuf
    port map (
            O => \N__12879\,
            I => \N__12873\
        );

    \I__2129\ : CascadeBuf
    port map (
            O => \N__12876\,
            I => \N__12870\
        );

    \I__2128\ : CascadeMux
    port map (
            O => \N__12873\,
            I => \N__12867\
        );

    \I__2127\ : CascadeMux
    port map (
            O => \N__12870\,
            I => \N__12864\
        );

    \I__2126\ : CascadeBuf
    port map (
            O => \N__12867\,
            I => \N__12861\
        );

    \I__2125\ : CascadeBuf
    port map (
            O => \N__12864\,
            I => \N__12858\
        );

    \I__2124\ : CascadeMux
    port map (
            O => \N__12861\,
            I => \N__12855\
        );

    \I__2123\ : CascadeMux
    port map (
            O => \N__12858\,
            I => \N__12852\
        );

    \I__2122\ : CascadeBuf
    port map (
            O => \N__12855\,
            I => \N__12849\
        );

    \I__2121\ : CascadeBuf
    port map (
            O => \N__12852\,
            I => \N__12846\
        );

    \I__2120\ : CascadeMux
    port map (
            O => \N__12849\,
            I => \N__12843\
        );

    \I__2119\ : CascadeMux
    port map (
            O => \N__12846\,
            I => \N__12840\
        );

    \I__2118\ : InMux
    port map (
            O => \N__12843\,
            I => \N__12837\
        );

    \I__2117\ : CascadeBuf
    port map (
            O => \N__12840\,
            I => \N__12834\
        );

    \I__2116\ : LocalMux
    port map (
            O => \N__12837\,
            I => \N__12831\
        );

    \I__2115\ : CascadeMux
    port map (
            O => \N__12834\,
            I => \N__12828\
        );

    \I__2114\ : Span4Mux_h
    port map (
            O => \N__12831\,
            I => \N__12825\
        );

    \I__2113\ : InMux
    port map (
            O => \N__12828\,
            I => \N__12822\
        );

    \I__2112\ : Span4Mux_h
    port map (
            O => \N__12825\,
            I => \N__12819\
        );

    \I__2111\ : LocalMux
    port map (
            O => \N__12822\,
            I => \N__12816\
        );

    \I__2110\ : Span4Mux_h
    port map (
            O => \N__12819\,
            I => \N__12813\
        );

    \I__2109\ : Span12Mux_s4_v
    port map (
            O => \N__12816\,
            I => \N__12810\
        );

    \I__2108\ : Odrv4
    port map (
            O => \N__12813\,
            I => n22
        );

    \I__2107\ : Odrv12
    port map (
            O => \N__12810\,
            I => n22
        );

    \I__2106\ : InMux
    port map (
            O => \N__12805\,
            I => \N__12802\
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__12802\,
            I => \N__12798\
        );

    \I__2104\ : InMux
    port map (
            O => \N__12801\,
            I => \N__12795\
        );

    \I__2103\ : Span12Mux_s4_v
    port map (
            O => \N__12798\,
            I => \N__12792\
        );

    \I__2102\ : LocalMux
    port map (
            O => \N__12795\,
            I => \N__12789\
        );

    \I__2101\ : Span12Mux_v
    port map (
            O => \N__12792\,
            I => \N__12786\
        );

    \I__2100\ : Odrv4
    port map (
            O => \N__12789\,
            I => \transmit_module.n109\
        );

    \I__2099\ : Odrv12
    port map (
            O => \N__12786\,
            I => \transmit_module.n109\
        );

    \I__2098\ : InMux
    port map (
            O => \N__12781\,
            I => \N__12778\
        );

    \I__2097\ : LocalMux
    port map (
            O => \N__12778\,
            I => \N__12774\
        );

    \I__2096\ : InMux
    port map (
            O => \N__12777\,
            I => \N__12771\
        );

    \I__2095\ : Span12Mux_s11_v
    port map (
            O => \N__12774\,
            I => \N__12768\
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__12771\,
            I => \transmit_module.n140\
        );

    \I__2093\ : Odrv12
    port map (
            O => \N__12768\,
            I => \transmit_module.n140\
        );

    \I__2092\ : CascadeMux
    port map (
            O => \N__12763\,
            I => \N__12759\
        );

    \I__2091\ : CascadeMux
    port map (
            O => \N__12762\,
            I => \N__12756\
        );

    \I__2090\ : CascadeBuf
    port map (
            O => \N__12759\,
            I => \N__12753\
        );

    \I__2089\ : CascadeBuf
    port map (
            O => \N__12756\,
            I => \N__12750\
        );

    \I__2088\ : CascadeMux
    port map (
            O => \N__12753\,
            I => \N__12747\
        );

    \I__2087\ : CascadeMux
    port map (
            O => \N__12750\,
            I => \N__12744\
        );

    \I__2086\ : CascadeBuf
    port map (
            O => \N__12747\,
            I => \N__12741\
        );

    \I__2085\ : CascadeBuf
    port map (
            O => \N__12744\,
            I => \N__12738\
        );

    \I__2084\ : CascadeMux
    port map (
            O => \N__12741\,
            I => \N__12735\
        );

    \I__2083\ : CascadeMux
    port map (
            O => \N__12738\,
            I => \N__12732\
        );

    \I__2082\ : CascadeBuf
    port map (
            O => \N__12735\,
            I => \N__12729\
        );

    \I__2081\ : CascadeBuf
    port map (
            O => \N__12732\,
            I => \N__12726\
        );

    \I__2080\ : CascadeMux
    port map (
            O => \N__12729\,
            I => \N__12723\
        );

    \I__2079\ : CascadeMux
    port map (
            O => \N__12726\,
            I => \N__12720\
        );

    \I__2078\ : CascadeBuf
    port map (
            O => \N__12723\,
            I => \N__12717\
        );

    \I__2077\ : CascadeBuf
    port map (
            O => \N__12720\,
            I => \N__12714\
        );

    \I__2076\ : CascadeMux
    port map (
            O => \N__12717\,
            I => \N__12711\
        );

    \I__2075\ : CascadeMux
    port map (
            O => \N__12714\,
            I => \N__12708\
        );

    \I__2074\ : CascadeBuf
    port map (
            O => \N__12711\,
            I => \N__12705\
        );

    \I__2073\ : CascadeBuf
    port map (
            O => \N__12708\,
            I => \N__12702\
        );

    \I__2072\ : CascadeMux
    port map (
            O => \N__12705\,
            I => \N__12699\
        );

    \I__2071\ : CascadeMux
    port map (
            O => \N__12702\,
            I => \N__12696\
        );

    \I__2070\ : CascadeBuf
    port map (
            O => \N__12699\,
            I => \N__12693\
        );

    \I__2069\ : CascadeBuf
    port map (
            O => \N__12696\,
            I => \N__12690\
        );

    \I__2068\ : CascadeMux
    port map (
            O => \N__12693\,
            I => \N__12687\
        );

    \I__2067\ : CascadeMux
    port map (
            O => \N__12690\,
            I => \N__12684\
        );

    \I__2066\ : CascadeBuf
    port map (
            O => \N__12687\,
            I => \N__12681\
        );

    \I__2065\ : CascadeBuf
    port map (
            O => \N__12684\,
            I => \N__12678\
        );

    \I__2064\ : CascadeMux
    port map (
            O => \N__12681\,
            I => \N__12675\
        );

    \I__2063\ : CascadeMux
    port map (
            O => \N__12678\,
            I => \N__12672\
        );

    \I__2062\ : CascadeBuf
    port map (
            O => \N__12675\,
            I => \N__12669\
        );

    \I__2061\ : CascadeBuf
    port map (
            O => \N__12672\,
            I => \N__12666\
        );

    \I__2060\ : CascadeMux
    port map (
            O => \N__12669\,
            I => \N__12663\
        );

    \I__2059\ : CascadeMux
    port map (
            O => \N__12666\,
            I => \N__12660\
        );

    \I__2058\ : CascadeBuf
    port map (
            O => \N__12663\,
            I => \N__12657\
        );

    \I__2057\ : CascadeBuf
    port map (
            O => \N__12660\,
            I => \N__12654\
        );

    \I__2056\ : CascadeMux
    port map (
            O => \N__12657\,
            I => \N__12651\
        );

    \I__2055\ : CascadeMux
    port map (
            O => \N__12654\,
            I => \N__12648\
        );

    \I__2054\ : CascadeBuf
    port map (
            O => \N__12651\,
            I => \N__12645\
        );

    \I__2053\ : CascadeBuf
    port map (
            O => \N__12648\,
            I => \N__12642\
        );

    \I__2052\ : CascadeMux
    port map (
            O => \N__12645\,
            I => \N__12639\
        );

    \I__2051\ : CascadeMux
    port map (
            O => \N__12642\,
            I => \N__12636\
        );

    \I__2050\ : CascadeBuf
    port map (
            O => \N__12639\,
            I => \N__12633\
        );

    \I__2049\ : CascadeBuf
    port map (
            O => \N__12636\,
            I => \N__12630\
        );

    \I__2048\ : CascadeMux
    port map (
            O => \N__12633\,
            I => \N__12627\
        );

    \I__2047\ : CascadeMux
    port map (
            O => \N__12630\,
            I => \N__12624\
        );

    \I__2046\ : CascadeBuf
    port map (
            O => \N__12627\,
            I => \N__12621\
        );

    \I__2045\ : CascadeBuf
    port map (
            O => \N__12624\,
            I => \N__12618\
        );

    \I__2044\ : CascadeMux
    port map (
            O => \N__12621\,
            I => \N__12615\
        );

    \I__2043\ : CascadeMux
    port map (
            O => \N__12618\,
            I => \N__12612\
        );

    \I__2042\ : CascadeBuf
    port map (
            O => \N__12615\,
            I => \N__12609\
        );

    \I__2041\ : CascadeBuf
    port map (
            O => \N__12612\,
            I => \N__12606\
        );

    \I__2040\ : CascadeMux
    port map (
            O => \N__12609\,
            I => \N__12603\
        );

    \I__2039\ : CascadeMux
    port map (
            O => \N__12606\,
            I => \N__12600\
        );

    \I__2038\ : CascadeBuf
    port map (
            O => \N__12603\,
            I => \N__12597\
        );

    \I__2037\ : CascadeBuf
    port map (
            O => \N__12600\,
            I => \N__12594\
        );

    \I__2036\ : CascadeMux
    port map (
            O => \N__12597\,
            I => \N__12591\
        );

    \I__2035\ : CascadeMux
    port map (
            O => \N__12594\,
            I => \N__12588\
        );

    \I__2034\ : CascadeBuf
    port map (
            O => \N__12591\,
            I => \N__12585\
        );

    \I__2033\ : CascadeBuf
    port map (
            O => \N__12588\,
            I => \N__12582\
        );

    \I__2032\ : CascadeMux
    port map (
            O => \N__12585\,
            I => \N__12579\
        );

    \I__2031\ : CascadeMux
    port map (
            O => \N__12582\,
            I => \N__12576\
        );

    \I__2030\ : InMux
    port map (
            O => \N__12579\,
            I => \N__12573\
        );

    \I__2029\ : InMux
    port map (
            O => \N__12576\,
            I => \N__12570\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__12573\,
            I => \N__12567\
        );

    \I__2027\ : LocalMux
    port map (
            O => \N__12570\,
            I => \N__12564\
        );

    \I__2026\ : Span12Mux_s9_h
    port map (
            O => \N__12567\,
            I => \N__12561\
        );

    \I__2025\ : Span4Mux_h
    port map (
            O => \N__12564\,
            I => \N__12558\
        );

    \I__2024\ : Odrv12
    port map (
            O => \N__12561\,
            I => n21
        );

    \I__2023\ : Odrv4
    port map (
            O => \N__12558\,
            I => n21
        );

    \I__2022\ : IoInMux
    port map (
            O => \N__12553\,
            I => \N__12550\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__12550\,
            I => \N__12547\
        );

    \I__2020\ : Span4Mux_s3_v
    port map (
            O => \N__12547\,
            I => \N__12544\
        );

    \I__2019\ : Span4Mux_h
    port map (
            O => \N__12544\,
            I => \N__12540\
        );

    \I__2018\ : InMux
    port map (
            O => \N__12543\,
            I => \N__12537\
        );

    \I__2017\ : Odrv4
    port map (
            O => \N__12540\,
            I => \LED_c\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__12537\,
            I => \LED_c\
        );

    \I__2015\ : CascadeMux
    port map (
            O => \N__12532\,
            I => \receive_module.rx_counter.n3628_cascade_\
        );

    \I__2014\ : InMux
    port map (
            O => \N__12529\,
            I => \N__12526\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__12526\,
            I => \receive_module.rx_counter.n7_adj_609\
        );

    \I__2012\ : InMux
    port map (
            O => \N__12523\,
            I => \N__12520\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__12520\,
            I => \receive_module.rx_counter.n11\
        );

    \I__2010\ : CascadeMux
    port map (
            O => \N__12517\,
            I => \receive_module.rx_counter.n11_cascade_\
        );

    \I__2009\ : InMux
    port map (
            O => \N__12514\,
            I => \N__12508\
        );

    \I__2008\ : InMux
    port map (
            O => \N__12513\,
            I => \N__12508\
        );

    \I__2007\ : LocalMux
    port map (
            O => \N__12508\,
            I => \receive_module.rx_counter.old_VS\
        );

    \I__2006\ : InMux
    port map (
            O => \N__12505\,
            I => \N__12502\
        );

    \I__2005\ : LocalMux
    port map (
            O => \N__12502\,
            I => \N__12499\
        );

    \I__2004\ : Odrv4
    port map (
            O => \N__12499\,
            I => \transmit_module.ADDR_Y_COMPONENT_6\
        );

    \I__2003\ : InMux
    port map (
            O => \N__12496\,
            I => \N__12492\
        );

    \I__2002\ : InMux
    port map (
            O => \N__12495\,
            I => \N__12489\
        );

    \I__2001\ : LocalMux
    port map (
            O => \N__12492\,
            I => \N__12486\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__12489\,
            I => \transmit_module.n106\
        );

    \I__1999\ : Odrv12
    port map (
            O => \N__12486\,
            I => \transmit_module.n106\
        );

    \I__1998\ : InMux
    port map (
            O => \N__12481\,
            I => \N__12478\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__12478\,
            I => \N__12475\
        );

    \I__1996\ : Odrv12
    port map (
            O => \N__12475\,
            I => \transmit_module.n137\
        );

    \I__1995\ : CascadeMux
    port map (
            O => \N__12472\,
            I => \N__12469\
        );

    \I__1994\ : CascadeBuf
    port map (
            O => \N__12469\,
            I => \N__12465\
        );

    \I__1993\ : CascadeMux
    port map (
            O => \N__12468\,
            I => \N__12462\
        );

    \I__1992\ : CascadeMux
    port map (
            O => \N__12465\,
            I => \N__12459\
        );

    \I__1991\ : CascadeBuf
    port map (
            O => \N__12462\,
            I => \N__12456\
        );

    \I__1990\ : CascadeBuf
    port map (
            O => \N__12459\,
            I => \N__12453\
        );

    \I__1989\ : CascadeMux
    port map (
            O => \N__12456\,
            I => \N__12450\
        );

    \I__1988\ : CascadeMux
    port map (
            O => \N__12453\,
            I => \N__12447\
        );

    \I__1987\ : CascadeBuf
    port map (
            O => \N__12450\,
            I => \N__12444\
        );

    \I__1986\ : CascadeBuf
    port map (
            O => \N__12447\,
            I => \N__12441\
        );

    \I__1985\ : CascadeMux
    port map (
            O => \N__12444\,
            I => \N__12438\
        );

    \I__1984\ : CascadeMux
    port map (
            O => \N__12441\,
            I => \N__12435\
        );

    \I__1983\ : CascadeBuf
    port map (
            O => \N__12438\,
            I => \N__12432\
        );

    \I__1982\ : CascadeBuf
    port map (
            O => \N__12435\,
            I => \N__12429\
        );

    \I__1981\ : CascadeMux
    port map (
            O => \N__12432\,
            I => \N__12426\
        );

    \I__1980\ : CascadeMux
    port map (
            O => \N__12429\,
            I => \N__12423\
        );

    \I__1979\ : CascadeBuf
    port map (
            O => \N__12426\,
            I => \N__12420\
        );

    \I__1978\ : CascadeBuf
    port map (
            O => \N__12423\,
            I => \N__12417\
        );

    \I__1977\ : CascadeMux
    port map (
            O => \N__12420\,
            I => \N__12414\
        );

    \I__1976\ : CascadeMux
    port map (
            O => \N__12417\,
            I => \N__12411\
        );

    \I__1975\ : CascadeBuf
    port map (
            O => \N__12414\,
            I => \N__12408\
        );

    \I__1974\ : CascadeBuf
    port map (
            O => \N__12411\,
            I => \N__12405\
        );

    \I__1973\ : CascadeMux
    port map (
            O => \N__12408\,
            I => \N__12402\
        );

    \I__1972\ : CascadeMux
    port map (
            O => \N__12405\,
            I => \N__12399\
        );

    \I__1971\ : CascadeBuf
    port map (
            O => \N__12402\,
            I => \N__12396\
        );

    \I__1970\ : CascadeBuf
    port map (
            O => \N__12399\,
            I => \N__12393\
        );

    \I__1969\ : CascadeMux
    port map (
            O => \N__12396\,
            I => \N__12390\
        );

    \I__1968\ : CascadeMux
    port map (
            O => \N__12393\,
            I => \N__12387\
        );

    \I__1967\ : CascadeBuf
    port map (
            O => \N__12390\,
            I => \N__12384\
        );

    \I__1966\ : CascadeBuf
    port map (
            O => \N__12387\,
            I => \N__12381\
        );

    \I__1965\ : CascadeMux
    port map (
            O => \N__12384\,
            I => \N__12378\
        );

    \I__1964\ : CascadeMux
    port map (
            O => \N__12381\,
            I => \N__12375\
        );

    \I__1963\ : CascadeBuf
    port map (
            O => \N__12378\,
            I => \N__12372\
        );

    \I__1962\ : CascadeBuf
    port map (
            O => \N__12375\,
            I => \N__12369\
        );

    \I__1961\ : CascadeMux
    port map (
            O => \N__12372\,
            I => \N__12366\
        );

    \I__1960\ : CascadeMux
    port map (
            O => \N__12369\,
            I => \N__12363\
        );

    \I__1959\ : CascadeBuf
    port map (
            O => \N__12366\,
            I => \N__12360\
        );

    \I__1958\ : CascadeBuf
    port map (
            O => \N__12363\,
            I => \N__12357\
        );

    \I__1957\ : CascadeMux
    port map (
            O => \N__12360\,
            I => \N__12354\
        );

    \I__1956\ : CascadeMux
    port map (
            O => \N__12357\,
            I => \N__12351\
        );

    \I__1955\ : CascadeBuf
    port map (
            O => \N__12354\,
            I => \N__12348\
        );

    \I__1954\ : CascadeBuf
    port map (
            O => \N__12351\,
            I => \N__12345\
        );

    \I__1953\ : CascadeMux
    port map (
            O => \N__12348\,
            I => \N__12342\
        );

    \I__1952\ : CascadeMux
    port map (
            O => \N__12345\,
            I => \N__12339\
        );

    \I__1951\ : CascadeBuf
    port map (
            O => \N__12342\,
            I => \N__12336\
        );

    \I__1950\ : CascadeBuf
    port map (
            O => \N__12339\,
            I => \N__12333\
        );

    \I__1949\ : CascadeMux
    port map (
            O => \N__12336\,
            I => \N__12330\
        );

    \I__1948\ : CascadeMux
    port map (
            O => \N__12333\,
            I => \N__12327\
        );

    \I__1947\ : CascadeBuf
    port map (
            O => \N__12330\,
            I => \N__12324\
        );

    \I__1946\ : CascadeBuf
    port map (
            O => \N__12327\,
            I => \N__12321\
        );

    \I__1945\ : CascadeMux
    port map (
            O => \N__12324\,
            I => \N__12318\
        );

    \I__1944\ : CascadeMux
    port map (
            O => \N__12321\,
            I => \N__12315\
        );

    \I__1943\ : CascadeBuf
    port map (
            O => \N__12318\,
            I => \N__12312\
        );

    \I__1942\ : CascadeBuf
    port map (
            O => \N__12315\,
            I => \N__12309\
        );

    \I__1941\ : CascadeMux
    port map (
            O => \N__12312\,
            I => \N__12306\
        );

    \I__1940\ : CascadeMux
    port map (
            O => \N__12309\,
            I => \N__12303\
        );

    \I__1939\ : CascadeBuf
    port map (
            O => \N__12306\,
            I => \N__12300\
        );

    \I__1938\ : CascadeBuf
    port map (
            O => \N__12303\,
            I => \N__12297\
        );

    \I__1937\ : CascadeMux
    port map (
            O => \N__12300\,
            I => \N__12294\
        );

    \I__1936\ : CascadeMux
    port map (
            O => \N__12297\,
            I => \N__12291\
        );

    \I__1935\ : CascadeBuf
    port map (
            O => \N__12294\,
            I => \N__12288\
        );

    \I__1934\ : InMux
    port map (
            O => \N__12291\,
            I => \N__12285\
        );

    \I__1933\ : CascadeMux
    port map (
            O => \N__12288\,
            I => \N__12282\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__12285\,
            I => \N__12279\
        );

    \I__1931\ : InMux
    port map (
            O => \N__12282\,
            I => \N__12276\
        );

    \I__1930\ : Span4Mux_v
    port map (
            O => \N__12279\,
            I => \N__12273\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__12276\,
            I => \N__12270\
        );

    \I__1928\ : Span4Mux_v
    port map (
            O => \N__12273\,
            I => \N__12267\
        );

    \I__1927\ : Span4Mux_v
    port map (
            O => \N__12270\,
            I => \N__12264\
        );

    \I__1926\ : Span4Mux_v
    port map (
            O => \N__12267\,
            I => \N__12261\
        );

    \I__1925\ : Span4Mux_v
    port map (
            O => \N__12264\,
            I => \N__12258\
        );

    \I__1924\ : Span4Mux_h
    port map (
            O => \N__12261\,
            I => \N__12255\
        );

    \I__1923\ : Span4Mux_v
    port map (
            O => \N__12258\,
            I => \N__12252\
        );

    \I__1922\ : Span4Mux_h
    port map (
            O => \N__12255\,
            I => \N__12247\
        );

    \I__1921\ : Span4Mux_h
    port map (
            O => \N__12252\,
            I => \N__12247\
        );

    \I__1920\ : Odrv4
    port map (
            O => \N__12247\,
            I => n18
        );

    \I__1919\ : InMux
    port map (
            O => \N__12244\,
            I => \N__12241\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__12241\,
            I => \transmit_module.ADDR_Y_COMPONENT_0\
        );

    \I__1917\ : InMux
    port map (
            O => \N__12238\,
            I => \N__12235\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__12235\,
            I => \line_buffer.n3722\
        );

    \I__1915\ : InMux
    port map (
            O => \N__12232\,
            I => \N__12229\
        );

    \I__1914\ : LocalMux
    port map (
            O => \N__12229\,
            I => \N__12226\
        );

    \I__1913\ : Odrv4
    port map (
            O => \N__12226\,
            I => \TX_DATA_6\
        );

    \I__1912\ : IoInMux
    port map (
            O => \N__12223\,
            I => \N__12220\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__12220\,
            I => \N__12216\
        );

    \I__1910\ : IoInMux
    port map (
            O => \N__12219\,
            I => \N__12212\
        );

    \I__1909\ : Span4Mux_s2_v
    port map (
            O => \N__12216\,
            I => \N__12209\
        );

    \I__1908\ : IoInMux
    port map (
            O => \N__12215\,
            I => \N__12206\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__12212\,
            I => \N__12203\
        );

    \I__1906\ : Span4Mux_h
    port map (
            O => \N__12209\,
            I => \N__12200\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__12206\,
            I => \N__12197\
        );

    \I__1904\ : Span4Mux_s2_v
    port map (
            O => \N__12203\,
            I => \N__12194\
        );

    \I__1903\ : Sp12to4
    port map (
            O => \N__12200\,
            I => \N__12191\
        );

    \I__1902\ : Span12Mux_s1_h
    port map (
            O => \N__12197\,
            I => \N__12188\
        );

    \I__1901\ : Span4Mux_h
    port map (
            O => \N__12194\,
            I => \N__12185\
        );

    \I__1900\ : Span12Mux_h
    port map (
            O => \N__12191\,
            I => \N__12180\
        );

    \I__1899\ : Span12Mux_h
    port map (
            O => \N__12188\,
            I => \N__12180\
        );

    \I__1898\ : Span4Mux_v
    port map (
            O => \N__12185\,
            I => \N__12177\
        );

    \I__1897\ : Odrv12
    port map (
            O => \N__12180\,
            I => n1792
        );

    \I__1896\ : Odrv4
    port map (
            O => \N__12177\,
            I => n1792
        );

    \I__1895\ : IoInMux
    port map (
            O => \N__12172\,
            I => \N__12169\
        );

    \I__1894\ : LocalMux
    port map (
            O => \N__12169\,
            I => \N__12164\
        );

    \I__1893\ : IoInMux
    port map (
            O => \N__12168\,
            I => \N__12161\
        );

    \I__1892\ : IoInMux
    port map (
            O => \N__12167\,
            I => \N__12158\
        );

    \I__1891\ : Span4Mux_s1_h
    port map (
            O => \N__12164\,
            I => \N__12155\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__12161\,
            I => \N__12152\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__12158\,
            I => \N__12149\
        );

    \I__1888\ : Span4Mux_h
    port map (
            O => \N__12155\,
            I => \N__12146\
        );

    \I__1887\ : IoSpan4Mux
    port map (
            O => \N__12152\,
            I => \N__12143\
        );

    \I__1886\ : Span12Mux_s8_v
    port map (
            O => \N__12149\,
            I => \N__12140\
        );

    \I__1885\ : Span4Mux_h
    port map (
            O => \N__12146\,
            I => \N__12137\
        );

    \I__1884\ : Span4Mux_s1_v
    port map (
            O => \N__12143\,
            I => \N__12134\
        );

    \I__1883\ : Span12Mux_h
    port map (
            O => \N__12140\,
            I => \N__12131\
        );

    \I__1882\ : Span4Mux_h
    port map (
            O => \N__12137\,
            I => \N__12126\
        );

    \I__1881\ : Span4Mux_v
    port map (
            O => \N__12134\,
            I => \N__12126\
        );

    \I__1880\ : Odrv12
    port map (
            O => \N__12131\,
            I => n1798
        );

    \I__1879\ : Odrv4
    port map (
            O => \N__12126\,
            I => n1798
        );

    \I__1878\ : InMux
    port map (
            O => \N__12121\,
            I => \N__12118\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__12118\,
            I => \N__12115\
        );

    \I__1876\ : Span4Mux_h
    port map (
            O => \N__12115\,
            I => \N__12112\
        );

    \I__1875\ : Span4Mux_h
    port map (
            O => \N__12112\,
            I => \N__12109\
        );

    \I__1874\ : Span4Mux_h
    port map (
            O => \N__12109\,
            I => \N__12106\
        );

    \I__1873\ : Odrv4
    port map (
            O => \N__12106\,
            I => \line_buffer.n448\
        );

    \I__1872\ : InMux
    port map (
            O => \N__12103\,
            I => \N__12100\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__12100\,
            I => \N__12097\
        );

    \I__1870\ : Span4Mux_v
    port map (
            O => \N__12097\,
            I => \N__12094\
        );

    \I__1869\ : Span4Mux_h
    port map (
            O => \N__12094\,
            I => \N__12091\
        );

    \I__1868\ : Odrv4
    port map (
            O => \N__12091\,
            I => \line_buffer.n440\
        );

    \I__1867\ : InMux
    port map (
            O => \N__12088\,
            I => \N__12085\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__12085\,
            I => \N__12082\
        );

    \I__1865\ : Odrv12
    port map (
            O => \N__12082\,
            I => \line_buffer.n3679\
        );

    \I__1864\ : InMux
    port map (
            O => \N__12079\,
            I => \N__12075\
        );

    \I__1863\ : InMux
    port map (
            O => \N__12078\,
            I => \N__12072\
        );

    \I__1862\ : LocalMux
    port map (
            O => \N__12075\,
            I => \N__12069\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__12072\,
            I => \N__12066\
        );

    \I__1860\ : Span4Mux_v
    port map (
            O => \N__12069\,
            I => \N__12063\
        );

    \I__1859\ : Span4Mux_v
    port map (
            O => \N__12066\,
            I => \N__12060\
        );

    \I__1858\ : Span4Mux_v
    port map (
            O => \N__12063\,
            I => \N__12057\
        );

    \I__1857\ : Odrv4
    port map (
            O => \N__12060\,
            I => \transmit_module.n116\
        );

    \I__1856\ : Odrv4
    port map (
            O => \N__12057\,
            I => \transmit_module.n116\
        );

    \I__1855\ : InMux
    port map (
            O => \N__12052\,
            I => \N__12048\
        );

    \I__1854\ : InMux
    port map (
            O => \N__12051\,
            I => \N__12045\
        );

    \I__1853\ : LocalMux
    port map (
            O => \N__12048\,
            I => \N__12042\
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__12045\,
            I => \N__12039\
        );

    \I__1851\ : Span12Mux_v
    port map (
            O => \N__12042\,
            I => \N__12036\
        );

    \I__1850\ : Odrv4
    port map (
            O => \N__12039\,
            I => \transmit_module.n147\
        );

    \I__1849\ : Odrv12
    port map (
            O => \N__12036\,
            I => \transmit_module.n147\
        );

    \I__1848\ : CascadeMux
    port map (
            O => \N__12031\,
            I => \N__12028\
        );

    \I__1847\ : CascadeBuf
    port map (
            O => \N__12028\,
            I => \N__12024\
        );

    \I__1846\ : CascadeMux
    port map (
            O => \N__12027\,
            I => \N__12021\
        );

    \I__1845\ : CascadeMux
    port map (
            O => \N__12024\,
            I => \N__12018\
        );

    \I__1844\ : CascadeBuf
    port map (
            O => \N__12021\,
            I => \N__12015\
        );

    \I__1843\ : CascadeBuf
    port map (
            O => \N__12018\,
            I => \N__12012\
        );

    \I__1842\ : CascadeMux
    port map (
            O => \N__12015\,
            I => \N__12009\
        );

    \I__1841\ : CascadeMux
    port map (
            O => \N__12012\,
            I => \N__12006\
        );

    \I__1840\ : CascadeBuf
    port map (
            O => \N__12009\,
            I => \N__12003\
        );

    \I__1839\ : CascadeBuf
    port map (
            O => \N__12006\,
            I => \N__12000\
        );

    \I__1838\ : CascadeMux
    port map (
            O => \N__12003\,
            I => \N__11997\
        );

    \I__1837\ : CascadeMux
    port map (
            O => \N__12000\,
            I => \N__11994\
        );

    \I__1836\ : CascadeBuf
    port map (
            O => \N__11997\,
            I => \N__11991\
        );

    \I__1835\ : CascadeBuf
    port map (
            O => \N__11994\,
            I => \N__11988\
        );

    \I__1834\ : CascadeMux
    port map (
            O => \N__11991\,
            I => \N__11985\
        );

    \I__1833\ : CascadeMux
    port map (
            O => \N__11988\,
            I => \N__11982\
        );

    \I__1832\ : CascadeBuf
    port map (
            O => \N__11985\,
            I => \N__11979\
        );

    \I__1831\ : CascadeBuf
    port map (
            O => \N__11982\,
            I => \N__11976\
        );

    \I__1830\ : CascadeMux
    port map (
            O => \N__11979\,
            I => \N__11973\
        );

    \I__1829\ : CascadeMux
    port map (
            O => \N__11976\,
            I => \N__11970\
        );

    \I__1828\ : CascadeBuf
    port map (
            O => \N__11973\,
            I => \N__11967\
        );

    \I__1827\ : CascadeBuf
    port map (
            O => \N__11970\,
            I => \N__11964\
        );

    \I__1826\ : CascadeMux
    port map (
            O => \N__11967\,
            I => \N__11961\
        );

    \I__1825\ : CascadeMux
    port map (
            O => \N__11964\,
            I => \N__11958\
        );

    \I__1824\ : CascadeBuf
    port map (
            O => \N__11961\,
            I => \N__11955\
        );

    \I__1823\ : CascadeBuf
    port map (
            O => \N__11958\,
            I => \N__11952\
        );

    \I__1822\ : CascadeMux
    port map (
            O => \N__11955\,
            I => \N__11949\
        );

    \I__1821\ : CascadeMux
    port map (
            O => \N__11952\,
            I => \N__11946\
        );

    \I__1820\ : CascadeBuf
    port map (
            O => \N__11949\,
            I => \N__11943\
        );

    \I__1819\ : CascadeBuf
    port map (
            O => \N__11946\,
            I => \N__11940\
        );

    \I__1818\ : CascadeMux
    port map (
            O => \N__11943\,
            I => \N__11937\
        );

    \I__1817\ : CascadeMux
    port map (
            O => \N__11940\,
            I => \N__11934\
        );

    \I__1816\ : CascadeBuf
    port map (
            O => \N__11937\,
            I => \N__11931\
        );

    \I__1815\ : CascadeBuf
    port map (
            O => \N__11934\,
            I => \N__11928\
        );

    \I__1814\ : CascadeMux
    port map (
            O => \N__11931\,
            I => \N__11925\
        );

    \I__1813\ : CascadeMux
    port map (
            O => \N__11928\,
            I => \N__11922\
        );

    \I__1812\ : CascadeBuf
    port map (
            O => \N__11925\,
            I => \N__11919\
        );

    \I__1811\ : CascadeBuf
    port map (
            O => \N__11922\,
            I => \N__11916\
        );

    \I__1810\ : CascadeMux
    port map (
            O => \N__11919\,
            I => \N__11913\
        );

    \I__1809\ : CascadeMux
    port map (
            O => \N__11916\,
            I => \N__11910\
        );

    \I__1808\ : CascadeBuf
    port map (
            O => \N__11913\,
            I => \N__11907\
        );

    \I__1807\ : CascadeBuf
    port map (
            O => \N__11910\,
            I => \N__11904\
        );

    \I__1806\ : CascadeMux
    port map (
            O => \N__11907\,
            I => \N__11901\
        );

    \I__1805\ : CascadeMux
    port map (
            O => \N__11904\,
            I => \N__11898\
        );

    \I__1804\ : CascadeBuf
    port map (
            O => \N__11901\,
            I => \N__11895\
        );

    \I__1803\ : CascadeBuf
    port map (
            O => \N__11898\,
            I => \N__11892\
        );

    \I__1802\ : CascadeMux
    port map (
            O => \N__11895\,
            I => \N__11889\
        );

    \I__1801\ : CascadeMux
    port map (
            O => \N__11892\,
            I => \N__11886\
        );

    \I__1800\ : CascadeBuf
    port map (
            O => \N__11889\,
            I => \N__11883\
        );

    \I__1799\ : CascadeBuf
    port map (
            O => \N__11886\,
            I => \N__11880\
        );

    \I__1798\ : CascadeMux
    port map (
            O => \N__11883\,
            I => \N__11877\
        );

    \I__1797\ : CascadeMux
    port map (
            O => \N__11880\,
            I => \N__11874\
        );

    \I__1796\ : CascadeBuf
    port map (
            O => \N__11877\,
            I => \N__11871\
        );

    \I__1795\ : CascadeBuf
    port map (
            O => \N__11874\,
            I => \N__11868\
        );

    \I__1794\ : CascadeMux
    port map (
            O => \N__11871\,
            I => \N__11865\
        );

    \I__1793\ : CascadeMux
    port map (
            O => \N__11868\,
            I => \N__11862\
        );

    \I__1792\ : CascadeBuf
    port map (
            O => \N__11865\,
            I => \N__11859\
        );

    \I__1791\ : CascadeBuf
    port map (
            O => \N__11862\,
            I => \N__11856\
        );

    \I__1790\ : CascadeMux
    port map (
            O => \N__11859\,
            I => \N__11853\
        );

    \I__1789\ : CascadeMux
    port map (
            O => \N__11856\,
            I => \N__11850\
        );

    \I__1788\ : CascadeBuf
    port map (
            O => \N__11853\,
            I => \N__11847\
        );

    \I__1787\ : InMux
    port map (
            O => \N__11850\,
            I => \N__11844\
        );

    \I__1786\ : CascadeMux
    port map (
            O => \N__11847\,
            I => \N__11841\
        );

    \I__1785\ : LocalMux
    port map (
            O => \N__11844\,
            I => \N__11838\
        );

    \I__1784\ : InMux
    port map (
            O => \N__11841\,
            I => \N__11835\
        );

    \I__1783\ : Span4Mux_v
    port map (
            O => \N__11838\,
            I => \N__11832\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__11835\,
            I => \N__11829\
        );

    \I__1781\ : Span4Mux_h
    port map (
            O => \N__11832\,
            I => \N__11826\
        );

    \I__1780\ : Span4Mux_h
    port map (
            O => \N__11829\,
            I => \N__11823\
        );

    \I__1779\ : Span4Mux_h
    port map (
            O => \N__11826\,
            I => \N__11820\
        );

    \I__1778\ : Span4Mux_v
    port map (
            O => \N__11823\,
            I => \N__11817\
        );

    \I__1777\ : Odrv4
    port map (
            O => \N__11820\,
            I => n28
        );

    \I__1776\ : Odrv4
    port map (
            O => \N__11817\,
            I => n28
        );

    \I__1775\ : InMux
    port map (
            O => \N__11812\,
            I => \N__11809\
        );

    \I__1774\ : LocalMux
    port map (
            O => \N__11809\,
            I => \transmit_module.n146\
        );

    \I__1773\ : CascadeMux
    port map (
            O => \N__11806\,
            I => \transmit_module.n146_cascade_\
        );

    \I__1772\ : InMux
    port map (
            O => \N__11803\,
            I => \N__11799\
        );

    \I__1771\ : InMux
    port map (
            O => \N__11802\,
            I => \N__11796\
        );

    \I__1770\ : LocalMux
    port map (
            O => \N__11799\,
            I => \N__11793\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__11796\,
            I => \transmit_module.n115\
        );

    \I__1768\ : Odrv4
    port map (
            O => \N__11793\,
            I => \transmit_module.n115\
        );

    \I__1767\ : CascadeMux
    port map (
            O => \N__11788\,
            I => \N__11785\
        );

    \I__1766\ : CascadeBuf
    port map (
            O => \N__11785\,
            I => \N__11781\
        );

    \I__1765\ : CascadeMux
    port map (
            O => \N__11784\,
            I => \N__11778\
        );

    \I__1764\ : CascadeMux
    port map (
            O => \N__11781\,
            I => \N__11775\
        );

    \I__1763\ : CascadeBuf
    port map (
            O => \N__11778\,
            I => \N__11772\
        );

    \I__1762\ : CascadeBuf
    port map (
            O => \N__11775\,
            I => \N__11769\
        );

    \I__1761\ : CascadeMux
    port map (
            O => \N__11772\,
            I => \N__11766\
        );

    \I__1760\ : CascadeMux
    port map (
            O => \N__11769\,
            I => \N__11763\
        );

    \I__1759\ : CascadeBuf
    port map (
            O => \N__11766\,
            I => \N__11760\
        );

    \I__1758\ : CascadeBuf
    port map (
            O => \N__11763\,
            I => \N__11757\
        );

    \I__1757\ : CascadeMux
    port map (
            O => \N__11760\,
            I => \N__11754\
        );

    \I__1756\ : CascadeMux
    port map (
            O => \N__11757\,
            I => \N__11751\
        );

    \I__1755\ : CascadeBuf
    port map (
            O => \N__11754\,
            I => \N__11748\
        );

    \I__1754\ : CascadeBuf
    port map (
            O => \N__11751\,
            I => \N__11745\
        );

    \I__1753\ : CascadeMux
    port map (
            O => \N__11748\,
            I => \N__11742\
        );

    \I__1752\ : CascadeMux
    port map (
            O => \N__11745\,
            I => \N__11739\
        );

    \I__1751\ : CascadeBuf
    port map (
            O => \N__11742\,
            I => \N__11736\
        );

    \I__1750\ : CascadeBuf
    port map (
            O => \N__11739\,
            I => \N__11733\
        );

    \I__1749\ : CascadeMux
    port map (
            O => \N__11736\,
            I => \N__11730\
        );

    \I__1748\ : CascadeMux
    port map (
            O => \N__11733\,
            I => \N__11727\
        );

    \I__1747\ : CascadeBuf
    port map (
            O => \N__11730\,
            I => \N__11724\
        );

    \I__1746\ : CascadeBuf
    port map (
            O => \N__11727\,
            I => \N__11721\
        );

    \I__1745\ : CascadeMux
    port map (
            O => \N__11724\,
            I => \N__11718\
        );

    \I__1744\ : CascadeMux
    port map (
            O => \N__11721\,
            I => \N__11715\
        );

    \I__1743\ : CascadeBuf
    port map (
            O => \N__11718\,
            I => \N__11712\
        );

    \I__1742\ : CascadeBuf
    port map (
            O => \N__11715\,
            I => \N__11709\
        );

    \I__1741\ : CascadeMux
    port map (
            O => \N__11712\,
            I => \N__11706\
        );

    \I__1740\ : CascadeMux
    port map (
            O => \N__11709\,
            I => \N__11703\
        );

    \I__1739\ : CascadeBuf
    port map (
            O => \N__11706\,
            I => \N__11700\
        );

    \I__1738\ : CascadeBuf
    port map (
            O => \N__11703\,
            I => \N__11697\
        );

    \I__1737\ : CascadeMux
    port map (
            O => \N__11700\,
            I => \N__11694\
        );

    \I__1736\ : CascadeMux
    port map (
            O => \N__11697\,
            I => \N__11691\
        );

    \I__1735\ : CascadeBuf
    port map (
            O => \N__11694\,
            I => \N__11688\
        );

    \I__1734\ : CascadeBuf
    port map (
            O => \N__11691\,
            I => \N__11685\
        );

    \I__1733\ : CascadeMux
    port map (
            O => \N__11688\,
            I => \N__11682\
        );

    \I__1732\ : CascadeMux
    port map (
            O => \N__11685\,
            I => \N__11679\
        );

    \I__1731\ : CascadeBuf
    port map (
            O => \N__11682\,
            I => \N__11676\
        );

    \I__1730\ : CascadeBuf
    port map (
            O => \N__11679\,
            I => \N__11673\
        );

    \I__1729\ : CascadeMux
    port map (
            O => \N__11676\,
            I => \N__11670\
        );

    \I__1728\ : CascadeMux
    port map (
            O => \N__11673\,
            I => \N__11667\
        );

    \I__1727\ : CascadeBuf
    port map (
            O => \N__11670\,
            I => \N__11664\
        );

    \I__1726\ : CascadeBuf
    port map (
            O => \N__11667\,
            I => \N__11661\
        );

    \I__1725\ : CascadeMux
    port map (
            O => \N__11664\,
            I => \N__11658\
        );

    \I__1724\ : CascadeMux
    port map (
            O => \N__11661\,
            I => \N__11655\
        );

    \I__1723\ : CascadeBuf
    port map (
            O => \N__11658\,
            I => \N__11652\
        );

    \I__1722\ : CascadeBuf
    port map (
            O => \N__11655\,
            I => \N__11649\
        );

    \I__1721\ : CascadeMux
    port map (
            O => \N__11652\,
            I => \N__11646\
        );

    \I__1720\ : CascadeMux
    port map (
            O => \N__11649\,
            I => \N__11643\
        );

    \I__1719\ : CascadeBuf
    port map (
            O => \N__11646\,
            I => \N__11640\
        );

    \I__1718\ : CascadeBuf
    port map (
            O => \N__11643\,
            I => \N__11637\
        );

    \I__1717\ : CascadeMux
    port map (
            O => \N__11640\,
            I => \N__11634\
        );

    \I__1716\ : CascadeMux
    port map (
            O => \N__11637\,
            I => \N__11631\
        );

    \I__1715\ : CascadeBuf
    port map (
            O => \N__11634\,
            I => \N__11628\
        );

    \I__1714\ : CascadeBuf
    port map (
            O => \N__11631\,
            I => \N__11625\
        );

    \I__1713\ : CascadeMux
    port map (
            O => \N__11628\,
            I => \N__11622\
        );

    \I__1712\ : CascadeMux
    port map (
            O => \N__11625\,
            I => \N__11619\
        );

    \I__1711\ : CascadeBuf
    port map (
            O => \N__11622\,
            I => \N__11616\
        );

    \I__1710\ : CascadeBuf
    port map (
            O => \N__11619\,
            I => \N__11613\
        );

    \I__1709\ : CascadeMux
    port map (
            O => \N__11616\,
            I => \N__11610\
        );

    \I__1708\ : CascadeMux
    port map (
            O => \N__11613\,
            I => \N__11607\
        );

    \I__1707\ : CascadeBuf
    port map (
            O => \N__11610\,
            I => \N__11604\
        );

    \I__1706\ : InMux
    port map (
            O => \N__11607\,
            I => \N__11601\
        );

    \I__1705\ : CascadeMux
    port map (
            O => \N__11604\,
            I => \N__11598\
        );

    \I__1704\ : LocalMux
    port map (
            O => \N__11601\,
            I => \N__11595\
        );

    \I__1703\ : InMux
    port map (
            O => \N__11598\,
            I => \N__11592\
        );

    \I__1702\ : Span4Mux_v
    port map (
            O => \N__11595\,
            I => \N__11589\
        );

    \I__1701\ : LocalMux
    port map (
            O => \N__11592\,
            I => \N__11586\
        );

    \I__1700\ : Span4Mux_v
    port map (
            O => \N__11589\,
            I => \N__11583\
        );

    \I__1699\ : Span4Mux_v
    port map (
            O => \N__11586\,
            I => \N__11580\
        );

    \I__1698\ : Span4Mux_v
    port map (
            O => \N__11583\,
            I => \N__11577\
        );

    \I__1697\ : Span4Mux_v
    port map (
            O => \N__11580\,
            I => \N__11574\
        );

    \I__1696\ : Span4Mux_v
    port map (
            O => \N__11577\,
            I => \N__11571\
        );

    \I__1695\ : Span4Mux_v
    port map (
            O => \N__11574\,
            I => \N__11568\
        );

    \I__1694\ : Span4Mux_h
    port map (
            O => \N__11571\,
            I => \N__11565\
        );

    \I__1693\ : Span4Mux_v
    port map (
            O => \N__11568\,
            I => \N__11562\
        );

    \I__1692\ : Span4Mux_h
    port map (
            O => \N__11565\,
            I => \N__11557\
        );

    \I__1691\ : Span4Mux_h
    port map (
            O => \N__11562\,
            I => \N__11557\
        );

    \I__1690\ : Odrv4
    port map (
            O => \N__11557\,
            I => n27
        );

    \I__1689\ : InMux
    port map (
            O => \N__11554\,
            I => \N__11551\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__11551\,
            I => \N__11548\
        );

    \I__1687\ : Odrv4
    port map (
            O => \N__11548\,
            I => \transmit_module.Y_DELTA_PATTERN_2\
        );

    \I__1686\ : InMux
    port map (
            O => \N__11545\,
            I => \N__11542\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__11542\,
            I => \transmit_module.Y_DELTA_PATTERN_1\
        );

    \I__1684\ : InMux
    port map (
            O => \N__11539\,
            I => \N__11536\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__11536\,
            I => \transmit_module.Y_DELTA_PATTERN_9\
        );

    \I__1682\ : InMux
    port map (
            O => \N__11533\,
            I => \N__11530\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__11530\,
            I => \N__11527\
        );

    \I__1680\ : Odrv12
    port map (
            O => \N__11527\,
            I => \transmit_module.Y_DELTA_PATTERN_8\
        );

    \I__1679\ : InMux
    port map (
            O => \N__11524\,
            I => \N__11521\
        );

    \I__1678\ : LocalMux
    port map (
            O => \N__11521\,
            I => \transmit_module.Y_DELTA_PATTERN_10\
        );

    \I__1677\ : InMux
    port map (
            O => \N__11518\,
            I => \N__11515\
        );

    \I__1676\ : LocalMux
    port map (
            O => \N__11515\,
            I => \N__11512\
        );

    \I__1675\ : Span4Mux_h
    port map (
            O => \N__11512\,
            I => \N__11509\
        );

    \I__1674\ : Span4Mux_h
    port map (
            O => \N__11509\,
            I => \N__11506\
        );

    \I__1673\ : Span4Mux_v
    port map (
            O => \N__11506\,
            I => \N__11503\
        );

    \I__1672\ : Span4Mux_v
    port map (
            O => \N__11503\,
            I => \N__11500\
        );

    \I__1671\ : Odrv4
    port map (
            O => \N__11500\,
            I => \line_buffer.n507\
        );

    \I__1670\ : CascadeMux
    port map (
            O => \N__11497\,
            I => \N__11494\
        );

    \I__1669\ : InMux
    port map (
            O => \N__11494\,
            I => \N__11491\
        );

    \I__1668\ : LocalMux
    port map (
            O => \N__11491\,
            I => \N__11488\
        );

    \I__1667\ : Span4Mux_v
    port map (
            O => \N__11488\,
            I => \N__11485\
        );

    \I__1666\ : Sp12to4
    port map (
            O => \N__11485\,
            I => \N__11482\
        );

    \I__1665\ : Span12Mux_h
    port map (
            O => \N__11482\,
            I => \N__11479\
        );

    \I__1664\ : Odrv12
    port map (
            O => \N__11479\,
            I => \line_buffer.n499\
        );

    \I__1663\ : InMux
    port map (
            O => \N__11476\,
            I => \N__11473\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__11473\,
            I => \line_buffer.n3752\
        );

    \I__1661\ : CascadeMux
    port map (
            O => \N__11470\,
            I => \transmit_module.n141_cascade_\
        );

    \I__1660\ : CascadeMux
    port map (
            O => \N__11467\,
            I => \transmit_module.n137_cascade_\
        );

    \I__1659\ : CascadeMux
    port map (
            O => \N__11464\,
            I => \N__11461\
        );

    \I__1658\ : InMux
    port map (
            O => \N__11461\,
            I => \N__11458\
        );

    \I__1657\ : LocalMux
    port map (
            O => \N__11458\,
            I => \transmit_module.ADDR_Y_COMPONENT_1\
        );

    \I__1656\ : CascadeMux
    port map (
            O => \N__11455\,
            I => \N__11452\
        );

    \I__1655\ : InMux
    port map (
            O => \N__11452\,
            I => \N__11449\
        );

    \I__1654\ : LocalMux
    port map (
            O => \N__11449\,
            I => \transmit_module.ADDR_Y_COMPONENT_10\
        );

    \I__1653\ : InMux
    port map (
            O => \N__11446\,
            I => \N__11443\
        );

    \I__1652\ : LocalMux
    port map (
            O => \N__11443\,
            I => \transmit_module.video_signal_controller.n3632\
        );

    \I__1651\ : InMux
    port map (
            O => \N__11440\,
            I => \N__11437\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__11437\,
            I => \N__11434\
        );

    \I__1649\ : Odrv4
    port map (
            O => \N__11434\,
            I => \transmit_module.video_signal_controller.n18_adj_616\
        );

    \I__1648\ : CascadeMux
    port map (
            O => \N__11431\,
            I => \N__11428\
        );

    \I__1647\ : InMux
    port map (
            O => \N__11428\,
            I => \N__11425\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__11425\,
            I => \transmit_module.video_signal_controller.n3614\
        );

    \I__1645\ : InMux
    port map (
            O => \N__11422\,
            I => \N__11419\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__11419\,
            I => \N__11416\
        );

    \I__1643\ : Span4Mux_h
    port map (
            O => \N__11416\,
            I => \N__11411\
        );

    \I__1642\ : InMux
    port map (
            O => \N__11415\,
            I => \N__11408\
        );

    \I__1641\ : InMux
    port map (
            O => \N__11414\,
            I => \N__11405\
        );

    \I__1640\ : Odrv4
    port map (
            O => \N__11411\,
            I => \transmit_module.video_signal_controller.VGA_Y_10\
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__11408\,
            I => \transmit_module.video_signal_controller.VGA_Y_10\
        );

    \I__1638\ : LocalMux
    port map (
            O => \N__11405\,
            I => \transmit_module.video_signal_controller.VGA_Y_10\
        );

    \I__1637\ : InMux
    port map (
            O => \N__11398\,
            I => \N__11395\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__11395\,
            I => \N__11392\
        );

    \I__1635\ : Span4Mux_h
    port map (
            O => \N__11392\,
            I => \N__11388\
        );

    \I__1634\ : InMux
    port map (
            O => \N__11391\,
            I => \N__11385\
        );

    \I__1633\ : Odrv4
    port map (
            O => \N__11388\,
            I => \transmit_module.video_signal_controller.VGA_Y_0\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__11385\,
            I => \transmit_module.video_signal_controller.VGA_Y_0\
        );

    \I__1631\ : InMux
    port map (
            O => \N__11380\,
            I => \N__11374\
        );

    \I__1630\ : InMux
    port map (
            O => \N__11379\,
            I => \N__11369\
        );

    \I__1629\ : InMux
    port map (
            O => \N__11378\,
            I => \N__11369\
        );

    \I__1628\ : InMux
    port map (
            O => \N__11377\,
            I => \N__11366\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__11374\,
            I => \N__11361\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__11369\,
            I => \N__11361\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__11366\,
            I => \transmit_module.video_signal_controller.VGA_Y_3\
        );

    \I__1624\ : Odrv4
    port map (
            O => \N__11361\,
            I => \transmit_module.video_signal_controller.VGA_Y_3\
        );

    \I__1623\ : CascadeMux
    port map (
            O => \N__11356\,
            I => \transmit_module.video_signal_controller.n3626_cascade_\
        );

    \I__1622\ : InMux
    port map (
            O => \N__11353\,
            I => \N__11349\
        );

    \I__1621\ : CascadeMux
    port map (
            O => \N__11352\,
            I => \N__11345\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__11349\,
            I => \N__11341\
        );

    \I__1619\ : InMux
    port map (
            O => \N__11348\,
            I => \N__11338\
        );

    \I__1618\ : InMux
    port map (
            O => \N__11345\,
            I => \N__11333\
        );

    \I__1617\ : InMux
    port map (
            O => \N__11344\,
            I => \N__11333\
        );

    \I__1616\ : Odrv4
    port map (
            O => \N__11341\,
            I => \transmit_module.video_signal_controller.VGA_Y_1\
        );

    \I__1615\ : LocalMux
    port map (
            O => \N__11338\,
            I => \transmit_module.video_signal_controller.VGA_Y_1\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__11333\,
            I => \transmit_module.video_signal_controller.VGA_Y_1\
        );

    \I__1613\ : InMux
    port map (
            O => \N__11326\,
            I => \N__11323\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__11323\,
            I => \N__11320\
        );

    \I__1611\ : Odrv4
    port map (
            O => \N__11320\,
            I => \transmit_module.n111\
        );

    \I__1610\ : InMux
    port map (
            O => \N__11317\,
            I => \N__11314\
        );

    \I__1609\ : LocalMux
    port map (
            O => \N__11314\,
            I => \N__11311\
        );

    \I__1608\ : Span4Mux_h
    port map (
            O => \N__11311\,
            I => \N__11308\
        );

    \I__1607\ : Odrv4
    port map (
            O => \N__11308\,
            I => \transmit_module.n143\
        );

    \I__1606\ : CascadeMux
    port map (
            O => \N__11305\,
            I => \transmit_module.n143_cascade_\
        );

    \I__1605\ : InMux
    port map (
            O => \N__11302\,
            I => \N__11299\
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__11299\,
            I => \transmit_module.n112\
        );

    \I__1603\ : InMux
    port map (
            O => \N__11296\,
            I => \N__11292\
        );

    \I__1602\ : InMux
    port map (
            O => \N__11295\,
            I => \N__11289\
        );

    \I__1601\ : LocalMux
    port map (
            O => \N__11292\,
            I => \transmit_module.n142\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__11289\,
            I => \transmit_module.n142\
        );

    \I__1599\ : InMux
    port map (
            O => \N__11284\,
            I => \N__11278\
        );

    \I__1598\ : InMux
    port map (
            O => \N__11283\,
            I => \N__11271\
        );

    \I__1597\ : InMux
    port map (
            O => \N__11282\,
            I => \N__11271\
        );

    \I__1596\ : InMux
    port map (
            O => \N__11281\,
            I => \N__11271\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__11278\,
            I => \receive_module.rx_counter.Y_3\
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__11271\,
            I => \receive_module.rx_counter.Y_3\
        );

    \I__1593\ : InMux
    port map (
            O => \N__11266\,
            I => \N__11260\
        );

    \I__1592\ : InMux
    port map (
            O => \N__11265\,
            I => \N__11253\
        );

    \I__1591\ : InMux
    port map (
            O => \N__11264\,
            I => \N__11253\
        );

    \I__1590\ : InMux
    port map (
            O => \N__11263\,
            I => \N__11253\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__11260\,
            I => \receive_module.rx_counter.Y_2\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__11253\,
            I => \receive_module.rx_counter.Y_2\
        );

    \I__1587\ : CascadeMux
    port map (
            O => \N__11248\,
            I => \N__11242\
        );

    \I__1586\ : InMux
    port map (
            O => \N__11247\,
            I => \N__11239\
        );

    \I__1585\ : InMux
    port map (
            O => \N__11246\,
            I => \N__11232\
        );

    \I__1584\ : InMux
    port map (
            O => \N__11245\,
            I => \N__11232\
        );

    \I__1583\ : InMux
    port map (
            O => \N__11242\,
            I => \N__11232\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__11239\,
            I => \receive_module.rx_counter.Y_1\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__11232\,
            I => \receive_module.rx_counter.Y_1\
        );

    \I__1580\ : InMux
    port map (
            O => \N__11227\,
            I => \N__11222\
        );

    \I__1579\ : InMux
    port map (
            O => \N__11226\,
            I => \N__11217\
        );

    \I__1578\ : InMux
    port map (
            O => \N__11225\,
            I => \N__11217\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__11222\,
            I => \receive_module.rx_counter.Y_5\
        );

    \I__1576\ : LocalMux
    port map (
            O => \N__11217\,
            I => \receive_module.rx_counter.Y_5\
        );

    \I__1575\ : InMux
    port map (
            O => \N__11212\,
            I => \N__11207\
        );

    \I__1574\ : InMux
    port map (
            O => \N__11211\,
            I => \N__11204\
        );

    \I__1573\ : InMux
    port map (
            O => \N__11210\,
            I => \N__11201\
        );

    \I__1572\ : LocalMux
    port map (
            O => \N__11207\,
            I => \receive_module.rx_counter.Y_6\
        );

    \I__1571\ : LocalMux
    port map (
            O => \N__11204\,
            I => \receive_module.rx_counter.Y_6\
        );

    \I__1570\ : LocalMux
    port map (
            O => \N__11201\,
            I => \receive_module.rx_counter.Y_6\
        );

    \I__1569\ : InMux
    port map (
            O => \N__11194\,
            I => \N__11191\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__11191\,
            I => \receive_module.rx_counter.n4_adj_604\
        );

    \I__1567\ : CascadeMux
    port map (
            O => \N__11188\,
            I => \receive_module.rx_counter.n5_cascade_\
        );

    \I__1566\ : InMux
    port map (
            O => \N__11185\,
            I => \N__11182\
        );

    \I__1565\ : LocalMux
    port map (
            O => \N__11182\,
            I => \receive_module.rx_counter.n3548\
        );

    \I__1564\ : InMux
    port map (
            O => \N__11179\,
            I => \N__11173\
        );

    \I__1563\ : InMux
    port map (
            O => \N__11178\,
            I => \N__11170\
        );

    \I__1562\ : InMux
    port map (
            O => \N__11177\,
            I => \N__11165\
        );

    \I__1561\ : InMux
    port map (
            O => \N__11176\,
            I => \N__11165\
        );

    \I__1560\ : LocalMux
    port map (
            O => \N__11173\,
            I => \receive_module.rx_counter.Y_0\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__11170\,
            I => \receive_module.rx_counter.Y_0\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__11165\,
            I => \receive_module.rx_counter.Y_0\
        );

    \I__1557\ : InMux
    port map (
            O => \N__11158\,
            I => \N__11155\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__11155\,
            I => \receive_module.rx_counter.n14_adj_611\
        );

    \I__1555\ : CascadeMux
    port map (
            O => \N__11152\,
            I => \N__11149\
        );

    \I__1554\ : InMux
    port map (
            O => \N__11149\,
            I => \N__11146\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__11146\,
            I => \receive_module.rx_counter.n10_adj_610\
        );

    \I__1552\ : InMux
    port map (
            O => \N__11143\,
            I => \N__11140\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__11140\,
            I => \transmit_module.ADDR_Y_COMPONENT_7\
        );

    \I__1550\ : InMux
    port map (
            O => \N__11137\,
            I => \N__11134\
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__11134\,
            I => \N__11131\
        );

    \I__1548\ : Odrv12
    port map (
            O => \N__11131\,
            I => \transmit_module.X_DELTA_PATTERN_1\
        );

    \I__1547\ : CEMux
    port map (
            O => \N__11128\,
            I => \N__11124\
        );

    \I__1546\ : CEMux
    port map (
            O => \N__11127\,
            I => \N__11119\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__11124\,
            I => \N__11116\
        );

    \I__1544\ : CEMux
    port map (
            O => \N__11123\,
            I => \N__11113\
        );

    \I__1543\ : CEMux
    port map (
            O => \N__11122\,
            I => \N__11110\
        );

    \I__1542\ : LocalMux
    port map (
            O => \N__11119\,
            I => \N__11107\
        );

    \I__1541\ : Span4Mux_h
    port map (
            O => \N__11116\,
            I => \N__11103\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__11113\,
            I => \N__11100\
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__11110\,
            I => \N__11097\
        );

    \I__1538\ : Span4Mux_v
    port map (
            O => \N__11107\,
            I => \N__11094\
        );

    \I__1537\ : CEMux
    port map (
            O => \N__11106\,
            I => \N__11091\
        );

    \I__1536\ : Span4Mux_h
    port map (
            O => \N__11103\,
            I => \N__11086\
        );

    \I__1535\ : Span4Mux_h
    port map (
            O => \N__11100\,
            I => \N__11086\
        );

    \I__1534\ : Span4Mux_h
    port map (
            O => \N__11097\,
            I => \N__11079\
        );

    \I__1533\ : Span4Mux_h
    port map (
            O => \N__11094\,
            I => \N__11079\
        );

    \I__1532\ : LocalMux
    port map (
            O => \N__11091\,
            I => \N__11079\
        );

    \I__1531\ : Odrv4
    port map (
            O => \N__11086\,
            I => \transmit_module.n2093\
        );

    \I__1530\ : Odrv4
    port map (
            O => \N__11079\,
            I => \transmit_module.n2093\
        );

    \I__1529\ : CEMux
    port map (
            O => \N__11074\,
            I => \N__11070\
        );

    \I__1528\ : CEMux
    port map (
            O => \N__11073\,
            I => \N__11066\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__11070\,
            I => \N__11061\
        );

    \I__1526\ : CEMux
    port map (
            O => \N__11069\,
            I => \N__11058\
        );

    \I__1525\ : LocalMux
    port map (
            O => \N__11066\,
            I => \N__11055\
        );

    \I__1524\ : CEMux
    port map (
            O => \N__11065\,
            I => \N__11052\
        );

    \I__1523\ : SRMux
    port map (
            O => \N__11064\,
            I => \N__11049\
        );

    \I__1522\ : Span4Mux_v
    port map (
            O => \N__11061\,
            I => \N__11044\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__11058\,
            I => \N__11044\
        );

    \I__1520\ : Span4Mux_v
    port map (
            O => \N__11055\,
            I => \N__11041\
        );

    \I__1519\ : LocalMux
    port map (
            O => \N__11052\,
            I => \N__11038\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__11049\,
            I => \N__11035\
        );

    \I__1517\ : Span4Mux_v
    port map (
            O => \N__11044\,
            I => \N__11032\
        );

    \I__1516\ : Span4Mux_h
    port map (
            O => \N__11041\,
            I => \N__11027\
        );

    \I__1515\ : Span4Mux_v
    port map (
            O => \N__11038\,
            I => \N__11027\
        );

    \I__1514\ : Span4Mux_v
    port map (
            O => \N__11035\,
            I => \N__11024\
        );

    \I__1513\ : Odrv4
    port map (
            O => \N__11032\,
            I => \transmit_module.n2147\
        );

    \I__1512\ : Odrv4
    port map (
            O => \N__11027\,
            I => \transmit_module.n2147\
        );

    \I__1511\ : Odrv4
    port map (
            O => \N__11024\,
            I => \transmit_module.n2147\
        );

    \I__1510\ : InMux
    port map (
            O => \N__11017\,
            I => \N__11013\
        );

    \I__1509\ : InMux
    port map (
            O => \N__11016\,
            I => \N__11008\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__11013\,
            I => \N__11005\
        );

    \I__1507\ : InMux
    port map (
            O => \N__11012\,
            I => \N__11000\
        );

    \I__1506\ : InMux
    port map (
            O => \N__11011\,
            I => \N__11000\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__11008\,
            I => \transmit_module.video_signal_controller.VGA_Y_4\
        );

    \I__1504\ : Odrv4
    port map (
            O => \N__11005\,
            I => \transmit_module.video_signal_controller.VGA_Y_4\
        );

    \I__1503\ : LocalMux
    port map (
            O => \N__11000\,
            I => \transmit_module.video_signal_controller.VGA_Y_4\
        );

    \I__1502\ : InMux
    port map (
            O => \N__10993\,
            I => \N__10989\
        );

    \I__1501\ : InMux
    port map (
            O => \N__10992\,
            I => \N__10985\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__10989\,
            I => \N__10982\
        );

    \I__1499\ : InMux
    port map (
            O => \N__10988\,
            I => \N__10978\
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__10985\,
            I => \N__10973\
        );

    \I__1497\ : Span4Mux_v
    port map (
            O => \N__10982\,
            I => \N__10973\
        );

    \I__1496\ : InMux
    port map (
            O => \N__10981\,
            I => \N__10970\
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__10978\,
            I => \transmit_module.video_signal_controller.VGA_Y_8\
        );

    \I__1494\ : Odrv4
    port map (
            O => \N__10973\,
            I => \transmit_module.video_signal_controller.VGA_Y_8\
        );

    \I__1493\ : LocalMux
    port map (
            O => \N__10970\,
            I => \transmit_module.video_signal_controller.VGA_Y_8\
        );

    \I__1492\ : InMux
    port map (
            O => \N__10963\,
            I => \N__10960\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__10960\,
            I => \transmit_module.ADDR_Y_COMPONENT_4\
        );

    \I__1490\ : InMux
    port map (
            O => \N__10957\,
            I => \N__10954\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__10954\,
            I => \transmit_module.ADDR_Y_COMPONENT_5\
        );

    \I__1488\ : InMux
    port map (
            O => \N__10951\,
            I => \N__10948\
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__10948\,
            I => \N__10945\
        );

    \I__1486\ : Span4Mux_v
    port map (
            O => \N__10945\,
            I => \N__10942\
        );

    \I__1485\ : Span4Mux_h
    port map (
            O => \N__10942\,
            I => \N__10939\
        );

    \I__1484\ : Odrv4
    port map (
            O => \N__10939\,
            I => \line_buffer.n571\
        );

    \I__1483\ : InMux
    port map (
            O => \N__10936\,
            I => \N__10933\
        );

    \I__1482\ : LocalMux
    port map (
            O => \N__10933\,
            I => \N__10930\
        );

    \I__1481\ : Span12Mux_v
    port map (
            O => \N__10930\,
            I => \N__10927\
        );

    \I__1480\ : Span12Mux_h
    port map (
            O => \N__10927\,
            I => \N__10924\
        );

    \I__1479\ : Odrv12
    port map (
            O => \N__10924\,
            I => \line_buffer.n563\
        );

    \I__1478\ : InMux
    port map (
            O => \N__10921\,
            I => \N__10918\
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__10918\,
            I => \N__10915\
        );

    \I__1476\ : Span4Mux_v
    port map (
            O => \N__10915\,
            I => \N__10912\
        );

    \I__1475\ : Span4Mux_h
    port map (
            O => \N__10912\,
            I => \N__10909\
        );

    \I__1474\ : Odrv4
    port map (
            O => \N__10909\,
            I => \line_buffer.n514\
        );

    \I__1473\ : CascadeMux
    port map (
            O => \N__10906\,
            I => \N__10903\
        );

    \I__1472\ : InMux
    port map (
            O => \N__10903\,
            I => \N__10900\
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__10900\,
            I => \N__10897\
        );

    \I__1470\ : Span12Mux_v
    port map (
            O => \N__10897\,
            I => \N__10894\
        );

    \I__1469\ : Span12Mux_v
    port map (
            O => \N__10894\,
            I => \N__10891\
        );

    \I__1468\ : Span12Mux_h
    port map (
            O => \N__10891\,
            I => \N__10888\
        );

    \I__1467\ : Odrv12
    port map (
            O => \N__10888\,
            I => \line_buffer.n506\
        );

    \I__1466\ : InMux
    port map (
            O => \N__10885\,
            I => \N__10882\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__10882\,
            I => \line_buffer.n3764\
        );

    \I__1464\ : InMux
    port map (
            O => \N__10879\,
            I => \N__10876\
        );

    \I__1463\ : LocalMux
    port map (
            O => \N__10876\,
            I => \N__10873\
        );

    \I__1462\ : Span4Mux_h
    port map (
            O => \N__10873\,
            I => \N__10870\
        );

    \I__1461\ : Span4Mux_h
    port map (
            O => \N__10870\,
            I => \N__10867\
        );

    \I__1460\ : Odrv4
    port map (
            O => \N__10867\,
            I => \line_buffer.n513\
        );

    \I__1459\ : InMux
    port map (
            O => \N__10864\,
            I => \N__10861\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__10861\,
            I => \N__10858\
        );

    \I__1457\ : Span12Mux_v
    port map (
            O => \N__10858\,
            I => \N__10855\
        );

    \I__1456\ : Span12Mux_v
    port map (
            O => \N__10855\,
            I => \N__10852\
        );

    \I__1455\ : Span12Mux_h
    port map (
            O => \N__10852\,
            I => \N__10849\
        );

    \I__1454\ : Odrv12
    port map (
            O => \N__10849\,
            I => \line_buffer.n505\
        );

    \I__1453\ : CascadeMux
    port map (
            O => \N__10846\,
            I => \line_buffer.n3646_cascade_\
        );

    \I__1452\ : InMux
    port map (
            O => \N__10843\,
            I => \N__10840\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__10840\,
            I => \line_buffer.n3647\
        );

    \I__1450\ : CascadeMux
    port map (
            O => \N__10837\,
            I => \transmit_module.n112_cascade_\
        );

    \I__1449\ : CascadeMux
    port map (
            O => \N__10834\,
            I => \N__10831\
        );

    \I__1448\ : CascadeBuf
    port map (
            O => \N__10831\,
            I => \N__10828\
        );

    \I__1447\ : CascadeMux
    port map (
            O => \N__10828\,
            I => \N__10824\
        );

    \I__1446\ : CascadeMux
    port map (
            O => \N__10827\,
            I => \N__10821\
        );

    \I__1445\ : CascadeBuf
    port map (
            O => \N__10824\,
            I => \N__10818\
        );

    \I__1444\ : CascadeBuf
    port map (
            O => \N__10821\,
            I => \N__10815\
        );

    \I__1443\ : CascadeMux
    port map (
            O => \N__10818\,
            I => \N__10812\
        );

    \I__1442\ : CascadeMux
    port map (
            O => \N__10815\,
            I => \N__10809\
        );

    \I__1441\ : CascadeBuf
    port map (
            O => \N__10812\,
            I => \N__10806\
        );

    \I__1440\ : CascadeBuf
    port map (
            O => \N__10809\,
            I => \N__10803\
        );

    \I__1439\ : CascadeMux
    port map (
            O => \N__10806\,
            I => \N__10800\
        );

    \I__1438\ : CascadeMux
    port map (
            O => \N__10803\,
            I => \N__10797\
        );

    \I__1437\ : CascadeBuf
    port map (
            O => \N__10800\,
            I => \N__10794\
        );

    \I__1436\ : CascadeBuf
    port map (
            O => \N__10797\,
            I => \N__10791\
        );

    \I__1435\ : CascadeMux
    port map (
            O => \N__10794\,
            I => \N__10788\
        );

    \I__1434\ : CascadeMux
    port map (
            O => \N__10791\,
            I => \N__10785\
        );

    \I__1433\ : CascadeBuf
    port map (
            O => \N__10788\,
            I => \N__10782\
        );

    \I__1432\ : CascadeBuf
    port map (
            O => \N__10785\,
            I => \N__10779\
        );

    \I__1431\ : CascadeMux
    port map (
            O => \N__10782\,
            I => \N__10776\
        );

    \I__1430\ : CascadeMux
    port map (
            O => \N__10779\,
            I => \N__10773\
        );

    \I__1429\ : CascadeBuf
    port map (
            O => \N__10776\,
            I => \N__10770\
        );

    \I__1428\ : CascadeBuf
    port map (
            O => \N__10773\,
            I => \N__10767\
        );

    \I__1427\ : CascadeMux
    port map (
            O => \N__10770\,
            I => \N__10764\
        );

    \I__1426\ : CascadeMux
    port map (
            O => \N__10767\,
            I => \N__10761\
        );

    \I__1425\ : CascadeBuf
    port map (
            O => \N__10764\,
            I => \N__10758\
        );

    \I__1424\ : CascadeBuf
    port map (
            O => \N__10761\,
            I => \N__10755\
        );

    \I__1423\ : CascadeMux
    port map (
            O => \N__10758\,
            I => \N__10752\
        );

    \I__1422\ : CascadeMux
    port map (
            O => \N__10755\,
            I => \N__10749\
        );

    \I__1421\ : CascadeBuf
    port map (
            O => \N__10752\,
            I => \N__10746\
        );

    \I__1420\ : CascadeBuf
    port map (
            O => \N__10749\,
            I => \N__10743\
        );

    \I__1419\ : CascadeMux
    port map (
            O => \N__10746\,
            I => \N__10740\
        );

    \I__1418\ : CascadeMux
    port map (
            O => \N__10743\,
            I => \N__10737\
        );

    \I__1417\ : CascadeBuf
    port map (
            O => \N__10740\,
            I => \N__10734\
        );

    \I__1416\ : CascadeBuf
    port map (
            O => \N__10737\,
            I => \N__10731\
        );

    \I__1415\ : CascadeMux
    port map (
            O => \N__10734\,
            I => \N__10728\
        );

    \I__1414\ : CascadeMux
    port map (
            O => \N__10731\,
            I => \N__10725\
        );

    \I__1413\ : CascadeBuf
    port map (
            O => \N__10728\,
            I => \N__10722\
        );

    \I__1412\ : CascadeBuf
    port map (
            O => \N__10725\,
            I => \N__10719\
        );

    \I__1411\ : CascadeMux
    port map (
            O => \N__10722\,
            I => \N__10716\
        );

    \I__1410\ : CascadeMux
    port map (
            O => \N__10719\,
            I => \N__10713\
        );

    \I__1409\ : CascadeBuf
    port map (
            O => \N__10716\,
            I => \N__10710\
        );

    \I__1408\ : CascadeBuf
    port map (
            O => \N__10713\,
            I => \N__10707\
        );

    \I__1407\ : CascadeMux
    port map (
            O => \N__10710\,
            I => \N__10704\
        );

    \I__1406\ : CascadeMux
    port map (
            O => \N__10707\,
            I => \N__10701\
        );

    \I__1405\ : CascadeBuf
    port map (
            O => \N__10704\,
            I => \N__10698\
        );

    \I__1404\ : CascadeBuf
    port map (
            O => \N__10701\,
            I => \N__10695\
        );

    \I__1403\ : CascadeMux
    port map (
            O => \N__10698\,
            I => \N__10692\
        );

    \I__1402\ : CascadeMux
    port map (
            O => \N__10695\,
            I => \N__10689\
        );

    \I__1401\ : CascadeBuf
    port map (
            O => \N__10692\,
            I => \N__10686\
        );

    \I__1400\ : CascadeBuf
    port map (
            O => \N__10689\,
            I => \N__10683\
        );

    \I__1399\ : CascadeMux
    port map (
            O => \N__10686\,
            I => \N__10680\
        );

    \I__1398\ : CascadeMux
    port map (
            O => \N__10683\,
            I => \N__10677\
        );

    \I__1397\ : CascadeBuf
    port map (
            O => \N__10680\,
            I => \N__10674\
        );

    \I__1396\ : CascadeBuf
    port map (
            O => \N__10677\,
            I => \N__10671\
        );

    \I__1395\ : CascadeMux
    port map (
            O => \N__10674\,
            I => \N__10668\
        );

    \I__1394\ : CascadeMux
    port map (
            O => \N__10671\,
            I => \N__10665\
        );

    \I__1393\ : CascadeBuf
    port map (
            O => \N__10668\,
            I => \N__10662\
        );

    \I__1392\ : CascadeBuf
    port map (
            O => \N__10665\,
            I => \N__10659\
        );

    \I__1391\ : CascadeMux
    port map (
            O => \N__10662\,
            I => \N__10656\
        );

    \I__1390\ : CascadeMux
    port map (
            O => \N__10659\,
            I => \N__10653\
        );

    \I__1389\ : InMux
    port map (
            O => \N__10656\,
            I => \N__10650\
        );

    \I__1388\ : CascadeBuf
    port map (
            O => \N__10653\,
            I => \N__10647\
        );

    \I__1387\ : LocalMux
    port map (
            O => \N__10650\,
            I => \N__10644\
        );

    \I__1386\ : CascadeMux
    port map (
            O => \N__10647\,
            I => \N__10641\
        );

    \I__1385\ : Span4Mux_s3_v
    port map (
            O => \N__10644\,
            I => \N__10638\
        );

    \I__1384\ : InMux
    port map (
            O => \N__10641\,
            I => \N__10635\
        );

    \I__1383\ : Span4Mux_h
    port map (
            O => \N__10638\,
            I => \N__10632\
        );

    \I__1382\ : LocalMux
    port map (
            O => \N__10635\,
            I => \N__10629\
        );

    \I__1381\ : Span4Mux_v
    port map (
            O => \N__10632\,
            I => \N__10626\
        );

    \I__1380\ : Span12Mux_s7_v
    port map (
            O => \N__10629\,
            I => \N__10623\
        );

    \I__1379\ : Sp12to4
    port map (
            O => \N__10626\,
            I => \N__10618\
        );

    \I__1378\ : Span12Mux_h
    port map (
            O => \N__10623\,
            I => \N__10618\
        );

    \I__1377\ : Odrv12
    port map (
            O => \N__10618\,
            I => n24
        );

    \I__1376\ : CascadeMux
    port map (
            O => \N__10615\,
            I => \N__10610\
        );

    \I__1375\ : InMux
    port map (
            O => \N__10614\,
            I => \N__10604\
        );

    \I__1374\ : InMux
    port map (
            O => \N__10613\,
            I => \N__10604\
        );

    \I__1373\ : InMux
    port map (
            O => \N__10610\,
            I => \N__10599\
        );

    \I__1372\ : InMux
    port map (
            O => \N__10609\,
            I => \N__10599\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__10604\,
            I => \transmit_module.old_VGA_HS\
        );

    \I__1370\ : LocalMux
    port map (
            O => \N__10599\,
            I => \transmit_module.old_VGA_HS\
        );

    \I__1369\ : CascadeMux
    port map (
            O => \N__10594\,
            I => \N__10591\
        );

    \I__1368\ : InMux
    port map (
            O => \N__10591\,
            I => \N__10585\
        );

    \I__1367\ : InMux
    port map (
            O => \N__10590\,
            I => \N__10585\
        );

    \I__1366\ : LocalMux
    port map (
            O => \N__10585\,
            I => \N__10580\
        );

    \I__1365\ : InMux
    port map (
            O => \N__10584\,
            I => \N__10575\
        );

    \I__1364\ : InMux
    port map (
            O => \N__10583\,
            I => \N__10575\
        );

    \I__1363\ : Odrv4
    port map (
            O => \N__10580\,
            I => \transmit_module.VGA_VISIBLE_Y\
        );

    \I__1362\ : LocalMux
    port map (
            O => \N__10575\,
            I => \transmit_module.VGA_VISIBLE_Y\
        );

    \I__1361\ : IoInMux
    port map (
            O => \N__10570\,
            I => \N__10567\
        );

    \I__1360\ : LocalMux
    port map (
            O => \N__10567\,
            I => \N__10564\
        );

    \I__1359\ : IoSpan4Mux
    port map (
            O => \N__10564\,
            I => \N__10561\
        );

    \I__1358\ : Span4Mux_s2_h
    port map (
            O => \N__10561\,
            I => \N__10558\
        );

    \I__1357\ : Span4Mux_h
    port map (
            O => \N__10558\,
            I => \N__10553\
        );

    \I__1356\ : InMux
    port map (
            O => \N__10557\,
            I => \N__10548\
        );

    \I__1355\ : InMux
    port map (
            O => \N__10556\,
            I => \N__10548\
        );

    \I__1354\ : Span4Mux_h
    port map (
            O => \N__10553\,
            I => \N__10542\
        );

    \I__1353\ : LocalMux
    port map (
            O => \N__10548\,
            I => \N__10539\
        );

    \I__1352\ : InMux
    port map (
            O => \N__10547\,
            I => \N__10532\
        );

    \I__1351\ : InMux
    port map (
            O => \N__10546\,
            I => \N__10532\
        );

    \I__1350\ : InMux
    port map (
            O => \N__10545\,
            I => \N__10532\
        );

    \I__1349\ : Odrv4
    port map (
            O => \N__10542\,
            I => \ADV_HSYNC_c\
        );

    \I__1348\ : Odrv4
    port map (
            O => \N__10539\,
            I => \ADV_HSYNC_c\
        );

    \I__1347\ : LocalMux
    port map (
            O => \N__10532\,
            I => \ADV_HSYNC_c\
        );

    \I__1346\ : InMux
    port map (
            O => \N__10525\,
            I => \N__10522\
        );

    \I__1345\ : LocalMux
    port map (
            O => \N__10522\,
            I => \N__10518\
        );

    \I__1344\ : InMux
    port map (
            O => \N__10521\,
            I => \N__10515\
        );

    \I__1343\ : Odrv4
    port map (
            O => \N__10518\,
            I => \transmit_module.video_signal_controller.n3486\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__10515\,
            I => \transmit_module.video_signal_controller.n3486\
        );

    \I__1341\ : InMux
    port map (
            O => \N__10510\,
            I => \N__10507\
        );

    \I__1340\ : LocalMux
    port map (
            O => \N__10507\,
            I => \N__10504\
        );

    \I__1339\ : Span4Mux_h
    port map (
            O => \N__10504\,
            I => \N__10501\
        );

    \I__1338\ : Odrv4
    port map (
            O => \N__10501\,
            I => \transmit_module.video_signal_controller.n7\
        );

    \I__1337\ : CascadeMux
    port map (
            O => \N__10498\,
            I => \N__10495\
        );

    \I__1336\ : InMux
    port map (
            O => \N__10495\,
            I => \N__10492\
        );

    \I__1335\ : LocalMux
    port map (
            O => \N__10492\,
            I => \N__10486\
        );

    \I__1334\ : InMux
    port map (
            O => \N__10491\,
            I => \N__10480\
        );

    \I__1333\ : InMux
    port map (
            O => \N__10490\,
            I => \N__10480\
        );

    \I__1332\ : InMux
    port map (
            O => \N__10489\,
            I => \N__10477\
        );

    \I__1331\ : Span4Mux_h
    port map (
            O => \N__10486\,
            I => \N__10474\
        );

    \I__1330\ : InMux
    port map (
            O => \N__10485\,
            I => \N__10471\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__10480\,
            I => \N__10468\
        );

    \I__1328\ : LocalMux
    port map (
            O => \N__10477\,
            I => \transmit_module.video_signal_controller.VGA_X_11\
        );

    \I__1327\ : Odrv4
    port map (
            O => \N__10474\,
            I => \transmit_module.video_signal_controller.VGA_X_11\
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__10471\,
            I => \transmit_module.video_signal_controller.VGA_X_11\
        );

    \I__1325\ : Odrv4
    port map (
            O => \N__10468\,
            I => \transmit_module.video_signal_controller.VGA_X_11\
        );

    \I__1324\ : InMux
    port map (
            O => \N__10459\,
            I => \N__10456\
        );

    \I__1323\ : LocalMux
    port map (
            O => \N__10456\,
            I => \N__10452\
        );

    \I__1322\ : InMux
    port map (
            O => \N__10455\,
            I => \N__10449\
        );

    \I__1321\ : Odrv4
    port map (
            O => \N__10452\,
            I => \transmit_module.video_signal_controller.VGA_VISIBLE_N_578\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__10449\,
            I => \transmit_module.video_signal_controller.VGA_VISIBLE_N_578\
        );

    \I__1319\ : CascadeMux
    port map (
            O => \N__10444\,
            I => \transmit_module.n111_cascade_\
        );

    \I__1318\ : CascadeMux
    port map (
            O => \N__10441\,
            I => \N__10438\
        );

    \I__1317\ : CascadeBuf
    port map (
            O => \N__10438\,
            I => \N__10435\
        );

    \I__1316\ : CascadeMux
    port map (
            O => \N__10435\,
            I => \N__10432\
        );

    \I__1315\ : CascadeBuf
    port map (
            O => \N__10432\,
            I => \N__10428\
        );

    \I__1314\ : CascadeMux
    port map (
            O => \N__10431\,
            I => \N__10425\
        );

    \I__1313\ : CascadeMux
    port map (
            O => \N__10428\,
            I => \N__10422\
        );

    \I__1312\ : CascadeBuf
    port map (
            O => \N__10425\,
            I => \N__10419\
        );

    \I__1311\ : CascadeBuf
    port map (
            O => \N__10422\,
            I => \N__10416\
        );

    \I__1310\ : CascadeMux
    port map (
            O => \N__10419\,
            I => \N__10413\
        );

    \I__1309\ : CascadeMux
    port map (
            O => \N__10416\,
            I => \N__10410\
        );

    \I__1308\ : CascadeBuf
    port map (
            O => \N__10413\,
            I => \N__10407\
        );

    \I__1307\ : CascadeBuf
    port map (
            O => \N__10410\,
            I => \N__10404\
        );

    \I__1306\ : CascadeMux
    port map (
            O => \N__10407\,
            I => \N__10401\
        );

    \I__1305\ : CascadeMux
    port map (
            O => \N__10404\,
            I => \N__10398\
        );

    \I__1304\ : CascadeBuf
    port map (
            O => \N__10401\,
            I => \N__10395\
        );

    \I__1303\ : CascadeBuf
    port map (
            O => \N__10398\,
            I => \N__10392\
        );

    \I__1302\ : CascadeMux
    port map (
            O => \N__10395\,
            I => \N__10389\
        );

    \I__1301\ : CascadeMux
    port map (
            O => \N__10392\,
            I => \N__10386\
        );

    \I__1300\ : CascadeBuf
    port map (
            O => \N__10389\,
            I => \N__10383\
        );

    \I__1299\ : CascadeBuf
    port map (
            O => \N__10386\,
            I => \N__10380\
        );

    \I__1298\ : CascadeMux
    port map (
            O => \N__10383\,
            I => \N__10377\
        );

    \I__1297\ : CascadeMux
    port map (
            O => \N__10380\,
            I => \N__10374\
        );

    \I__1296\ : CascadeBuf
    port map (
            O => \N__10377\,
            I => \N__10371\
        );

    \I__1295\ : CascadeBuf
    port map (
            O => \N__10374\,
            I => \N__10368\
        );

    \I__1294\ : CascadeMux
    port map (
            O => \N__10371\,
            I => \N__10365\
        );

    \I__1293\ : CascadeMux
    port map (
            O => \N__10368\,
            I => \N__10362\
        );

    \I__1292\ : CascadeBuf
    port map (
            O => \N__10365\,
            I => \N__10359\
        );

    \I__1291\ : CascadeBuf
    port map (
            O => \N__10362\,
            I => \N__10356\
        );

    \I__1290\ : CascadeMux
    port map (
            O => \N__10359\,
            I => \N__10353\
        );

    \I__1289\ : CascadeMux
    port map (
            O => \N__10356\,
            I => \N__10350\
        );

    \I__1288\ : CascadeBuf
    port map (
            O => \N__10353\,
            I => \N__10347\
        );

    \I__1287\ : CascadeBuf
    port map (
            O => \N__10350\,
            I => \N__10344\
        );

    \I__1286\ : CascadeMux
    port map (
            O => \N__10347\,
            I => \N__10341\
        );

    \I__1285\ : CascadeMux
    port map (
            O => \N__10344\,
            I => \N__10338\
        );

    \I__1284\ : CascadeBuf
    port map (
            O => \N__10341\,
            I => \N__10335\
        );

    \I__1283\ : CascadeBuf
    port map (
            O => \N__10338\,
            I => \N__10332\
        );

    \I__1282\ : CascadeMux
    port map (
            O => \N__10335\,
            I => \N__10329\
        );

    \I__1281\ : CascadeMux
    port map (
            O => \N__10332\,
            I => \N__10326\
        );

    \I__1280\ : CascadeBuf
    port map (
            O => \N__10329\,
            I => \N__10323\
        );

    \I__1279\ : CascadeBuf
    port map (
            O => \N__10326\,
            I => \N__10320\
        );

    \I__1278\ : CascadeMux
    port map (
            O => \N__10323\,
            I => \N__10317\
        );

    \I__1277\ : CascadeMux
    port map (
            O => \N__10320\,
            I => \N__10314\
        );

    \I__1276\ : CascadeBuf
    port map (
            O => \N__10317\,
            I => \N__10311\
        );

    \I__1275\ : CascadeBuf
    port map (
            O => \N__10314\,
            I => \N__10308\
        );

    \I__1274\ : CascadeMux
    port map (
            O => \N__10311\,
            I => \N__10305\
        );

    \I__1273\ : CascadeMux
    port map (
            O => \N__10308\,
            I => \N__10302\
        );

    \I__1272\ : CascadeBuf
    port map (
            O => \N__10305\,
            I => \N__10299\
        );

    \I__1271\ : CascadeBuf
    port map (
            O => \N__10302\,
            I => \N__10296\
        );

    \I__1270\ : CascadeMux
    port map (
            O => \N__10299\,
            I => \N__10293\
        );

    \I__1269\ : CascadeMux
    port map (
            O => \N__10296\,
            I => \N__10290\
        );

    \I__1268\ : CascadeBuf
    port map (
            O => \N__10293\,
            I => \N__10287\
        );

    \I__1267\ : CascadeBuf
    port map (
            O => \N__10290\,
            I => \N__10284\
        );

    \I__1266\ : CascadeMux
    port map (
            O => \N__10287\,
            I => \N__10281\
        );

    \I__1265\ : CascadeMux
    port map (
            O => \N__10284\,
            I => \N__10278\
        );

    \I__1264\ : CascadeBuf
    port map (
            O => \N__10281\,
            I => \N__10275\
        );

    \I__1263\ : CascadeBuf
    port map (
            O => \N__10278\,
            I => \N__10272\
        );

    \I__1262\ : CascadeMux
    port map (
            O => \N__10275\,
            I => \N__10269\
        );

    \I__1261\ : CascadeMux
    port map (
            O => \N__10272\,
            I => \N__10266\
        );

    \I__1260\ : CascadeBuf
    port map (
            O => \N__10269\,
            I => \N__10263\
        );

    \I__1259\ : InMux
    port map (
            O => \N__10266\,
            I => \N__10260\
        );

    \I__1258\ : CascadeMux
    port map (
            O => \N__10263\,
            I => \N__10257\
        );

    \I__1257\ : LocalMux
    port map (
            O => \N__10260\,
            I => \N__10254\
        );

    \I__1256\ : CascadeBuf
    port map (
            O => \N__10257\,
            I => \N__10251\
        );

    \I__1255\ : Span4Mux_v
    port map (
            O => \N__10254\,
            I => \N__10248\
        );

    \I__1254\ : CascadeMux
    port map (
            O => \N__10251\,
            I => \N__10245\
        );

    \I__1253\ : Span4Mux_v
    port map (
            O => \N__10248\,
            I => \N__10242\
        );

    \I__1252\ : InMux
    port map (
            O => \N__10245\,
            I => \N__10239\
        );

    \I__1251\ : Span4Mux_v
    port map (
            O => \N__10242\,
            I => \N__10236\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__10239\,
            I => \N__10233\
        );

    \I__1249\ : Span4Mux_h
    port map (
            O => \N__10236\,
            I => \N__10230\
        );

    \I__1248\ : Span4Mux_v
    port map (
            O => \N__10233\,
            I => \N__10227\
        );

    \I__1247\ : Span4Mux_h
    port map (
            O => \N__10230\,
            I => \N__10224\
        );

    \I__1246\ : Span4Mux_v
    port map (
            O => \N__10227\,
            I => \N__10221\
        );

    \I__1245\ : Span4Mux_h
    port map (
            O => \N__10224\,
            I => \N__10216\
        );

    \I__1244\ : Span4Mux_h
    port map (
            O => \N__10221\,
            I => \N__10216\
        );

    \I__1243\ : Sp12to4
    port map (
            O => \N__10216\,
            I => \N__10213\
        );

    \I__1242\ : Odrv12
    port map (
            O => \N__10213\,
            I => n23
        );

    \I__1241\ : InMux
    port map (
            O => \N__10210\,
            I => \N__10207\
        );

    \I__1240\ : LocalMux
    port map (
            O => \N__10207\,
            I => \transmit_module.video_signal_controller.n8\
        );

    \I__1239\ : CascadeMux
    port map (
            O => \N__10204\,
            I => \transmit_module.video_signal_controller.n7_adj_615_cascade_\
        );

    \I__1238\ : CascadeMux
    port map (
            O => \N__10201\,
            I => \transmit_module.video_signal_controller.n2_cascade_\
        );

    \I__1237\ : InMux
    port map (
            O => \N__10198\,
            I => \N__10195\
        );

    \I__1236\ : LocalMux
    port map (
            O => \N__10195\,
            I => \transmit_module.video_signal_controller.n3785\
        );

    \I__1235\ : CascadeMux
    port map (
            O => \N__10192\,
            I => \transmit_module.video_signal_controller.n3577_cascade_\
        );

    \I__1234\ : InMux
    port map (
            O => \N__10189\,
            I => \N__10183\
        );

    \I__1233\ : InMux
    port map (
            O => \N__10188\,
            I => \N__10183\
        );

    \I__1232\ : LocalMux
    port map (
            O => \N__10183\,
            I => \transmit_module.video_signal_controller.n3485\
        );

    \I__1231\ : InMux
    port map (
            O => \N__10180\,
            I => \N__10172\
        );

    \I__1230\ : InMux
    port map (
            O => \N__10179\,
            I => \N__10172\
        );

    \I__1229\ : InMux
    port map (
            O => \N__10178\,
            I => \N__10169\
        );

    \I__1228\ : InMux
    port map (
            O => \N__10177\,
            I => \N__10166\
        );

    \I__1227\ : LocalMux
    port map (
            O => \N__10172\,
            I => \N__10163\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__10169\,
            I => \transmit_module.video_signal_controller.VGA_Y_9\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__10166\,
            I => \transmit_module.video_signal_controller.VGA_Y_9\
        );

    \I__1224\ : Odrv4
    port map (
            O => \N__10163\,
            I => \transmit_module.video_signal_controller.VGA_Y_9\
        );

    \I__1223\ : InMux
    port map (
            O => \N__10156\,
            I => \N__10150\
        );

    \I__1222\ : InMux
    port map (
            O => \N__10155\,
            I => \N__10147\
        );

    \I__1221\ : InMux
    port map (
            O => \N__10154\,
            I => \N__10142\
        );

    \I__1220\ : InMux
    port map (
            O => \N__10153\,
            I => \N__10142\
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__10150\,
            I => \transmit_module.video_signal_controller.VGA_Y_6\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__10147\,
            I => \transmit_module.video_signal_controller.VGA_Y_6\
        );

    \I__1217\ : LocalMux
    port map (
            O => \N__10142\,
            I => \transmit_module.video_signal_controller.VGA_Y_6\
        );

    \I__1216\ : InMux
    port map (
            O => \N__10135\,
            I => \N__10130\
        );

    \I__1215\ : InMux
    port map (
            O => \N__10134\,
            I => \N__10125\
        );

    \I__1214\ : InMux
    port map (
            O => \N__10133\,
            I => \N__10125\
        );

    \I__1213\ : LocalMux
    port map (
            O => \N__10130\,
            I => \transmit_module.video_signal_controller.VGA_Y_11\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__10125\,
            I => \transmit_module.video_signal_controller.VGA_Y_11\
        );

    \I__1211\ : InMux
    port map (
            O => \N__10120\,
            I => \N__10114\
        );

    \I__1210\ : InMux
    port map (
            O => \N__10119\,
            I => \N__10111\
        );

    \I__1209\ : InMux
    port map (
            O => \N__10118\,
            I => \N__10106\
        );

    \I__1208\ : InMux
    port map (
            O => \N__10117\,
            I => \N__10106\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__10114\,
            I => \transmit_module.video_signal_controller.VGA_Y_7\
        );

    \I__1206\ : LocalMux
    port map (
            O => \N__10111\,
            I => \transmit_module.video_signal_controller.VGA_Y_7\
        );

    \I__1205\ : LocalMux
    port map (
            O => \N__10106\,
            I => \transmit_module.video_signal_controller.VGA_Y_7\
        );

    \I__1204\ : CascadeMux
    port map (
            O => \N__10099\,
            I => \N__10096\
        );

    \I__1203\ : InMux
    port map (
            O => \N__10096\,
            I => \N__10090\
        );

    \I__1202\ : InMux
    port map (
            O => \N__10095\,
            I => \N__10087\
        );

    \I__1201\ : InMux
    port map (
            O => \N__10094\,
            I => \N__10082\
        );

    \I__1200\ : InMux
    port map (
            O => \N__10093\,
            I => \N__10082\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__10090\,
            I => \transmit_module.video_signal_controller.VGA_Y_5\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__10087\,
            I => \transmit_module.video_signal_controller.VGA_Y_5\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__10082\,
            I => \transmit_module.video_signal_controller.VGA_Y_5\
        );

    \I__1196\ : InMux
    port map (
            O => \N__10075\,
            I => \N__10069\
        );

    \I__1195\ : InMux
    port map (
            O => \N__10074\,
            I => \N__10066\
        );

    \I__1194\ : InMux
    port map (
            O => \N__10073\,
            I => \N__10061\
        );

    \I__1193\ : InMux
    port map (
            O => \N__10072\,
            I => \N__10061\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__10069\,
            I => \transmit_module.video_signal_controller.VGA_Y_2\
        );

    \I__1191\ : LocalMux
    port map (
            O => \N__10066\,
            I => \transmit_module.video_signal_controller.VGA_Y_2\
        );

    \I__1190\ : LocalMux
    port map (
            O => \N__10061\,
            I => \transmit_module.video_signal_controller.VGA_Y_2\
        );

    \I__1189\ : CEMux
    port map (
            O => \N__10054\,
            I => \N__10046\
        );

    \I__1188\ : CEMux
    port map (
            O => \N__10053\,
            I => \N__10043\
        );

    \I__1187\ : CEMux
    port map (
            O => \N__10052\,
            I => \N__10040\
        );

    \I__1186\ : CEMux
    port map (
            O => \N__10051\,
            I => \N__10036\
        );

    \I__1185\ : CEMux
    port map (
            O => \N__10050\,
            I => \N__10032\
        );

    \I__1184\ : CEMux
    port map (
            O => \N__10049\,
            I => \N__10029\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__10046\,
            I => \N__10025\
        );

    \I__1182\ : LocalMux
    port map (
            O => \N__10043\,
            I => \N__10021\
        );

    \I__1181\ : LocalMux
    port map (
            O => \N__10040\,
            I => \N__10018\
        );

    \I__1180\ : CEMux
    port map (
            O => \N__10039\,
            I => \N__10015\
        );

    \I__1179\ : LocalMux
    port map (
            O => \N__10036\,
            I => \N__10012\
        );

    \I__1178\ : CEMux
    port map (
            O => \N__10035\,
            I => \N__10009\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__10032\,
            I => \N__10006\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__10029\,
            I => \N__10003\
        );

    \I__1175\ : CEMux
    port map (
            O => \N__10028\,
            I => \N__10000\
        );

    \I__1174\ : Span4Mux_h
    port map (
            O => \N__10025\,
            I => \N__9997\
        );

    \I__1173\ : CEMux
    port map (
            O => \N__10024\,
            I => \N__9994\
        );

    \I__1172\ : Span4Mux_v
    port map (
            O => \N__10021\,
            I => \N__9989\
        );

    \I__1171\ : Span4Mux_v
    port map (
            O => \N__10018\,
            I => \N__9989\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__10015\,
            I => \N__9986\
        );

    \I__1169\ : Span4Mux_v
    port map (
            O => \N__10012\,
            I => \N__9981\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__10009\,
            I => \N__9981\
        );

    \I__1167\ : Span4Mux_v
    port map (
            O => \N__10006\,
            I => \N__9976\
        );

    \I__1166\ : Span4Mux_h
    port map (
            O => \N__10003\,
            I => \N__9976\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__10000\,
            I => \N__9973\
        );

    \I__1164\ : Span4Mux_h
    port map (
            O => \N__9997\,
            I => \N__9968\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__9994\,
            I => \N__9968\
        );

    \I__1162\ : Span4Mux_v
    port map (
            O => \N__9989\,
            I => \N__9965\
        );

    \I__1161\ : Span12Mux_h
    port map (
            O => \N__9986\,
            I => \N__9962\
        );

    \I__1160\ : Span4Mux_h
    port map (
            O => \N__9981\,
            I => \N__9959\
        );

    \I__1159\ : Span4Mux_h
    port map (
            O => \N__9976\,
            I => \N__9954\
        );

    \I__1158\ : Span4Mux_h
    port map (
            O => \N__9973\,
            I => \N__9954\
        );

    \I__1157\ : Span4Mux_h
    port map (
            O => \N__9968\,
            I => \N__9951\
        );

    \I__1156\ : Odrv4
    port map (
            O => \N__9965\,
            I => \transmit_module.n3798\
        );

    \I__1155\ : Odrv12
    port map (
            O => \N__9962\,
            I => \transmit_module.n3798\
        );

    \I__1154\ : Odrv4
    port map (
            O => \N__9959\,
            I => \transmit_module.n3798\
        );

    \I__1153\ : Odrv4
    port map (
            O => \N__9954\,
            I => \transmit_module.n3798\
        );

    \I__1152\ : Odrv4
    port map (
            O => \N__9951\,
            I => \transmit_module.n3798\
        );

    \I__1151\ : InMux
    port map (
            O => \N__9940\,
            I => \receive_module.rx_counter.n3275\
        );

    \I__1150\ : InMux
    port map (
            O => \N__9937\,
            I => \receive_module.rx_counter.n3276\
        );

    \I__1149\ : InMux
    port map (
            O => \N__9934\,
            I => \receive_module.rx_counter.n3277\
        );

    \I__1148\ : InMux
    port map (
            O => \N__9931\,
            I => \bfn_13_11_0_\
        );

    \I__1147\ : CascadeMux
    port map (
            O => \N__9928\,
            I => \transmit_module.video_signal_controller.n3786_cascade_\
        );

    \I__1146\ : InMux
    port map (
            O => \N__9925\,
            I => \N__9922\
        );

    \I__1145\ : LocalMux
    port map (
            O => \N__9922\,
            I => \transmit_module.Y_DELTA_PATTERN_4\
        );

    \I__1144\ : InMux
    port map (
            O => \N__9919\,
            I => \N__9916\
        );

    \I__1143\ : LocalMux
    port map (
            O => \N__9916\,
            I => \transmit_module.Y_DELTA_PATTERN_3\
        );

    \I__1142\ : InMux
    port map (
            O => \N__9913\,
            I => \N__9910\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__9910\,
            I => \N__9907\
        );

    \I__1140\ : Span12Mux_v
    port map (
            O => \N__9907\,
            I => \N__9904\
        );

    \I__1139\ : Odrv12
    port map (
            O => \N__9904\,
            I => \line_buffer.n578\
        );

    \I__1138\ : InMux
    port map (
            O => \N__9901\,
            I => \N__9898\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__9898\,
            I => \N__9895\
        );

    \I__1136\ : Span4Mux_h
    port map (
            O => \N__9895\,
            I => \N__9892\
        );

    \I__1135\ : Odrv4
    port map (
            O => \N__9892\,
            I => \line_buffer.n570\
        );

    \I__1134\ : InMux
    port map (
            O => \N__9889\,
            I => \N__9886\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__9886\,
            I => \N__9883\
        );

    \I__1132\ : Span12Mux_v
    port map (
            O => \N__9883\,
            I => \N__9880\
        );

    \I__1131\ : Odrv12
    port map (
            O => \N__9880\,
            I => \line_buffer.n577\
        );

    \I__1130\ : InMux
    port map (
            O => \N__9877\,
            I => \N__9874\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__9874\,
            I => \N__9871\
        );

    \I__1128\ : Span12Mux_v
    port map (
            O => \N__9871\,
            I => \N__9868\
        );

    \I__1127\ : Odrv12
    port map (
            O => \N__9868\,
            I => \line_buffer.n569\
        );

    \I__1126\ : InMux
    port map (
            O => \N__9865\,
            I => \bfn_13_10_0_\
        );

    \I__1125\ : InMux
    port map (
            O => \N__9862\,
            I => \receive_module.rx_counter.n3271\
        );

    \I__1124\ : InMux
    port map (
            O => \N__9859\,
            I => \receive_module.rx_counter.n3272\
        );

    \I__1123\ : InMux
    port map (
            O => \N__9856\,
            I => \receive_module.rx_counter.n3273\
        );

    \I__1122\ : InMux
    port map (
            O => \N__9853\,
            I => \receive_module.rx_counter.n3274\
        );

    \I__1121\ : SRMux
    port map (
            O => \N__9850\,
            I => \N__9846\
        );

    \I__1120\ : SRMux
    port map (
            O => \N__9849\,
            I => \N__9843\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__9846\,
            I => \transmit_module.video_signal_controller.n2361\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__9843\,
            I => \transmit_module.video_signal_controller.n2361\
        );

    \I__1117\ : CascadeMux
    port map (
            O => \N__9838\,
            I => \transmit_module.n3787_cascade_\
        );

    \I__1116\ : InMux
    port map (
            O => \N__9835\,
            I => \N__9832\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__9832\,
            I => \transmit_module.Y_DELTA_PATTERN_7\
        );

    \I__1114\ : InMux
    port map (
            O => \N__9829\,
            I => \N__9826\
        );

    \I__1113\ : LocalMux
    port map (
            O => \N__9826\,
            I => \transmit_module.Y_DELTA_PATTERN_6\
        );

    \I__1112\ : InMux
    port map (
            O => \N__9823\,
            I => \N__9820\
        );

    \I__1111\ : LocalMux
    port map (
            O => \N__9820\,
            I => \transmit_module.Y_DELTA_PATTERN_5\
        );

    \I__1110\ : InMux
    port map (
            O => \N__9817\,
            I => \transmit_module.video_signal_controller.n3292\
        );

    \I__1109\ : InMux
    port map (
            O => \N__9814\,
            I => \transmit_module.video_signal_controller.n3293\
        );

    \I__1108\ : InMux
    port map (
            O => \N__9811\,
            I => \transmit_module.video_signal_controller.n3294\
        );

    \I__1107\ : InMux
    port map (
            O => \N__9808\,
            I => \transmit_module.video_signal_controller.n3295\
        );

    \I__1106\ : InMux
    port map (
            O => \N__9805\,
            I => \transmit_module.video_signal_controller.n3296\
        );

    \I__1105\ : InMux
    port map (
            O => \N__9802\,
            I => \bfn_12_14_0_\
        );

    \I__1104\ : InMux
    port map (
            O => \N__9799\,
            I => \transmit_module.video_signal_controller.n3298\
        );

    \I__1103\ : InMux
    port map (
            O => \N__9796\,
            I => \transmit_module.video_signal_controller.n3299\
        );

    \I__1102\ : InMux
    port map (
            O => \N__9793\,
            I => \transmit_module.video_signal_controller.n3300\
        );

    \I__1101\ : SRMux
    port map (
            O => \N__9790\,
            I => \N__9787\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__9787\,
            I => \N__9783\
        );

    \I__1099\ : SRMux
    port map (
            O => \N__9786\,
            I => \N__9779\
        );

    \I__1098\ : Span4Mux_v
    port map (
            O => \N__9783\,
            I => \N__9775\
        );

    \I__1097\ : CEMux
    port map (
            O => \N__9782\,
            I => \N__9772\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__9779\,
            I => \N__9769\
        );

    \I__1095\ : CEMux
    port map (
            O => \N__9778\,
            I => \N__9766\
        );

    \I__1094\ : Span4Mux_h
    port map (
            O => \N__9775\,
            I => \N__9759\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__9772\,
            I => \N__9759\
        );

    \I__1092\ : Span4Mux_v
    port map (
            O => \N__9769\,
            I => \N__9759\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__9766\,
            I => \transmit_module.video_signal_controller.n2010\
        );

    \I__1090\ : Odrv4
    port map (
            O => \N__9759\,
            I => \transmit_module.video_signal_controller.n2010\
        );

    \I__1089\ : InMux
    port map (
            O => \N__9754\,
            I => \N__9751\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__9751\,
            I => \transmit_module.Y_DELTA_PATTERN_60\
        );

    \I__1087\ : InMux
    port map (
            O => \N__9748\,
            I => \N__9745\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__9745\,
            I => \transmit_module.Y_DELTA_PATTERN_59\
        );

    \I__1085\ : InMux
    port map (
            O => \N__9742\,
            I => \N__9739\
        );

    \I__1084\ : LocalMux
    port map (
            O => \N__9739\,
            I => \transmit_module.Y_DELTA_PATTERN_98\
        );

    \I__1083\ : InMux
    port map (
            O => \N__9736\,
            I => \N__9733\
        );

    \I__1082\ : LocalMux
    port map (
            O => \N__9733\,
            I => \N__9730\
        );

    \I__1081\ : Odrv4
    port map (
            O => \N__9730\,
            I => \transmit_module.Y_DELTA_PATTERN_86\
        );

    \I__1080\ : InMux
    port map (
            O => \N__9727\,
            I => \N__9724\
        );

    \I__1079\ : LocalMux
    port map (
            O => \N__9724\,
            I => \transmit_module.Y_DELTA_PATTERN_85\
        );

    \I__1078\ : InMux
    port map (
            O => \N__9721\,
            I => \N__9718\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__9718\,
            I => \transmit_module.Y_DELTA_PATTERN_84\
        );

    \I__1076\ : InMux
    port map (
            O => \N__9715\,
            I => \N__9712\
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__9712\,
            I => \transmit_module.Y_DELTA_PATTERN_83\
        );

    \I__1074\ : InMux
    port map (
            O => \N__9709\,
            I => \N__9706\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__9706\,
            I => \transmit_module.Y_DELTA_PATTERN_99\
        );

    \I__1072\ : InMux
    port map (
            O => \N__9703\,
            I => \bfn_12_13_0_\
        );

    \I__1071\ : InMux
    port map (
            O => \N__9700\,
            I => \transmit_module.video_signal_controller.n3290\
        );

    \I__1070\ : InMux
    port map (
            O => \N__9697\,
            I => \transmit_module.video_signal_controller.n3291\
        );

    \I__1069\ : CascadeMux
    port map (
            O => \N__9694\,
            I => \N__9691\
        );

    \I__1068\ : InMux
    port map (
            O => \N__9691\,
            I => \N__9683\
        );

    \I__1067\ : InMux
    port map (
            O => \N__9690\,
            I => \N__9683\
        );

    \I__1066\ : InMux
    port map (
            O => \N__9689\,
            I => \N__9680\
        );

    \I__1065\ : InMux
    port map (
            O => \N__9688\,
            I => \N__9677\
        );

    \I__1064\ : LocalMux
    port map (
            O => \N__9683\,
            I => \N__9674\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__9680\,
            I => \transmit_module.video_signal_controller.VGA_X_8\
        );

    \I__1062\ : LocalMux
    port map (
            O => \N__9677\,
            I => \transmit_module.video_signal_controller.VGA_X_8\
        );

    \I__1061\ : Odrv4
    port map (
            O => \N__9674\,
            I => \transmit_module.video_signal_controller.VGA_X_8\
        );

    \I__1060\ : CascadeMux
    port map (
            O => \N__9667\,
            I => \transmit_module.video_signal_controller.n4_adj_617_cascade_\
        );

    \I__1059\ : InMux
    port map (
            O => \N__9664\,
            I => \N__9658\
        );

    \I__1058\ : InMux
    port map (
            O => \N__9663\,
            I => \N__9655\
        );

    \I__1057\ : InMux
    port map (
            O => \N__9662\,
            I => \N__9652\
        );

    \I__1056\ : InMux
    port map (
            O => \N__9661\,
            I => \N__9649\
        );

    \I__1055\ : LocalMux
    port map (
            O => \N__9658\,
            I => \transmit_module.video_signal_controller.VGA_X_6\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__9655\,
            I => \transmit_module.video_signal_controller.VGA_X_6\
        );

    \I__1053\ : LocalMux
    port map (
            O => \N__9652\,
            I => \transmit_module.video_signal_controller.VGA_X_6\
        );

    \I__1052\ : LocalMux
    port map (
            O => \N__9649\,
            I => \transmit_module.video_signal_controller.VGA_X_6\
        );

    \I__1051\ : CascadeMux
    port map (
            O => \N__9640\,
            I => \N__9636\
        );

    \I__1050\ : InMux
    port map (
            O => \N__9639\,
            I => \N__9630\
        );

    \I__1049\ : InMux
    port map (
            O => \N__9636\,
            I => \N__9630\
        );

    \I__1048\ : InMux
    port map (
            O => \N__9635\,
            I => \N__9626\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__9630\,
            I => \N__9623\
        );

    \I__1046\ : InMux
    port map (
            O => \N__9629\,
            I => \N__9620\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__9626\,
            I => \transmit_module.video_signal_controller.VGA_X_9\
        );

    \I__1044\ : Odrv4
    port map (
            O => \N__9623\,
            I => \transmit_module.video_signal_controller.VGA_X_9\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__9620\,
            I => \transmit_module.video_signal_controller.VGA_X_9\
        );

    \I__1042\ : InMux
    port map (
            O => \N__9613\,
            I => \N__9607\
        );

    \I__1041\ : InMux
    port map (
            O => \N__9612\,
            I => \N__9607\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__9607\,
            I => \N__9603\
        );

    \I__1039\ : InMux
    port map (
            O => \N__9606\,
            I => \N__9599\
        );

    \I__1038\ : Span4Mux_v
    port map (
            O => \N__9603\,
            I => \N__9596\
        );

    \I__1037\ : InMux
    port map (
            O => \N__9602\,
            I => \N__9593\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__9599\,
            I => \transmit_module.video_signal_controller.VGA_X_10\
        );

    \I__1035\ : Odrv4
    port map (
            O => \N__9596\,
            I => \transmit_module.video_signal_controller.VGA_X_10\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__9593\,
            I => \transmit_module.video_signal_controller.VGA_X_10\
        );

    \I__1033\ : InMux
    port map (
            O => \N__9586\,
            I => \N__9583\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__9583\,
            I => \transmit_module.video_signal_controller.n4\
        );

    \I__1031\ : CascadeMux
    port map (
            O => \N__9580\,
            I => \N__9577\
        );

    \I__1030\ : InMux
    port map (
            O => \N__9577\,
            I => \N__9569\
        );

    \I__1029\ : InMux
    port map (
            O => \N__9576\,
            I => \N__9569\
        );

    \I__1028\ : InMux
    port map (
            O => \N__9575\,
            I => \N__9566\
        );

    \I__1027\ : InMux
    port map (
            O => \N__9574\,
            I => \N__9563\
        );

    \I__1026\ : LocalMux
    port map (
            O => \N__9569\,
            I => \transmit_module.video_signal_controller.VGA_X_7\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__9566\,
            I => \transmit_module.video_signal_controller.VGA_X_7\
        );

    \I__1024\ : LocalMux
    port map (
            O => \N__9563\,
            I => \transmit_module.video_signal_controller.VGA_X_7\
        );

    \I__1023\ : CascadeMux
    port map (
            O => \N__9556\,
            I => \transmit_module.video_signal_controller.n3794_cascade_\
        );

    \I__1022\ : InMux
    port map (
            O => \N__9553\,
            I => \N__9545\
        );

    \I__1021\ : InMux
    port map (
            O => \N__9552\,
            I => \N__9545\
        );

    \I__1020\ : InMux
    port map (
            O => \N__9551\,
            I => \N__9542\
        );

    \I__1019\ : InMux
    port map (
            O => \N__9550\,
            I => \N__9539\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__9545\,
            I => \transmit_module.video_signal_controller.VGA_X_4\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__9542\,
            I => \transmit_module.video_signal_controller.VGA_X_4\
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__9539\,
            I => \transmit_module.video_signal_controller.VGA_X_4\
        );

    \I__1015\ : InMux
    port map (
            O => \N__9532\,
            I => \N__9529\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__9529\,
            I => \transmit_module.video_signal_controller.n3618\
        );

    \I__1013\ : InMux
    port map (
            O => \N__9526\,
            I => \N__9523\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__9523\,
            I => \transmit_module.Y_DELTA_PATTERN_61\
        );

    \I__1011\ : InMux
    port map (
            O => \N__9520\,
            I => \N__9517\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__9517\,
            I => \transmit_module.Y_DELTA_PATTERN_37\
        );

    \I__1009\ : InMux
    port map (
            O => \N__9514\,
            I => \N__9511\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__9511\,
            I => \transmit_module.Y_DELTA_PATTERN_39\
        );

    \I__1007\ : InMux
    port map (
            O => \N__9508\,
            I => \N__9505\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__9505\,
            I => \transmit_module.Y_DELTA_PATTERN_38\
        );

    \I__1005\ : InMux
    port map (
            O => \N__9502\,
            I => \N__9499\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__9499\,
            I => \transmit_module.Y_DELTA_PATTERN_58\
        );

    \I__1003\ : InMux
    port map (
            O => \N__9496\,
            I => \N__9493\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__9493\,
            I => \transmit_module.Y_DELTA_PATTERN_57\
        );

    \I__1001\ : InMux
    port map (
            O => \N__9490\,
            I => \N__9487\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__9487\,
            I => \transmit_module.Y_DELTA_PATTERN_71\
        );

    \I__999\ : InMux
    port map (
            O => \N__9484\,
            I => \N__9481\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__9481\,
            I => \transmit_module.Y_DELTA_PATTERN_70\
        );

    \I__997\ : InMux
    port map (
            O => \N__9478\,
            I => \N__9475\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__9475\,
            I => \transmit_module.Y_DELTA_PATTERN_68\
        );

    \I__995\ : InMux
    port map (
            O => \N__9472\,
            I => \N__9469\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__9469\,
            I => \N__9466\
        );

    \I__993\ : Odrv4
    port map (
            O => \N__9466\,
            I => \transmit_module.Y_DELTA_PATTERN_67\
        );

    \I__992\ : InMux
    port map (
            O => \N__9463\,
            I => \N__9460\
        );

    \I__991\ : LocalMux
    port map (
            O => \N__9460\,
            I => \transmit_module.video_signal_controller.n2886\
        );

    \I__990\ : CascadeMux
    port map (
            O => \N__9457\,
            I => \transmit_module.video_signal_controller.n1983_cascade_\
        );

    \I__989\ : InMux
    port map (
            O => \N__9454\,
            I => \N__9451\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__9451\,
            I => \transmit_module.video_signal_controller.n2926\
        );

    \I__987\ : CascadeMux
    port map (
            O => \N__9448\,
            I => \transmit_module.video_signal_controller.n2010_cascade_\
        );

    \I__986\ : InMux
    port map (
            O => \N__9445\,
            I => \N__9442\
        );

    \I__985\ : LocalMux
    port map (
            O => \N__9442\,
            I => \transmit_module.video_signal_controller.n1983\
        );

    \I__984\ : InMux
    port map (
            O => \N__9439\,
            I => \N__9436\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__9436\,
            I => \transmit_module.video_signal_controller.n3789\
        );

    \I__982\ : InMux
    port map (
            O => \N__9433\,
            I => \N__9427\
        );

    \I__981\ : InMux
    port map (
            O => \N__9432\,
            I => \N__9427\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__9427\,
            I => \transmit_module.video_signal_controller.n3467\
        );

    \I__979\ : CascadeMux
    port map (
            O => \N__9424\,
            I => \transmit_module.video_signal_controller.n18_cascade_\
        );

    \I__978\ : InMux
    port map (
            O => \N__9421\,
            I => \N__9416\
        );

    \I__977\ : InMux
    port map (
            O => \N__9420\,
            I => \N__9412\
        );

    \I__976\ : InMux
    port map (
            O => \N__9419\,
            I => \N__9409\
        );

    \I__975\ : LocalMux
    port map (
            O => \N__9416\,
            I => \N__9406\
        );

    \I__974\ : InMux
    port map (
            O => \N__9415\,
            I => \N__9403\
        );

    \I__973\ : LocalMux
    port map (
            O => \N__9412\,
            I => \transmit_module.video_signal_controller.VGA_X_3\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__9409\,
            I => \transmit_module.video_signal_controller.VGA_X_3\
        );

    \I__971\ : Odrv4
    port map (
            O => \N__9406\,
            I => \transmit_module.video_signal_controller.VGA_X_3\
        );

    \I__970\ : LocalMux
    port map (
            O => \N__9403\,
            I => \transmit_module.video_signal_controller.VGA_X_3\
        );

    \I__969\ : InMux
    port map (
            O => \N__9394\,
            I => \N__9388\
        );

    \I__968\ : InMux
    port map (
            O => \N__9393\,
            I => \N__9385\
        );

    \I__967\ : InMux
    port map (
            O => \N__9392\,
            I => \N__9382\
        );

    \I__966\ : InMux
    port map (
            O => \N__9391\,
            I => \N__9379\
        );

    \I__965\ : LocalMux
    port map (
            O => \N__9388\,
            I => \transmit_module.video_signal_controller.VGA_X_5\
        );

    \I__964\ : LocalMux
    port map (
            O => \N__9385\,
            I => \transmit_module.video_signal_controller.VGA_X_5\
        );

    \I__963\ : LocalMux
    port map (
            O => \N__9382\,
            I => \transmit_module.video_signal_controller.VGA_X_5\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__9379\,
            I => \transmit_module.video_signal_controller.VGA_X_5\
        );

    \I__961\ : InMux
    port map (
            O => \N__9370\,
            I => \N__9367\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__9367\,
            I => \transmit_module.Y_DELTA_PATTERN_81\
        );

    \I__959\ : InMux
    port map (
            O => \N__9364\,
            I => \N__9361\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__9361\,
            I => \transmit_module.Y_DELTA_PATTERN_50\
        );

    \I__957\ : InMux
    port map (
            O => \N__9358\,
            I => \N__9355\
        );

    \I__956\ : LocalMux
    port map (
            O => \N__9355\,
            I => \transmit_module.Y_DELTA_PATTERN_49\
        );

    \I__955\ : InMux
    port map (
            O => \N__9352\,
            I => \N__9349\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__9349\,
            I => \N__9346\
        );

    \I__953\ : Odrv4
    port map (
            O => \N__9346\,
            I => \transmit_module.Y_DELTA_PATTERN_35\
        );

    \I__952\ : InMux
    port map (
            O => \N__9343\,
            I => \N__9340\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__9340\,
            I => \transmit_module.Y_DELTA_PATTERN_34\
        );

    \I__950\ : InMux
    port map (
            O => \N__9337\,
            I => \N__9334\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__9334\,
            I => \transmit_module.Y_DELTA_PATTERN_72\
        );

    \I__948\ : InMux
    port map (
            O => \N__9331\,
            I => \N__9328\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__9328\,
            I => \transmit_module.Y_DELTA_PATTERN_82\
        );

    \I__946\ : InMux
    port map (
            O => \N__9325\,
            I => \N__9322\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__9322\,
            I => \transmit_module.Y_DELTA_PATTERN_69\
        );

    \I__944\ : InMux
    port map (
            O => \N__9319\,
            I => \N__9316\
        );

    \I__943\ : LocalMux
    port map (
            O => \N__9316\,
            I => \N__9313\
        );

    \I__942\ : Span4Mux_h
    port map (
            O => \N__9313\,
            I => \N__9310\
        );

    \I__941\ : Odrv4
    port map (
            O => \N__9310\,
            I => \transmit_module.Y_DELTA_PATTERN_78\
        );

    \I__940\ : InMux
    port map (
            O => \N__9307\,
            I => \N__9304\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__9304\,
            I => \transmit_module.Y_DELTA_PATTERN_80\
        );

    \I__938\ : InMux
    port map (
            O => \N__9301\,
            I => \N__9298\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__9298\,
            I => \transmit_module.Y_DELTA_PATTERN_79\
        );

    \I__936\ : InMux
    port map (
            O => \N__9295\,
            I => \N__9292\
        );

    \I__935\ : LocalMux
    port map (
            O => \N__9292\,
            I => \transmit_module.Y_DELTA_PATTERN_36\
        );

    \I__934\ : InMux
    port map (
            O => \N__9289\,
            I => \N__9286\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__9286\,
            I => \transmit_module.Y_DELTA_PATTERN_62\
        );

    \I__932\ : InMux
    port map (
            O => \N__9283\,
            I => \N__9280\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__9280\,
            I => \transmit_module.Y_DELTA_PATTERN_66\
        );

    \I__930\ : InMux
    port map (
            O => \N__9277\,
            I => \N__9274\
        );

    \I__929\ : LocalMux
    port map (
            O => \N__9274\,
            I => \N__9271\
        );

    \I__928\ : Odrv12
    port map (
            O => \N__9271\,
            I => \transmit_module.Y_DELTA_PATTERN_53\
        );

    \I__927\ : InMux
    port map (
            O => \N__9268\,
            I => \N__9265\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__9265\,
            I => \transmit_module.Y_DELTA_PATTERN_52\
        );

    \I__925\ : InMux
    port map (
            O => \N__9262\,
            I => \N__9259\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__9259\,
            I => \transmit_module.Y_DELTA_PATTERN_51\
        );

    \I__923\ : InMux
    port map (
            O => \N__9256\,
            I => \bfn_10_16_0_\
        );

    \I__922\ : InMux
    port map (
            O => \N__9253\,
            I => \transmit_module.video_signal_controller.n3287\
        );

    \I__921\ : InMux
    port map (
            O => \N__9250\,
            I => \transmit_module.video_signal_controller.n3288\
        );

    \I__920\ : InMux
    port map (
            O => \N__9247\,
            I => \transmit_module.video_signal_controller.n3289\
        );

    \I__919\ : InMux
    port map (
            O => \N__9244\,
            I => \N__9241\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__9241\,
            I => \transmit_module.Y_DELTA_PATTERN_55\
        );

    \I__917\ : InMux
    port map (
            O => \N__9238\,
            I => \N__9235\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__9235\,
            I => \transmit_module.Y_DELTA_PATTERN_54\
        );

    \I__915\ : InMux
    port map (
            O => \N__9232\,
            I => \N__9229\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__9229\,
            I => \transmit_module.Y_DELTA_PATTERN_40\
        );

    \I__913\ : InMux
    port map (
            O => \N__9226\,
            I => \N__9223\
        );

    \I__912\ : LocalMux
    port map (
            O => \N__9223\,
            I => \transmit_module.Y_DELTA_PATTERN_56\
        );

    \I__911\ : InMux
    port map (
            O => \N__9220\,
            I => \N__9217\
        );

    \I__910\ : LocalMux
    port map (
            O => \N__9217\,
            I => \N__9214\
        );

    \I__909\ : Span4Mux_h
    port map (
            O => \N__9214\,
            I => \N__9211\
        );

    \I__908\ : Odrv4
    port map (
            O => \N__9211\,
            I => \transmit_module.Y_DELTA_PATTERN_97\
        );

    \I__907\ : InMux
    port map (
            O => \N__9208\,
            I => \N__9203\
        );

    \I__906\ : InMux
    port map (
            O => \N__9207\,
            I => \N__9198\
        );

    \I__905\ : InMux
    port map (
            O => \N__9206\,
            I => \N__9198\
        );

    \I__904\ : LocalMux
    port map (
            O => \N__9203\,
            I => \transmit_module.video_signal_controller.VGA_X_0\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__9198\,
            I => \transmit_module.video_signal_controller.VGA_X_0\
        );

    \I__902\ : InMux
    port map (
            O => \N__9193\,
            I => \bfn_10_15_0_\
        );

    \I__901\ : CascadeMux
    port map (
            O => \N__9190\,
            I => \N__9184\
        );

    \I__900\ : InMux
    port map (
            O => \N__9189\,
            I => \N__9181\
        );

    \I__899\ : InMux
    port map (
            O => \N__9188\,
            I => \N__9174\
        );

    \I__898\ : InMux
    port map (
            O => \N__9187\,
            I => \N__9174\
        );

    \I__897\ : InMux
    port map (
            O => \N__9184\,
            I => \N__9174\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__9181\,
            I => \transmit_module.video_signal_controller.VGA_X_1\
        );

    \I__895\ : LocalMux
    port map (
            O => \N__9174\,
            I => \transmit_module.video_signal_controller.VGA_X_1\
        );

    \I__894\ : InMux
    port map (
            O => \N__9169\,
            I => \transmit_module.video_signal_controller.n3279\
        );

    \I__893\ : InMux
    port map (
            O => \N__9166\,
            I => \N__9160\
        );

    \I__892\ : InMux
    port map (
            O => \N__9165\,
            I => \N__9153\
        );

    \I__891\ : InMux
    port map (
            O => \N__9164\,
            I => \N__9153\
        );

    \I__890\ : InMux
    port map (
            O => \N__9163\,
            I => \N__9153\
        );

    \I__889\ : LocalMux
    port map (
            O => \N__9160\,
            I => \transmit_module.video_signal_controller.VGA_X_2\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__9153\,
            I => \transmit_module.video_signal_controller.VGA_X_2\
        );

    \I__887\ : InMux
    port map (
            O => \N__9148\,
            I => \transmit_module.video_signal_controller.n3280\
        );

    \I__886\ : InMux
    port map (
            O => \N__9145\,
            I => \transmit_module.video_signal_controller.n3281\
        );

    \I__885\ : InMux
    port map (
            O => \N__9142\,
            I => \transmit_module.video_signal_controller.n3282\
        );

    \I__884\ : InMux
    port map (
            O => \N__9139\,
            I => \transmit_module.video_signal_controller.n3283\
        );

    \I__883\ : InMux
    port map (
            O => \N__9136\,
            I => \transmit_module.video_signal_controller.n3284\
        );

    \I__882\ : InMux
    port map (
            O => \N__9133\,
            I => \transmit_module.video_signal_controller.n3285\
        );

    \I__881\ : InMux
    port map (
            O => \N__9130\,
            I => \N__9127\
        );

    \I__880\ : LocalMux
    port map (
            O => \N__9127\,
            I => \N__9124\
        );

    \I__879\ : Odrv4
    port map (
            O => \N__9124\,
            I => \transmit_module.Y_DELTA_PATTERN_42\
        );

    \I__878\ : InMux
    port map (
            O => \N__9121\,
            I => \N__9118\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__9118\,
            I => \transmit_module.Y_DELTA_PATTERN_96\
        );

    \I__876\ : InMux
    port map (
            O => \N__9115\,
            I => \N__9112\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__9112\,
            I => \transmit_module.Y_DELTA_PATTERN_45\
        );

    \I__874\ : InMux
    port map (
            O => \N__9109\,
            I => \N__9106\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__9106\,
            I => \transmit_module.Y_DELTA_PATTERN_44\
        );

    \I__872\ : InMux
    port map (
            O => \N__9103\,
            I => \N__9100\
        );

    \I__871\ : LocalMux
    port map (
            O => \N__9100\,
            I => \transmit_module.Y_DELTA_PATTERN_43\
        );

    \I__870\ : CascadeMux
    port map (
            O => \N__9097\,
            I => \transmit_module.video_signal_controller.n3788_cascade_\
        );

    \I__869\ : InMux
    port map (
            O => \N__9094\,
            I => \N__9091\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__9091\,
            I => \transmit_module.video_signal_controller.n2876\
        );

    \I__867\ : InMux
    port map (
            O => \N__9088\,
            I => \N__9085\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__9085\,
            I => \transmit_module.Y_DELTA_PATTERN_63\
        );

    \I__865\ : InMux
    port map (
            O => \N__9082\,
            I => \N__9079\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__9079\,
            I => \transmit_module.Y_DELTA_PATTERN_74\
        );

    \I__863\ : InMux
    port map (
            O => \N__9076\,
            I => \N__9073\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__9073\,
            I => \transmit_module.Y_DELTA_PATTERN_76\
        );

    \I__861\ : InMux
    port map (
            O => \N__9070\,
            I => \N__9067\
        );

    \I__860\ : LocalMux
    port map (
            O => \N__9067\,
            I => \transmit_module.Y_DELTA_PATTERN_75\
        );

    \I__859\ : InMux
    port map (
            O => \N__9064\,
            I => \N__9061\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__9061\,
            I => \transmit_module.Y_DELTA_PATTERN_73\
        );

    \I__857\ : InMux
    port map (
            O => \N__9058\,
            I => \N__9055\
        );

    \I__856\ : LocalMux
    port map (
            O => \N__9055\,
            I => \transmit_module.Y_DELTA_PATTERN_48\
        );

    \I__855\ : InMux
    port map (
            O => \N__9052\,
            I => \N__9049\
        );

    \I__854\ : LocalMux
    port map (
            O => \N__9049\,
            I => \transmit_module.Y_DELTA_PATTERN_47\
        );

    \I__853\ : InMux
    port map (
            O => \N__9046\,
            I => \N__9043\
        );

    \I__852\ : LocalMux
    port map (
            O => \N__9043\,
            I => \transmit_module.Y_DELTA_PATTERN_46\
        );

    \I__851\ : InMux
    port map (
            O => \N__9040\,
            I => \N__9037\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__9037\,
            I => \transmit_module.X_DELTA_PATTERN_15\
        );

    \I__849\ : InMux
    port map (
            O => \N__9034\,
            I => \N__9031\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__9031\,
            I => \transmit_module.X_DELTA_PATTERN_12\
        );

    \I__847\ : InMux
    port map (
            O => \N__9028\,
            I => \N__9025\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__9025\,
            I => \transmit_module.X_DELTA_PATTERN_11\
        );

    \I__845\ : InMux
    port map (
            O => \N__9022\,
            I => \N__9019\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__9019\,
            I => \transmit_module.X_DELTA_PATTERN_14\
        );

    \I__843\ : InMux
    port map (
            O => \N__9016\,
            I => \N__9013\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__9013\,
            I => \transmit_module.X_DELTA_PATTERN_13\
        );

    \I__841\ : InMux
    port map (
            O => \N__9010\,
            I => \N__9007\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__9007\,
            I => \transmit_module.Y_DELTA_PATTERN_64\
        );

    \I__839\ : InMux
    port map (
            O => \N__9004\,
            I => \N__9001\
        );

    \I__838\ : LocalMux
    port map (
            O => \N__9001\,
            I => \transmit_module.Y_DELTA_PATTERN_65\
        );

    \I__837\ : InMux
    port map (
            O => \N__8998\,
            I => \N__8995\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__8995\,
            I => \transmit_module.Y_DELTA_PATTERN_41\
        );

    \I__835\ : InMux
    port map (
            O => \N__8992\,
            I => \N__8989\
        );

    \I__834\ : LocalMux
    port map (
            O => \N__8989\,
            I => \transmit_module.Y_DELTA_PATTERN_92\
        );

    \I__833\ : InMux
    port map (
            O => \N__8986\,
            I => \N__8983\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__8983\,
            I => \transmit_module.Y_DELTA_PATTERN_93\
        );

    \I__831\ : InMux
    port map (
            O => \N__8980\,
            I => \N__8977\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__8977\,
            I => \transmit_module.Y_DELTA_PATTERN_95\
        );

    \I__829\ : InMux
    port map (
            O => \N__8974\,
            I => \N__8971\
        );

    \I__828\ : LocalMux
    port map (
            O => \N__8971\,
            I => \transmit_module.Y_DELTA_PATTERN_94\
        );

    \I__827\ : InMux
    port map (
            O => \N__8968\,
            I => \N__8965\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__8965\,
            I => \N__8962\
        );

    \I__825\ : Odrv4
    port map (
            O => \N__8962\,
            I => \transmit_module.X_DELTA_PATTERN_8\
        );

    \I__824\ : InMux
    port map (
            O => \N__8959\,
            I => \N__8956\
        );

    \I__823\ : LocalMux
    port map (
            O => \N__8956\,
            I => \transmit_module.X_DELTA_PATTERN_7\
        );

    \I__822\ : InMux
    port map (
            O => \N__8953\,
            I => \N__8950\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__8950\,
            I => \N__8947\
        );

    \I__820\ : Odrv4
    port map (
            O => \N__8947\,
            I => \transmit_module.X_DELTA_PATTERN_10\
        );

    \I__819\ : InMux
    port map (
            O => \N__8944\,
            I => \N__8941\
        );

    \I__818\ : LocalMux
    port map (
            O => \N__8941\,
            I => \transmit_module.X_DELTA_PATTERN_6\
        );

    \I__817\ : InMux
    port map (
            O => \N__8938\,
            I => \N__8935\
        );

    \I__816\ : LocalMux
    port map (
            O => \N__8935\,
            I => \N__8932\
        );

    \I__815\ : Odrv12
    port map (
            O => \N__8932\,
            I => \transmit_module.X_DELTA_PATTERN_5\
        );

    \I__814\ : InMux
    port map (
            O => \N__8929\,
            I => \N__8926\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__8926\,
            I => \transmit_module.X_DELTA_PATTERN_4\
        );

    \I__812\ : InMux
    port map (
            O => \N__8923\,
            I => \N__8920\
        );

    \I__811\ : LocalMux
    port map (
            O => \N__8920\,
            I => \transmit_module.X_DELTA_PATTERN_9\
        );

    \I__810\ : InMux
    port map (
            O => \N__8917\,
            I => \N__8914\
        );

    \I__809\ : LocalMux
    port map (
            O => \N__8914\,
            I => \transmit_module.Y_DELTA_PATTERN_87\
        );

    \I__808\ : InMux
    port map (
            O => \N__8911\,
            I => \N__8908\
        );

    \I__807\ : LocalMux
    port map (
            O => \N__8908\,
            I => \transmit_module.Y_DELTA_PATTERN_89\
        );

    \I__806\ : InMux
    port map (
            O => \N__8905\,
            I => \N__8902\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__8902\,
            I => \transmit_module.Y_DELTA_PATTERN_88\
        );

    \I__804\ : InMux
    port map (
            O => \N__8899\,
            I => \N__8896\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__8896\,
            I => \transmit_module.Y_DELTA_PATTERN_90\
        );

    \I__802\ : InMux
    port map (
            O => \N__8893\,
            I => \N__8890\
        );

    \I__801\ : LocalMux
    port map (
            O => \N__8890\,
            I => \transmit_module.Y_DELTA_PATTERN_91\
        );

    \I__800\ : InMux
    port map (
            O => \N__8887\,
            I => \N__8884\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__8884\,
            I => \transmit_module.Y_DELTA_PATTERN_77\
        );

    \I__798\ : InMux
    port map (
            O => \N__8881\,
            I => \N__8878\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__8878\,
            I => \N__8875\
        );

    \I__796\ : Span4Mux_s2_v
    port map (
            O => \N__8875\,
            I => \N__8871\
        );

    \I__795\ : InMux
    port map (
            O => \N__8874\,
            I => \N__8868\
        );

    \I__794\ : Span4Mux_v
    port map (
            O => \N__8871\,
            I => \N__8863\
        );

    \I__793\ : LocalMux
    port map (
            O => \N__8868\,
            I => \N__8863\
        );

    \I__792\ : Span4Mux_v
    port map (
            O => \N__8863\,
            I => \N__8859\
        );

    \I__791\ : InMux
    port map (
            O => \N__8862\,
            I => \N__8856\
        );

    \I__790\ : Span4Mux_v
    port map (
            O => \N__8859\,
            I => \N__8850\
        );

    \I__789\ : LocalMux
    port map (
            O => \N__8856\,
            I => \N__8850\
        );

    \I__788\ : InMux
    port map (
            O => \N__8855\,
            I => \N__8847\
        );

    \I__787\ : Span4Mux_v
    port map (
            O => \N__8850\,
            I => \N__8842\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__8847\,
            I => \N__8842\
        );

    \I__785\ : Span4Mux_v
    port map (
            O => \N__8842\,
            I => \N__8837\
        );

    \I__784\ : InMux
    port map (
            O => \N__8841\,
            I => \N__8834\
        );

    \I__783\ : InMux
    port map (
            O => \N__8840\,
            I => \N__8831\
        );

    \I__782\ : Span4Mux_v
    port map (
            O => \N__8837\,
            I => \N__8826\
        );

    \I__781\ : LocalMux
    port map (
            O => \N__8834\,
            I => \N__8826\
        );

    \I__780\ : LocalMux
    port map (
            O => \N__8831\,
            I => \N__8823\
        );

    \I__779\ : Span4Mux_h
    port map (
            O => \N__8826\,
            I => \N__8819\
        );

    \I__778\ : Span4Mux_h
    port map (
            O => \N__8823\,
            I => \N__8816\
        );

    \I__777\ : InMux
    port map (
            O => \N__8822\,
            I => \N__8813\
        );

    \I__776\ : Span4Mux_h
    port map (
            O => \N__8819\,
            I => \N__8810\
        );

    \I__775\ : Span4Mux_v
    port map (
            O => \N__8816\,
            I => \N__8806\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__8813\,
            I => \N__8803\
        );

    \I__773\ : Span4Mux_h
    port map (
            O => \N__8810\,
            I => \N__8800\
        );

    \I__772\ : InMux
    port map (
            O => \N__8809\,
            I => \N__8797\
        );

    \I__771\ : Span4Mux_v
    port map (
            O => \N__8806\,
            I => \N__8792\
        );

    \I__770\ : Span4Mux_h
    port map (
            O => \N__8803\,
            I => \N__8792\
        );

    \I__769\ : Span4Mux_h
    port map (
            O => \N__8800\,
            I => \N__8787\
        );

    \I__768\ : LocalMux
    port map (
            O => \N__8797\,
            I => \N__8787\
        );

    \I__767\ : Span4Mux_v
    port map (
            O => \N__8792\,
            I => \N__8784\
        );

    \I__766\ : Span4Mux_h
    port map (
            O => \N__8787\,
            I => \N__8781\
        );

    \I__765\ : Span4Mux_v
    port map (
            O => \N__8784\,
            I => \N__8778\
        );

    \I__764\ : Span4Mux_v
    port map (
            O => \N__8781\,
            I => \N__8775\
        );

    \I__763\ : Odrv4
    port map (
            O => \N__8778\,
            I => \TVP_VIDEO_c_2\
        );

    \I__762\ : Odrv4
    port map (
            O => \N__8775\,
            I => \TVP_VIDEO_c_2\
        );

    \I__761\ : InMux
    port map (
            O => \N__8770\,
            I => \N__8767\
        );

    \I__760\ : LocalMux
    port map (
            O => \N__8767\,
            I => \transmit_module.X_DELTA_PATTERN_3\
        );

    \I__759\ : InMux
    port map (
            O => \N__8764\,
            I => \N__8761\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__8761\,
            I => \N__8758\
        );

    \I__757\ : Odrv4
    port map (
            O => \N__8758\,
            I => \transmit_module.X_DELTA_PATTERN_2\
        );

    \I__756\ : InMux
    port map (
            O => \N__8755\,
            I => \N__8750\
        );

    \I__755\ : InMux
    port map (
            O => \N__8754\,
            I => \N__8747\
        );

    \I__754\ : InMux
    port map (
            O => \N__8753\,
            I => \N__8744\
        );

    \I__753\ : LocalMux
    port map (
            O => \N__8750\,
            I => \N__8741\
        );

    \I__752\ : LocalMux
    port map (
            O => \N__8747\,
            I => \N__8734\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__8744\,
            I => \N__8734\
        );

    \I__750\ : Span4Mux_v
    port map (
            O => \N__8741\,
            I => \N__8731\
        );

    \I__749\ : InMux
    port map (
            O => \N__8740\,
            I => \N__8728\
        );

    \I__748\ : InMux
    port map (
            O => \N__8739\,
            I => \N__8724\
        );

    \I__747\ : Span4Mux_v
    port map (
            O => \N__8734\,
            I => \N__8721\
        );

    \I__746\ : Span4Mux_v
    port map (
            O => \N__8731\,
            I => \N__8716\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__8728\,
            I => \N__8716\
        );

    \I__744\ : InMux
    port map (
            O => \N__8727\,
            I => \N__8713\
        );

    \I__743\ : LocalMux
    port map (
            O => \N__8724\,
            I => \N__8708\
        );

    \I__742\ : Span4Mux_v
    port map (
            O => \N__8721\,
            I => \N__8701\
        );

    \I__741\ : Span4Mux_v
    port map (
            O => \N__8716\,
            I => \N__8701\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__8713\,
            I => \N__8701\
        );

    \I__739\ : InMux
    port map (
            O => \N__8712\,
            I => \N__8698\
        );

    \I__738\ : InMux
    port map (
            O => \N__8711\,
            I => \N__8695\
        );

    \I__737\ : Span4Mux_v
    port map (
            O => \N__8708\,
            I => \N__8692\
        );

    \I__736\ : Span4Mux_v
    port map (
            O => \N__8701\,
            I => \N__8689\
        );

    \I__735\ : LocalMux
    port map (
            O => \N__8698\,
            I => \N__8686\
        );

    \I__734\ : LocalMux
    port map (
            O => \N__8695\,
            I => \N__8683\
        );

    \I__733\ : Sp12to4
    port map (
            O => \N__8692\,
            I => \N__8680\
        );

    \I__732\ : Span4Mux_v
    port map (
            O => \N__8689\,
            I => \N__8677\
        );

    \I__731\ : Span4Mux_h
    port map (
            O => \N__8686\,
            I => \N__8674\
        );

    \I__730\ : Span4Mux_h
    port map (
            O => \N__8683\,
            I => \N__8671\
        );

    \I__729\ : Span12Mux_h
    port map (
            O => \N__8680\,
            I => \N__8668\
        );

    \I__728\ : Sp12to4
    port map (
            O => \N__8677\,
            I => \N__8665\
        );

    \I__727\ : IoSpan4Mux
    port map (
            O => \N__8674\,
            I => \N__8662\
        );

    \I__726\ : Span4Mux_h
    port map (
            O => \N__8671\,
            I => \N__8659\
        );

    \I__725\ : Span12Mux_v
    port map (
            O => \N__8668\,
            I => \N__8654\
        );

    \I__724\ : Span12Mux_h
    port map (
            O => \N__8665\,
            I => \N__8654\
        );

    \I__723\ : IoSpan4Mux
    port map (
            O => \N__8662\,
            I => \N__8649\
        );

    \I__722\ : IoSpan4Mux
    port map (
            O => \N__8659\,
            I => \N__8649\
        );

    \I__721\ : Odrv12
    port map (
            O => \N__8654\,
            I => \TVP_VIDEO_c_8\
        );

    \I__720\ : Odrv4
    port map (
            O => \N__8649\,
            I => \TVP_VIDEO_c_8\
        );

    \I__719\ : InMux
    port map (
            O => \N__8644\,
            I => \N__8641\
        );

    \I__718\ : LocalMux
    port map (
            O => \N__8641\,
            I => \N__8636\
        );

    \I__717\ : InMux
    port map (
            O => \N__8640\,
            I => \N__8633\
        );

    \I__716\ : InMux
    port map (
            O => \N__8639\,
            I => \N__8630\
        );

    \I__715\ : Span4Mux_v
    port map (
            O => \N__8636\,
            I => \N__8621\
        );

    \I__714\ : LocalMux
    port map (
            O => \N__8633\,
            I => \N__8621\
        );

    \I__713\ : LocalMux
    port map (
            O => \N__8630\,
            I => \N__8621\
        );

    \I__712\ : InMux
    port map (
            O => \N__8629\,
            I => \N__8618\
        );

    \I__711\ : InMux
    port map (
            O => \N__8628\,
            I => \N__8615\
        );

    \I__710\ : Span4Mux_v
    port map (
            O => \N__8621\,
            I => \N__8609\
        );

    \I__709\ : LocalMux
    port map (
            O => \N__8618\,
            I => \N__8609\
        );

    \I__708\ : LocalMux
    port map (
            O => \N__8615\,
            I => \N__8606\
        );

    \I__707\ : InMux
    port map (
            O => \N__8614\,
            I => \N__8603\
        );

    \I__706\ : Span4Mux_h
    port map (
            O => \N__8609\,
            I => \N__8600\
        );

    \I__705\ : Span4Mux_h
    port map (
            O => \N__8606\,
            I => \N__8597\
        );

    \I__704\ : LocalMux
    port map (
            O => \N__8603\,
            I => \N__8594\
        );

    \I__703\ : Sp12to4
    port map (
            O => \N__8600\,
            I => \N__8588\
        );

    \I__702\ : Sp12to4
    port map (
            O => \N__8597\,
            I => \N__8588\
        );

    \I__701\ : Span12Mux_s8_h
    port map (
            O => \N__8594\,
            I => \N__8585\
        );

    \I__700\ : InMux
    port map (
            O => \N__8593\,
            I => \N__8582\
        );

    \I__699\ : Span12Mux_v
    port map (
            O => \N__8588\,
            I => \N__8579\
        );

    \I__698\ : Span12Mux_v
    port map (
            O => \N__8585\,
            I => \N__8576\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__8582\,
            I => \N__8573\
        );

    \I__696\ : Span12Mux_h
    port map (
            O => \N__8579\,
            I => \N__8569\
        );

    \I__695\ : Span12Mux_v
    port map (
            O => \N__8576\,
            I => \N__8566\
        );

    \I__694\ : Span4Mux_h
    port map (
            O => \N__8573\,
            I => \N__8563\
        );

    \I__693\ : InMux
    port map (
            O => \N__8572\,
            I => \N__8560\
        );

    \I__692\ : Odrv12
    port map (
            O => \N__8569\,
            I => \TVP_VIDEO_c_9\
        );

    \I__691\ : Odrv12
    port map (
            O => \N__8566\,
            I => \TVP_VIDEO_c_9\
        );

    \I__690\ : Odrv4
    port map (
            O => \N__8563\,
            I => \TVP_VIDEO_c_9\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__8560\,
            I => \TVP_VIDEO_c_9\
        );

    \I__688\ : InMux
    port map (
            O => \N__8551\,
            I => \N__8548\
        );

    \I__687\ : LocalMux
    port map (
            O => \N__8548\,
            I => \N__8545\
        );

    \I__686\ : Span4Mux_v
    port map (
            O => \N__8545\,
            I => \N__8541\
        );

    \I__685\ : InMux
    port map (
            O => \N__8544\,
            I => \N__8538\
        );

    \I__684\ : Span4Mux_v
    port map (
            O => \N__8541\,
            I => \N__8534\
        );

    \I__683\ : LocalMux
    port map (
            O => \N__8538\,
            I => \N__8529\
        );

    \I__682\ : InMux
    port map (
            O => \N__8537\,
            I => \N__8526\
        );

    \I__681\ : Span4Mux_v
    port map (
            O => \N__8534\,
            I => \N__8523\
        );

    \I__680\ : InMux
    port map (
            O => \N__8533\,
            I => \N__8520\
        );

    \I__679\ : InMux
    port map (
            O => \N__8532\,
            I => \N__8517\
        );

    \I__678\ : Span12Mux_h
    port map (
            O => \N__8529\,
            I => \N__8513\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__8526\,
            I => \N__8510\
        );

    \I__676\ : Span4Mux_v
    port map (
            O => \N__8523\,
            I => \N__8505\
        );

    \I__675\ : LocalMux
    port map (
            O => \N__8520\,
            I => \N__8505\
        );

    \I__674\ : LocalMux
    port map (
            O => \N__8517\,
            I => \N__8502\
        );

    \I__673\ : InMux
    port map (
            O => \N__8516\,
            I => \N__8497\
        );

    \I__672\ : Span12Mux_v
    port map (
            O => \N__8513\,
            I => \N__8494\
        );

    \I__671\ : Span4Mux_v
    port map (
            O => \N__8510\,
            I => \N__8491\
        );

    \I__670\ : Span4Mux_v
    port map (
            O => \N__8505\,
            I => \N__8488\
        );

    \I__669\ : Span12Mux_h
    port map (
            O => \N__8502\,
            I => \N__8485\
        );

    \I__668\ : InMux
    port map (
            O => \N__8501\,
            I => \N__8482\
        );

    \I__667\ : InMux
    port map (
            O => \N__8500\,
            I => \N__8479\
        );

    \I__666\ : LocalMux
    port map (
            O => \N__8497\,
            I => \N__8476\
        );

    \I__665\ : Span12Mux_v
    port map (
            O => \N__8494\,
            I => \N__8473\
        );

    \I__664\ : Sp12to4
    port map (
            O => \N__8491\,
            I => \N__8470\
        );

    \I__663\ : Sp12to4
    port map (
            O => \N__8488\,
            I => \N__8467\
        );

    \I__662\ : Span12Mux_v
    port map (
            O => \N__8485\,
            I => \N__8462\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__8482\,
            I => \N__8462\
        );

    \I__660\ : LocalMux
    port map (
            O => \N__8479\,
            I => \N__8459\
        );

    \I__659\ : Span4Mux_h
    port map (
            O => \N__8476\,
            I => \N__8456\
        );

    \I__658\ : Span12Mux_h
    port map (
            O => \N__8473\,
            I => \N__8453\
        );

    \I__657\ : Span12Mux_h
    port map (
            O => \N__8470\,
            I => \N__8448\
        );

    \I__656\ : Span12Mux_h
    port map (
            O => \N__8467\,
            I => \N__8448\
        );

    \I__655\ : Span12Mux_h
    port map (
            O => \N__8462\,
            I => \N__8443\
        );

    \I__654\ : Span12Mux_h
    port map (
            O => \N__8459\,
            I => \N__8443\
        );

    \I__653\ : Span4Mux_h
    port map (
            O => \N__8456\,
            I => \N__8440\
        );

    \I__652\ : Odrv12
    port map (
            O => \N__8453\,
            I => \TVP_VIDEO_c_7\
        );

    \I__651\ : Odrv12
    port map (
            O => \N__8448\,
            I => \TVP_VIDEO_c_7\
        );

    \I__650\ : Odrv12
    port map (
            O => \N__8443\,
            I => \TVP_VIDEO_c_7\
        );

    \I__649\ : Odrv4
    port map (
            O => \N__8440\,
            I => \TVP_VIDEO_c_7\
        );

    \I__648\ : InMux
    port map (
            O => \N__8431\,
            I => \N__8427\
        );

    \I__647\ : InMux
    port map (
            O => \N__8430\,
            I => \N__8424\
        );

    \I__646\ : LocalMux
    port map (
            O => \N__8427\,
            I => \N__8421\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__8424\,
            I => \N__8417\
        );

    \I__644\ : Span4Mux_v
    port map (
            O => \N__8421\,
            I => \N__8414\
        );

    \I__643\ : InMux
    port map (
            O => \N__8420\,
            I => \N__8411\
        );

    \I__642\ : Span4Mux_v
    port map (
            O => \N__8417\,
            I => \N__8407\
        );

    \I__641\ : Span4Mux_v
    port map (
            O => \N__8414\,
            I => \N__8402\
        );

    \I__640\ : LocalMux
    port map (
            O => \N__8411\,
            I => \N__8402\
        );

    \I__639\ : InMux
    port map (
            O => \N__8410\,
            I => \N__8399\
        );

    \I__638\ : Span4Mux_v
    port map (
            O => \N__8407\,
            I => \N__8396\
        );

    \I__637\ : Span4Mux_v
    port map (
            O => \N__8402\,
            I => \N__8390\
        );

    \I__636\ : LocalMux
    port map (
            O => \N__8399\,
            I => \N__8390\
        );

    \I__635\ : Span4Mux_v
    port map (
            O => \N__8396\,
            I => \N__8386\
        );

    \I__634\ : InMux
    port map (
            O => \N__8395\,
            I => \N__8383\
        );

    \I__633\ : Span4Mux_v
    port map (
            O => \N__8390\,
            I => \N__8379\
        );

    \I__632\ : InMux
    port map (
            O => \N__8389\,
            I => \N__8376\
        );

    \I__631\ : Span4Mux_v
    port map (
            O => \N__8386\,
            I => \N__8371\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__8383\,
            I => \N__8371\
        );

    \I__629\ : InMux
    port map (
            O => \N__8382\,
            I => \N__8368\
        );

    \I__628\ : Span4Mux_v
    port map (
            O => \N__8379\,
            I => \N__8363\
        );

    \I__627\ : LocalMux
    port map (
            O => \N__8376\,
            I => \N__8363\
        );

    \I__626\ : Span4Mux_v
    port map (
            O => \N__8371\,
            I => \N__8358\
        );

    \I__625\ : LocalMux
    port map (
            O => \N__8368\,
            I => \N__8358\
        );

    \I__624\ : Span4Mux_v
    port map (
            O => \N__8363\,
            I => \N__8354\
        );

    \I__623\ : Span4Mux_v
    port map (
            O => \N__8358\,
            I => \N__8351\
        );

    \I__622\ : InMux
    port map (
            O => \N__8357\,
            I => \N__8348\
        );

    \I__621\ : Sp12to4
    port map (
            O => \N__8354\,
            I => \N__8345\
        );

    \I__620\ : Span4Mux_v
    port map (
            O => \N__8351\,
            I => \N__8340\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__8348\,
            I => \N__8340\
        );

    \I__618\ : Span12Mux_h
    port map (
            O => \N__8345\,
            I => \N__8337\
        );

    \I__617\ : Span4Mux_h
    port map (
            O => \N__8340\,
            I => \N__8334\
        );

    \I__616\ : Odrv12
    port map (
            O => \N__8337\,
            I => \TVP_VIDEO_c_6\
        );

    \I__615\ : Odrv4
    port map (
            O => \N__8334\,
            I => \TVP_VIDEO_c_6\
        );

    \I__614\ : InMux
    port map (
            O => \N__8329\,
            I => \N__8326\
        );

    \I__613\ : LocalMux
    port map (
            O => \N__8326\,
            I => \N__8322\
        );

    \I__612\ : InMux
    port map (
            O => \N__8325\,
            I => \N__8318\
        );

    \I__611\ : Span4Mux_v
    port map (
            O => \N__8322\,
            I => \N__8315\
        );

    \I__610\ : InMux
    port map (
            O => \N__8321\,
            I => \N__8311\
        );

    \I__609\ : LocalMux
    port map (
            O => \N__8318\,
            I => \N__8308\
        );

    \I__608\ : Span4Mux_v
    port map (
            O => \N__8315\,
            I => \N__8304\
        );

    \I__607\ : InMux
    port map (
            O => \N__8314\,
            I => \N__8301\
        );

    \I__606\ : LocalMux
    port map (
            O => \N__8311\,
            I => \N__8298\
        );

    \I__605\ : Span4Mux_v
    port map (
            O => \N__8308\,
            I => \N__8295\
        );

    \I__604\ : InMux
    port map (
            O => \N__8307\,
            I => \N__8292\
        );

    \I__603\ : Span4Mux_v
    port map (
            O => \N__8304\,
            I => \N__8286\
        );

    \I__602\ : LocalMux
    port map (
            O => \N__8301\,
            I => \N__8286\
        );

    \I__601\ : Span4Mux_h
    port map (
            O => \N__8298\,
            I => \N__8282\
        );

    \I__600\ : Span4Mux_v
    port map (
            O => \N__8295\,
            I => \N__8277\
        );

    \I__599\ : LocalMux
    port map (
            O => \N__8292\,
            I => \N__8277\
        );

    \I__598\ : InMux
    port map (
            O => \N__8291\,
            I => \N__8274\
        );

    \I__597\ : Span4Mux_v
    port map (
            O => \N__8286\,
            I => \N__8271\
        );

    \I__596\ : InMux
    port map (
            O => \N__8285\,
            I => \N__8268\
        );

    \I__595\ : Sp12to4
    port map (
            O => \N__8282\,
            I => \N__8265\
        );

    \I__594\ : Span4Mux_v
    port map (
            O => \N__8277\,
            I => \N__8260\
        );

    \I__593\ : LocalMux
    port map (
            O => \N__8274\,
            I => \N__8260\
        );

    \I__592\ : Span4Mux_v
    port map (
            O => \N__8271\,
            I => \N__8255\
        );

    \I__591\ : LocalMux
    port map (
            O => \N__8268\,
            I => \N__8255\
        );

    \I__590\ : Span12Mux_v
    port map (
            O => \N__8265\,
            I => \N__8251\
        );

    \I__589\ : Span4Mux_v
    port map (
            O => \N__8260\,
            I => \N__8248\
        );

    \I__588\ : Span4Mux_v
    port map (
            O => \N__8255\,
            I => \N__8245\
        );

    \I__587\ : InMux
    port map (
            O => \N__8254\,
            I => \N__8242\
        );

    \I__586\ : Span12Mux_v
    port map (
            O => \N__8251\,
            I => \N__8237\
        );

    \I__585\ : Sp12to4
    port map (
            O => \N__8248\,
            I => \N__8237\
        );

    \I__584\ : Span4Mux_v
    port map (
            O => \N__8245\,
            I => \N__8232\
        );

    \I__583\ : LocalMux
    port map (
            O => \N__8242\,
            I => \N__8232\
        );

    \I__582\ : Span12Mux_h
    port map (
            O => \N__8237\,
            I => \N__8229\
        );

    \I__581\ : Span4Mux_h
    port map (
            O => \N__8232\,
            I => \N__8226\
        );

    \I__580\ : Odrv12
    port map (
            O => \N__8229\,
            I => \TVP_VIDEO_c_5\
        );

    \I__579\ : Odrv4
    port map (
            O => \N__8226\,
            I => \TVP_VIDEO_c_5\
        );

    \I__578\ : InMux
    port map (
            O => \N__8221\,
            I => \N__8218\
        );

    \I__577\ : LocalMux
    port map (
            O => \N__8218\,
            I => \N__8215\
        );

    \I__576\ : Span4Mux_v
    port map (
            O => \N__8215\,
            I => \N__8209\
        );

    \I__575\ : InMux
    port map (
            O => \N__8214\,
            I => \N__8206\
        );

    \I__574\ : InMux
    port map (
            O => \N__8213\,
            I => \N__8202\
        );

    \I__573\ : InMux
    port map (
            O => \N__8212\,
            I => \N__8198\
        );

    \I__572\ : Span4Mux_v
    port map (
            O => \N__8209\,
            I => \N__8193\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__8206\,
            I => \N__8193\
        );

    \I__570\ : InMux
    port map (
            O => \N__8205\,
            I => \N__8190\
        );

    \I__569\ : LocalMux
    port map (
            O => \N__8202\,
            I => \N__8187\
        );

    \I__568\ : InMux
    port map (
            O => \N__8201\,
            I => \N__8184\
        );

    \I__567\ : LocalMux
    port map (
            O => \N__8198\,
            I => \N__8181\
        );

    \I__566\ : Span4Mux_v
    port map (
            O => \N__8193\,
            I => \N__8176\
        );

    \I__565\ : LocalMux
    port map (
            O => \N__8190\,
            I => \N__8176\
        );

    \I__564\ : Span4Mux_h
    port map (
            O => \N__8187\,
            I => \N__8173\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__8184\,
            I => \N__8170\
        );

    \I__562\ : Span4Mux_s1_v
    port map (
            O => \N__8181\,
            I => \N__8166\
        );

    \I__561\ : Span4Mux_v
    port map (
            O => \N__8176\,
            I => \N__8163\
        );

    \I__560\ : Span4Mux_h
    port map (
            O => \N__8173\,
            I => \N__8160\
        );

    \I__559\ : Span4Mux_h
    port map (
            O => \N__8170\,
            I => \N__8157\
        );

    \I__558\ : InMux
    port map (
            O => \N__8169\,
            I => \N__8154\
        );

    \I__557\ : Sp12to4
    port map (
            O => \N__8166\,
            I => \N__8151\
        );

    \I__556\ : Span4Mux_h
    port map (
            O => \N__8163\,
            I => \N__8148\
        );

    \I__555\ : Span4Mux_h
    port map (
            O => \N__8160\,
            I => \N__8145\
        );

    \I__554\ : Span4Mux_v
    port map (
            O => \N__8157\,
            I => \N__8142\
        );

    \I__553\ : LocalMux
    port map (
            O => \N__8154\,
            I => \N__8139\
        );

    \I__552\ : Span12Mux_s10_h
    port map (
            O => \N__8151\,
            I => \N__8135\
        );

    \I__551\ : Sp12to4
    port map (
            O => \N__8148\,
            I => \N__8132\
        );

    \I__550\ : Span4Mux_h
    port map (
            O => \N__8145\,
            I => \N__8125\
        );

    \I__549\ : Span4Mux_v
    port map (
            O => \N__8142\,
            I => \N__8125\
        );

    \I__548\ : Span4Mux_h
    port map (
            O => \N__8139\,
            I => \N__8125\
        );

    \I__547\ : InMux
    port map (
            O => \N__8138\,
            I => \N__8122\
        );

    \I__546\ : Span12Mux_v
    port map (
            O => \N__8135\,
            I => \N__8119\
        );

    \I__545\ : Span12Mux_h
    port map (
            O => \N__8132\,
            I => \N__8116\
        );

    \I__544\ : Span4Mux_v
    port map (
            O => \N__8125\,
            I => \N__8113\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__8122\,
            I => \N__8110\
        );

    \I__542\ : Span12Mux_v
    port map (
            O => \N__8119\,
            I => \N__8107\
        );

    \I__541\ : Span12Mux_v
    port map (
            O => \N__8116\,
            I => \N__8104\
        );

    \I__540\ : Span4Mux_v
    port map (
            O => \N__8113\,
            I => \N__8101\
        );

    \I__539\ : Span4Mux_h
    port map (
            O => \N__8110\,
            I => \N__8098\
        );

    \I__538\ : Odrv12
    port map (
            O => \N__8107\,
            I => \TVP_VIDEO_c_4\
        );

    \I__537\ : Odrv12
    port map (
            O => \N__8104\,
            I => \TVP_VIDEO_c_4\
        );

    \I__536\ : Odrv4
    port map (
            O => \N__8101\,
            I => \TVP_VIDEO_c_4\
        );

    \I__535\ : Odrv4
    port map (
            O => \N__8098\,
            I => \TVP_VIDEO_c_4\
        );

    \I__534\ : InMux
    port map (
            O => \N__8089\,
            I => \N__8085\
        );

    \I__533\ : InMux
    port map (
            O => \N__8088\,
            I => \N__8082\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__8085\,
            I => \N__8078\
        );

    \I__531\ : LocalMux
    port map (
            O => \N__8082\,
            I => \N__8075\
        );

    \I__530\ : InMux
    port map (
            O => \N__8081\,
            I => \N__8072\
        );

    \I__529\ : Sp12to4
    port map (
            O => \N__8078\,
            I => \N__8068\
        );

    \I__528\ : Span4Mux_h
    port map (
            O => \N__8075\,
            I => \N__8065\
        );

    \I__527\ : LocalMux
    port map (
            O => \N__8072\,
            I => \N__8062\
        );

    \I__526\ : InMux
    port map (
            O => \N__8071\,
            I => \N__8058\
        );

    \I__525\ : Span12Mux_h
    port map (
            O => \N__8068\,
            I => \N__8053\
        );

    \I__524\ : Span4Mux_h
    port map (
            O => \N__8065\,
            I => \N__8050\
        );

    \I__523\ : Span4Mux_v
    port map (
            O => \N__8062\,
            I => \N__8047\
        );

    \I__522\ : InMux
    port map (
            O => \N__8061\,
            I => \N__8044\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__8058\,
            I => \N__8041\
        );

    \I__520\ : InMux
    port map (
            O => \N__8057\,
            I => \N__8038\
        );

    \I__519\ : InMux
    port map (
            O => \N__8056\,
            I => \N__8034\
        );

    \I__518\ : Span12Mux_v
    port map (
            O => \N__8053\,
            I => \N__8029\
        );

    \I__517\ : Sp12to4
    port map (
            O => \N__8050\,
            I => \N__8029\
        );

    \I__516\ : Sp12to4
    port map (
            O => \N__8047\,
            I => \N__8026\
        );

    \I__515\ : LocalMux
    port map (
            O => \N__8044\,
            I => \N__8023\
        );

    \I__514\ : Span12Mux_h
    port map (
            O => \N__8041\,
            I => \N__8020\
        );

    \I__513\ : LocalMux
    port map (
            O => \N__8038\,
            I => \N__8017\
        );

    \I__512\ : InMux
    port map (
            O => \N__8037\,
            I => \N__8014\
        );

    \I__511\ : LocalMux
    port map (
            O => \N__8034\,
            I => \N__8011\
        );

    \I__510\ : Span12Mux_v
    port map (
            O => \N__8029\,
            I => \N__8006\
        );

    \I__509\ : Span12Mux_h
    port map (
            O => \N__8026\,
            I => \N__8006\
        );

    \I__508\ : Span12Mux_h
    port map (
            O => \N__8023\,
            I => \N__8003\
        );

    \I__507\ : Span12Mux_v
    port map (
            O => \N__8020\,
            I => \N__7996\
        );

    \I__506\ : Span12Mux_h
    port map (
            O => \N__8017\,
            I => \N__7996\
        );

    \I__505\ : LocalMux
    port map (
            O => \N__8014\,
            I => \N__7996\
        );

    \I__504\ : Span4Mux_h
    port map (
            O => \N__8011\,
            I => \N__7993\
        );

    \I__503\ : Span12Mux_h
    port map (
            O => \N__8006\,
            I => \N__7988\
        );

    \I__502\ : Span12Mux_v
    port map (
            O => \N__8003\,
            I => \N__7988\
        );

    \I__501\ : Span12Mux_h
    port map (
            O => \N__7996\,
            I => \N__7985\
        );

    \I__500\ : Span4Mux_v
    port map (
            O => \N__7993\,
            I => \N__7982\
        );

    \I__499\ : Odrv12
    port map (
            O => \N__7988\,
            I => \TVP_VIDEO_c_3\
        );

    \I__498\ : Odrv12
    port map (
            O => \N__7985\,
            I => \TVP_VIDEO_c_3\
        );

    \I__497\ : Odrv4
    port map (
            O => \N__7982\,
            I => \TVP_VIDEO_c_3\
        );

    \INVsync_buffer.WIRE_OUT_8C\ : INV
    port map (
            O => \INVsync_buffer.WIRE_OUT_8C_net\,
            I => \N__22997\
        );

    \IN_MUX_bfv_12_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_13_0_\
        );

    \IN_MUX_bfv_12_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \transmit_module.video_signal_controller.n3297\,
            carryinitout => \bfn_12_14_0_\
        );

    \IN_MUX_bfv_10_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_15_0_\
        );

    \IN_MUX_bfv_10_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \transmit_module.video_signal_controller.n3286\,
            carryinitout => \bfn_10_16_0_\
        );

    \IN_MUX_bfv_15_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_13_0_\
        );

    \IN_MUX_bfv_15_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \transmit_module.n3265\,
            carryinitout => \bfn_15_14_0_\
        );

    \IN_MUX_bfv_13_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_10_0_\
        );

    \IN_MUX_bfv_13_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \receive_module.rx_counter.n3278\,
            carryinitout => \bfn_13_11_0_\
        );

    \IN_MUX_bfv_17_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_10_0_\
        );

    \IN_MUX_bfv_17_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \receive_module.rx_counter.n3308\,
            carryinitout => \bfn_17_11_0_\
        );

    \IN_MUX_bfv_16_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_5_0_\
        );

    \IN_MUX_bfv_15_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_11_0_\
        );

    \IN_MUX_bfv_15_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \receive_module.n3252\,
            carryinitout => \bfn_15_12_0_\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \transmit_module.X_DELTA_PATTERN_i1_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8764\,
            lcout => \transmit_module.X_DELTA_PATTERN_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23190\,
            ce => \N__11128\,
            sr => \N__21488\
        );

    \transmit_module.X_DELTA_PATTERN_i3_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8929\,
            lcout => \transmit_module.X_DELTA_PATTERN_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23224\,
            ce => \N__11122\,
            sr => \N__21458\
        );

    \transmit_module.X_DELTA_PATTERN_i2_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8770\,
            lcout => \transmit_module.X_DELTA_PATTERN_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23224\,
            ce => \N__11122\,
            sr => \N__21458\
        );

    \transmit_module.X_DELTA_PATTERN_i8_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8923\,
            lcout => \transmit_module.X_DELTA_PATTERN_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23224\,
            ce => \N__11122\,
            sr => \N__21458\
        );

    \transmit_module.X_DELTA_PATTERN_i4_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8938\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.X_DELTA_PATTERN_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23224\,
            ce => \N__11122\,
            sr => \N__21458\
        );

    \transmit_module.X_DELTA_PATTERN_i9_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8953\,
            lcout => \transmit_module.X_DELTA_PATTERN_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23224\,
            ce => \N__11122\,
            sr => \N__21458\
        );

    \transmit_module.Y_DELTA_PATTERN_i89_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8899\,
            lcout => \transmit_module.Y_DELTA_PATTERN_89\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23268\,
            ce => \N__11074\,
            sr => \N__21320\
        );

    \transmit_module.Y_DELTA_PATTERN_i86_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8917\,
            lcout => \transmit_module.Y_DELTA_PATTERN_86\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23268\,
            ce => \N__11074\,
            sr => \N__21320\
        );

    \transmit_module.Y_DELTA_PATTERN_i87_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8905\,
            lcout => \transmit_module.Y_DELTA_PATTERN_87\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23268\,
            ce => \N__11074\,
            sr => \N__21320\
        );

    \transmit_module.Y_DELTA_PATTERN_i88_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8911\,
            lcout => \transmit_module.Y_DELTA_PATTERN_88\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23268\,
            ce => \N__11074\,
            sr => \N__21320\
        );

    \transmit_module.Y_DELTA_PATTERN_i76_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8887\,
            lcout => \transmit_module.Y_DELTA_PATTERN_76\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23225\,
            ce => \N__11073\,
            sr => \N__21348\
        );

    \transmit_module.Y_DELTA_PATTERN_i90_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8893\,
            lcout => \transmit_module.Y_DELTA_PATTERN_90\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23225\,
            ce => \N__11073\,
            sr => \N__21348\
        );

    \transmit_module.Y_DELTA_PATTERN_i91_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8992\,
            lcout => \transmit_module.Y_DELTA_PATTERN_91\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23225\,
            ce => \N__11073\,
            sr => \N__21348\
        );

    \transmit_module.Y_DELTA_PATTERN_i77_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9319\,
            lcout => \transmit_module.Y_DELTA_PATTERN_77\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23225\,
            ce => \N__11073\,
            sr => \N__21348\
        );

    \transmit_module.Y_DELTA_PATTERN_i92_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8986\,
            lcout => \transmit_module.Y_DELTA_PATTERN_92\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23225\,
            ce => \N__11073\,
            sr => \N__21348\
        );

    \transmit_module.Y_DELTA_PATTERN_i93_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8974\,
            lcout => \transmit_module.Y_DELTA_PATTERN_93\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23160\,
            ce => \N__11069\,
            sr => \N__21351\
        );

    \transmit_module.Y_DELTA_PATTERN_i95_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9121\,
            lcout => \transmit_module.Y_DELTA_PATTERN_95\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23160\,
            ce => \N__11069\,
            sr => \N__21351\
        );

    \transmit_module.Y_DELTA_PATTERN_i94_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8980\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.Y_DELTA_PATTERN_94\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23080\,
            ce => \N__21460\,
            sr => \N__21304\
        );

    \transmit_module.X_DELTA_PATTERN_i7_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8968\,
            lcout => \transmit_module.X_DELTA_PATTERN_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23175\,
            ce => \N__11106\,
            sr => \N__21457\
        );

    \transmit_module.X_DELTA_PATTERN_i6_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8959\,
            lcout => \transmit_module.X_DELTA_PATTERN_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23175\,
            ce => \N__11106\,
            sr => \N__21457\
        );

    \transmit_module.X_DELTA_PATTERN_i15_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13426\,
            lcout => \transmit_module.X_DELTA_PATTERN_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23175\,
            ce => \N__11106\,
            sr => \N__21457\
        );

    \transmit_module.X_DELTA_PATTERN_i10_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9028\,
            lcout => \transmit_module.X_DELTA_PATTERN_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23175\,
            ce => \N__11106\,
            sr => \N__21457\
        );

    \transmit_module.X_DELTA_PATTERN_i5_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8944\,
            lcout => \transmit_module.X_DELTA_PATTERN_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23175\,
            ce => \N__11106\,
            sr => \N__21457\
        );

    \transmit_module.X_DELTA_PATTERN_i14_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9040\,
            lcout => \transmit_module.X_DELTA_PATTERN_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23175\,
            ce => \N__11106\,
            sr => \N__21457\
        );

    \transmit_module.X_DELTA_PATTERN_i12_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9016\,
            lcout => \transmit_module.X_DELTA_PATTERN_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23055\,
            ce => \N__11127\,
            sr => \N__21474\
        );

    \transmit_module.X_DELTA_PATTERN_i11_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9034\,
            lcout => \transmit_module.X_DELTA_PATTERN_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23055\,
            ce => \N__11127\,
            sr => \N__21474\
        );

    \transmit_module.X_DELTA_PATTERN_i13_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9022\,
            lcout => \transmit_module.X_DELTA_PATTERN_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23055\,
            ce => \N__11127\,
            sr => \N__21474\
        );

    \transmit_module.Y_DELTA_PATTERN_i40_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8998\,
            lcout => \transmit_module.Y_DELTA_PATTERN_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23151\,
            ce => \N__10051\,
            sr => \N__21350\
        );

    \transmit_module.Y_DELTA_PATTERN_i64_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9004\,
            lcout => \transmit_module.Y_DELTA_PATTERN_64\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23292\,
            ce => \N__10039\,
            sr => \N__21325\
        );

    \transmit_module.Y_DELTA_PATTERN_i63_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9010\,
            lcout => \transmit_module.Y_DELTA_PATTERN_63\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23292\,
            ce => \N__10039\,
            sr => \N__21325\
        );

    \transmit_module.Y_DELTA_PATTERN_i65_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9283\,
            lcout => \transmit_module.Y_DELTA_PATTERN_65\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23292\,
            ce => \N__10039\,
            sr => \N__21325\
        );

    \transmit_module.Y_DELTA_PATTERN_i41_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9130\,
            lcout => \transmit_module.Y_DELTA_PATTERN_41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23292\,
            ce => \N__10039\,
            sr => \N__21325\
        );

    \transmit_module.Y_DELTA_PATTERN_i62_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9088\,
            lcout => \transmit_module.Y_DELTA_PATTERN_62\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23292\,
            ce => \N__10039\,
            sr => \N__21325\
        );

    \transmit_module.Y_DELTA_PATTERN_i73_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9082\,
            lcout => \transmit_module.Y_DELTA_PATTERN_73\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23134\,
            ce => \N__10049\,
            sr => \N__21349\
        );

    \transmit_module.Y_DELTA_PATTERN_i74_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9070\,
            lcout => \transmit_module.Y_DELTA_PATTERN_74\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23134\,
            ce => \N__10049\,
            sr => \N__21349\
        );

    \transmit_module.Y_DELTA_PATTERN_i75_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9076\,
            lcout => \transmit_module.Y_DELTA_PATTERN_75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23134\,
            ce => \N__10049\,
            sr => \N__21349\
        );

    \transmit_module.Y_DELTA_PATTERN_i72_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9064\,
            lcout => \transmit_module.Y_DELTA_PATTERN_72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23134\,
            ce => \N__10049\,
            sr => \N__21349\
        );

    \transmit_module.Y_DELTA_PATTERN_i48_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9358\,
            lcout => \transmit_module.Y_DELTA_PATTERN_48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23134\,
            ce => \N__10049\,
            sr => \N__21349\
        );

    \transmit_module.Y_DELTA_PATTERN_i46_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9052\,
            lcout => \transmit_module.Y_DELTA_PATTERN_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23134\,
            ce => \N__10049\,
            sr => \N__21349\
        );

    \transmit_module.Y_DELTA_PATTERN_i47_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9058\,
            lcout => \transmit_module.Y_DELTA_PATTERN_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23134\,
            ce => \N__10049\,
            sr => \N__21349\
        );

    \transmit_module.Y_DELTA_PATTERN_i45_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9046\,
            lcout => \transmit_module.Y_DELTA_PATTERN_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23134\,
            ce => \N__10049\,
            sr => \N__21349\
        );

    \transmit_module.Y_DELTA_PATTERN_i42_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9103\,
            lcout => \transmit_module.Y_DELTA_PATTERN_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23201\,
            ce => \N__10054\,
            sr => \N__21347\
        );

    \transmit_module.Y_DELTA_PATTERN_i96_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9220\,
            lcout => \transmit_module.Y_DELTA_PATTERN_96\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23201\,
            ce => \N__10054\,
            sr => \N__21347\
        );

    \transmit_module.Y_DELTA_PATTERN_i44_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9115\,
            lcout => \transmit_module.Y_DELTA_PATTERN_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23201\,
            ce => \N__10054\,
            sr => \N__21347\
        );

    \transmit_module.Y_DELTA_PATTERN_i43_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9109\,
            lcout => \transmit_module.Y_DELTA_PATTERN_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23201\,
            ce => \N__10054\,
            sr => \N__21347\
        );

    \transmit_module.video_signal_controller.i1653_2_lut_3_lut_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9163\,
            in2 => \N__9190\,
            in3 => \N__9206\,
            lcout => \transmit_module.video_signal_controller.n2886\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_2_lut_adj_23_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9550\,
            in2 => \_gnd_net_\,
            in3 => \N__9415\,
            lcout => \transmit_module.video_signal_controller.n3467\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1643_2_lut_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__9207\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9188\,
            lcout => \transmit_module.video_signal_controller.n2876\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_2_lut_rep_21_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9662\,
            in2 => \_gnd_net_\,
            in3 => \N__9392\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n3788_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_4_lut_adj_25_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__9165\,
            in1 => \N__9421\,
            in2 => \N__9097\,
            in3 => \N__9094\,
            lcout => \transmit_module.video_signal_controller.n4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i495_2_lut_rep_22_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__9187\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9164\,
            lcout => \transmit_module.video_signal_controller.n3789\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.VGA_X_i0_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9208\,
            in2 => \_gnd_net_\,
            in3 => \N__9193\,
            lcout => \transmit_module.video_signal_controller.VGA_X_0\,
            ltout => OPEN,
            carryin => \bfn_10_15_0_\,
            carryout => \transmit_module.video_signal_controller.n3279\,
            clk => \N__23174\,
            ce => 'H',
            sr => \N__9790\
        );

    \transmit_module.video_signal_controller.VGA_X_i1_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9189\,
            in2 => \_gnd_net_\,
            in3 => \N__9169\,
            lcout => \transmit_module.video_signal_controller.VGA_X_1\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3279\,
            carryout => \transmit_module.video_signal_controller.n3280\,
            clk => \N__23174\,
            ce => 'H',
            sr => \N__9790\
        );

    \transmit_module.video_signal_controller.VGA_X_i2_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9166\,
            in2 => \_gnd_net_\,
            in3 => \N__9148\,
            lcout => \transmit_module.video_signal_controller.VGA_X_2\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3280\,
            carryout => \transmit_module.video_signal_controller.n3281\,
            clk => \N__23174\,
            ce => 'H',
            sr => \N__9790\
        );

    \transmit_module.video_signal_controller.VGA_X_i3_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9419\,
            in2 => \_gnd_net_\,
            in3 => \N__9145\,
            lcout => \transmit_module.video_signal_controller.VGA_X_3\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3281\,
            carryout => \transmit_module.video_signal_controller.n3282\,
            clk => \N__23174\,
            ce => 'H',
            sr => \N__9790\
        );

    \transmit_module.video_signal_controller.VGA_X_i4_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9551\,
            in2 => \_gnd_net_\,
            in3 => \N__9142\,
            lcout => \transmit_module.video_signal_controller.VGA_X_4\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3282\,
            carryout => \transmit_module.video_signal_controller.n3283\,
            clk => \N__23174\,
            ce => 'H',
            sr => \N__9790\
        );

    \transmit_module.video_signal_controller.VGA_X_i5_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9393\,
            in2 => \_gnd_net_\,
            in3 => \N__9139\,
            lcout => \transmit_module.video_signal_controller.VGA_X_5\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3283\,
            carryout => \transmit_module.video_signal_controller.n3284\,
            clk => \N__23174\,
            ce => 'H',
            sr => \N__9790\
        );

    \transmit_module.video_signal_controller.VGA_X_i6_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9663\,
            in2 => \_gnd_net_\,
            in3 => \N__9136\,
            lcout => \transmit_module.video_signal_controller.VGA_X_6\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3284\,
            carryout => \transmit_module.video_signal_controller.n3285\,
            clk => \N__23174\,
            ce => 'H',
            sr => \N__9790\
        );

    \transmit_module.video_signal_controller.VGA_X_i7_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9575\,
            in2 => \_gnd_net_\,
            in3 => \N__9133\,
            lcout => \transmit_module.video_signal_controller.VGA_X_7\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3285\,
            carryout => \transmit_module.video_signal_controller.n3286\,
            clk => \N__23174\,
            ce => 'H',
            sr => \N__9790\
        );

    \transmit_module.video_signal_controller.VGA_X_i8_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9688\,
            in2 => \_gnd_net_\,
            in3 => \N__9256\,
            lcout => \transmit_module.video_signal_controller.VGA_X_8\,
            ltout => OPEN,
            carryin => \bfn_10_16_0_\,
            carryout => \transmit_module.video_signal_controller.n3287\,
            clk => \N__23189\,
            ce => 'H',
            sr => \N__9786\
        );

    \transmit_module.video_signal_controller.VGA_X_i9_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9635\,
            in2 => \_gnd_net_\,
            in3 => \N__9253\,
            lcout => \transmit_module.video_signal_controller.VGA_X_9\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3287\,
            carryout => \transmit_module.video_signal_controller.n3288\,
            clk => \N__23189\,
            ce => 'H',
            sr => \N__9786\
        );

    \transmit_module.video_signal_controller.VGA_X_i10_LC_10_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9606\,
            in2 => \_gnd_net_\,
            in3 => \N__9250\,
            lcout => \transmit_module.video_signal_controller.VGA_X_10\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3288\,
            carryout => \transmit_module.video_signal_controller.n3289\,
            clk => \N__23189\,
            ce => 'H',
            sr => \N__9786\
        );

    \transmit_module.video_signal_controller.VGA_X_i11_LC_10_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10489\,
            in2 => \_gnd_net_\,
            in3 => \N__9247\,
            lcout => \transmit_module.video_signal_controller.VGA_X_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23189\,
            ce => 'H',
            sr => \N__9786\
        );

    \transmit_module.Y_DELTA_PATTERN_i53_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9238\,
            lcout => \transmit_module.Y_DELTA_PATTERN_53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23079\,
            ce => \N__10053\,
            sr => \N__21324\
        );

    \transmit_module.Y_DELTA_PATTERN_i55_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9226\,
            lcout => \transmit_module.Y_DELTA_PATTERN_55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23079\,
            ce => \N__10053\,
            sr => \N__21324\
        );

    \transmit_module.Y_DELTA_PATTERN_i54_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9244\,
            lcout => \transmit_module.Y_DELTA_PATTERN_54\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23079\,
            ce => \N__10053\,
            sr => \N__21324\
        );

    \transmit_module.Y_DELTA_PATTERN_i39_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9232\,
            lcout => \transmit_module.Y_DELTA_PATTERN_39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23199\,
            ce => \N__10052\,
            sr => \N__21330\
        );

    \transmit_module.Y_DELTA_PATTERN_i56_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__9496\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.Y_DELTA_PATTERN_56\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23199\,
            ce => \N__10052\,
            sr => \N__21330\
        );

    \transmit_module.Y_DELTA_PATTERN_i97_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9742\,
            lcout => \transmit_module.Y_DELTA_PATTERN_97\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23199\,
            ce => \N__10052\,
            sr => \N__21330\
        );

    \transmit_module.Y_DELTA_PATTERN_i35_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9295\,
            lcout => \transmit_module.Y_DELTA_PATTERN_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23199\,
            ce => \N__10052\,
            sr => \N__21330\
        );

    \transmit_module.Y_DELTA_PATTERN_i36_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9520\,
            lcout => \transmit_module.Y_DELTA_PATTERN_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23199\,
            ce => \N__10052\,
            sr => \N__21330\
        );

    \transmit_module.Y_DELTA_PATTERN_i61_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__9289\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.Y_DELTA_PATTERN_61\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23081\,
            ce => \N__10035\,
            sr => \N__21329\
        );

    \transmit_module.Y_DELTA_PATTERN_i66_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9472\,
            lcout => \transmit_module.Y_DELTA_PATTERN_66\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23081\,
            ce => \N__10035\,
            sr => \N__21329\
        );

    \transmit_module.Y_DELTA_PATTERN_i52_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9277\,
            lcout => \transmit_module.Y_DELTA_PATTERN_52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23081\,
            ce => \N__10035\,
            sr => \N__21329\
        );

    \transmit_module.Y_DELTA_PATTERN_i50_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9262\,
            lcout => \transmit_module.Y_DELTA_PATTERN_50\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23081\,
            ce => \N__10035\,
            sr => \N__21329\
        );

    \transmit_module.Y_DELTA_PATTERN_i51_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9268\,
            lcout => \transmit_module.Y_DELTA_PATTERN_51\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23081\,
            ce => \N__10035\,
            sr => \N__21329\
        );

    \transmit_module.Y_DELTA_PATTERN_i33_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9343\,
            lcout => \transmit_module.Y_DELTA_PATTERN_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23086\,
            ce => \N__10028\,
            sr => \N__21276\
        );

    \transmit_module.Y_DELTA_PATTERN_i81_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9331\,
            lcout => \transmit_module.Y_DELTA_PATTERN_81\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23086\,
            ce => \N__10028\,
            sr => \N__21276\
        );

    \transmit_module.Y_DELTA_PATTERN_i80_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9370\,
            lcout => \transmit_module.Y_DELTA_PATTERN_80\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23086\,
            ce => \N__10028\,
            sr => \N__21276\
        );

    \transmit_module.Y_DELTA_PATTERN_i49_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9364\,
            lcout => \transmit_module.Y_DELTA_PATTERN_49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23086\,
            ce => \N__10028\,
            sr => \N__21276\
        );

    \transmit_module.Y_DELTA_PATTERN_i34_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9352\,
            lcout => \transmit_module.Y_DELTA_PATTERN_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23086\,
            ce => \N__10028\,
            sr => \N__21276\
        );

    \transmit_module.Y_DELTA_PATTERN_i71_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9337\,
            lcout => \transmit_module.Y_DELTA_PATTERN_71\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23086\,
            ce => \N__10028\,
            sr => \N__21276\
        );

    \transmit_module.Y_DELTA_PATTERN_i82_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__9715\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.Y_DELTA_PATTERN_82\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23086\,
            ce => \N__10028\,
            sr => \N__21276\
        );

    \transmit_module.Y_DELTA_PATTERN_i69_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9484\,
            lcout => \transmit_module.Y_DELTA_PATTERN_69\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23077\,
            ce => \N__10024\,
            sr => \N__21331\
        );

    \transmit_module.Y_DELTA_PATTERN_i68_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9325\,
            lcout => \transmit_module.Y_DELTA_PATTERN_68\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23077\,
            ce => \N__10024\,
            sr => \N__21331\
        );

    \transmit_module.Y_DELTA_PATTERN_i78_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9301\,
            lcout => \transmit_module.Y_DELTA_PATTERN_78\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23077\,
            ce => \N__10024\,
            sr => \N__21331\
        );

    \transmit_module.Y_DELTA_PATTERN_i79_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9307\,
            lcout => \transmit_module.Y_DELTA_PATTERN_79\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23077\,
            ce => \N__10024\,
            sr => \N__21331\
        );

    \transmit_module.Y_DELTA_PATTERN_i70_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9490\,
            lcout => \transmit_module.Y_DELTA_PATTERN_70\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23077\,
            ce => \N__10024\,
            sr => \N__21331\
        );

    \transmit_module.Y_DELTA_PATTERN_i67_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9478\,
            lcout => \transmit_module.Y_DELTA_PATTERN_67\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23077\,
            ce => \N__10024\,
            sr => \N__21331\
        );

    \transmit_module.video_signal_controller.i1_2_lut_3_lut_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__9661\,
            in1 => \N__9391\,
            in2 => \_gnd_net_\,
            in3 => \N__9574\,
            lcout => \transmit_module.video_signal_controller.n1983\,
            ltout => \transmit_module.video_signal_controller.n1983_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1693_4_lut_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010100000"
        )
    port map (
            in0 => \N__9690\,
            in1 => \N__9463\,
            in2 => \N__9457\,
            in3 => \N__9432\,
            lcout => \transmit_module.video_signal_controller.n2926\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1699_4_lut_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101100"
        )
    port map (
            in0 => \N__9612\,
            in1 => \N__10490\,
            in2 => \N__9640\,
            in3 => \N__9454\,
            lcout => \transmit_module.video_signal_controller.n2010\,
            ltout => \transmit_module.video_signal_controller.n2010_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1136_2_lut_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17401\,
            in2 => \N__9448\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.video_signal_controller.n2361\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i483_4_lut_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000010100000"
        )
    port map (
            in0 => \N__9445\,
            in1 => \N__9439\,
            in2 => \N__9694\,
            in3 => \N__9433\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i2_4_lut_4_lut_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001111111110"
        )
    port map (
            in0 => \N__10491\,
            in1 => \N__9639\,
            in2 => \N__9424\,
            in3 => \N__9613\,
            lcout => \transmit_module.video_signal_controller.n7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_4_lut_adj_26_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110000"
        )
    port map (
            in0 => \N__9553\,
            in1 => \N__9420\,
            in2 => \N__9580\,
            in3 => \N__9394\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n4_adj_617_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.VGA_HS_66_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011101111"
        )
    port map (
            in0 => \N__9689\,
            in1 => \N__9532\,
            in2 => \N__9667\,
            in3 => \N__9664\,
            lcout => \ADV_HSYNC_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22972\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i2_3_lut_rep_27_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__9629\,
            in1 => \N__9602\,
            in2 => \_gnd_net_\,
            in3 => \N__10485\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n3794_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i2292_4_lut_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111000"
        )
    port map (
            in0 => \N__9586\,
            in1 => \N__9576\,
            in2 => \N__9556\,
            in3 => \N__9552\,
            lcout => \transmit_module.video_signal_controller.n3618\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.Y_DELTA_PATTERN_i60_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9526\,
            lcout => \transmit_module.Y_DELTA_PATTERN_60\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23082\,
            ce => \N__10050\,
            sr => \N__21319\
        );

    \transmit_module.Y_DELTA_PATTERN_i37_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9508\,
            lcout => \transmit_module.Y_DELTA_PATTERN_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23082\,
            ce => \N__10050\,
            sr => \N__21319\
        );

    \transmit_module.Y_DELTA_PATTERN_i38_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9514\,
            lcout => \transmit_module.Y_DELTA_PATTERN_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23082\,
            ce => \N__10050\,
            sr => \N__21319\
        );

    \transmit_module.Y_DELTA_PATTERN_i58_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9748\,
            lcout => \transmit_module.Y_DELTA_PATTERN_58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23082\,
            ce => \N__10050\,
            sr => \N__21319\
        );

    \transmit_module.Y_DELTA_PATTERN_i57_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9502\,
            lcout => \transmit_module.Y_DELTA_PATTERN_57\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23082\,
            ce => \N__10050\,
            sr => \N__21319\
        );

    \transmit_module.Y_DELTA_PATTERN_i59_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9754\,
            lcout => \transmit_module.Y_DELTA_PATTERN_59\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23082\,
            ce => \N__10050\,
            sr => \N__21319\
        );

    \transmit_module.Y_DELTA_PATTERN_i98_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9709\,
            lcout => \transmit_module.Y_DELTA_PATTERN_98\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22968\,
            ce => \N__11065\,
            sr => \N__21284\
        );

    \transmit_module.Y_DELTA_PATTERN_i85_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9736\,
            lcout => \transmit_module.Y_DELTA_PATTERN_85\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22968\,
            ce => \N__11065\,
            sr => \N__21284\
        );

    \transmit_module.Y_DELTA_PATTERN_i84_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9727\,
            lcout => \transmit_module.Y_DELTA_PATTERN_84\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22968\,
            ce => \N__11065\,
            sr => \N__21284\
        );

    \transmit_module.Y_DELTA_PATTERN_i83_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9721\,
            lcout => \transmit_module.Y_DELTA_PATTERN_83\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22968\,
            ce => \N__11065\,
            sr => \N__21284\
        );

    \transmit_module.Y_DELTA_PATTERN_i99_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17938\,
            lcout => \transmit_module.Y_DELTA_PATTERN_99\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23144\,
            ce => \N__21478\,
            sr => \N__21275\
        );

    \transmit_module.video_signal_controller.VGA_Y_i0_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11391\,
            in2 => \_gnd_net_\,
            in3 => \N__9703\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_0\,
            ltout => OPEN,
            carryin => \bfn_12_13_0_\,
            carryout => \transmit_module.video_signal_controller.n3290\,
            clk => \N__23101\,
            ce => \N__9778\,
            sr => \N__9850\
        );

    \transmit_module.video_signal_controller.VGA_Y_i1_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11348\,
            in2 => \_gnd_net_\,
            in3 => \N__9700\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_1\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3290\,
            carryout => \transmit_module.video_signal_controller.n3291\,
            clk => \N__23101\,
            ce => \N__9778\,
            sr => \N__9850\
        );

    \transmit_module.video_signal_controller.VGA_Y_i2_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10074\,
            in2 => \_gnd_net_\,
            in3 => \N__9697\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_2\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3291\,
            carryout => \transmit_module.video_signal_controller.n3292\,
            clk => \N__23101\,
            ce => \N__9778\,
            sr => \N__9850\
        );

    \transmit_module.video_signal_controller.VGA_Y_i3_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11377\,
            in2 => \_gnd_net_\,
            in3 => \N__9817\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_3\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3292\,
            carryout => \transmit_module.video_signal_controller.n3293\,
            clk => \N__23101\,
            ce => \N__9778\,
            sr => \N__9850\
        );

    \transmit_module.video_signal_controller.VGA_Y_i4_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11016\,
            in2 => \_gnd_net_\,
            in3 => \N__9814\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_4\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3293\,
            carryout => \transmit_module.video_signal_controller.n3294\,
            clk => \N__23101\,
            ce => \N__9778\,
            sr => \N__9850\
        );

    \transmit_module.video_signal_controller.VGA_Y_i5_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10095\,
            in2 => \_gnd_net_\,
            in3 => \N__9811\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_5\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3294\,
            carryout => \transmit_module.video_signal_controller.n3295\,
            clk => \N__23101\,
            ce => \N__9778\,
            sr => \N__9850\
        );

    \transmit_module.video_signal_controller.VGA_Y_i6_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10155\,
            in2 => \_gnd_net_\,
            in3 => \N__9808\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_6\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3295\,
            carryout => \transmit_module.video_signal_controller.n3296\,
            clk => \N__23101\,
            ce => \N__9778\,
            sr => \N__9850\
        );

    \transmit_module.video_signal_controller.VGA_Y_i7_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10119\,
            in2 => \_gnd_net_\,
            in3 => \N__9805\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_7\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3296\,
            carryout => \transmit_module.video_signal_controller.n3297\,
            clk => \N__23101\,
            ce => \N__9778\,
            sr => \N__9850\
        );

    \transmit_module.video_signal_controller.VGA_Y_i8_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10992\,
            in2 => \_gnd_net_\,
            in3 => \N__9802\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_8\,
            ltout => OPEN,
            carryin => \bfn_12_14_0_\,
            carryout => \transmit_module.video_signal_controller.n3298\,
            clk => \N__22990\,
            ce => \N__9782\,
            sr => \N__9849\
        );

    \transmit_module.video_signal_controller.VGA_Y_i9_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10178\,
            in2 => \_gnd_net_\,
            in3 => \N__9799\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_9\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3298\,
            carryout => \transmit_module.video_signal_controller.n3299\,
            clk => \N__22990\,
            ce => \N__9782\,
            sr => \N__9849\
        );

    \transmit_module.video_signal_controller.VGA_Y_i10_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11415\,
            in2 => \_gnd_net_\,
            in3 => \N__9796\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_10\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3299\,
            carryout => \transmit_module.video_signal_controller.n3300\,
            clk => \N__22990\,
            ce => \N__9782\,
            sr => \N__9849\
        );

    \transmit_module.video_signal_controller.VGA_Y_i11_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__10135\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9793\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22990\,
            ce => \N__9782\,
            sr => \N__9849\
        );

    \transmit_module.i2_3_lut_rep_20_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__10583\,
            in1 => \N__10609\,
            in2 => \_gnd_net_\,
            in3 => \N__10545\,
            lcout => \transmit_module.n3787\,
            ltout => \transmit_module.n3787_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i2_3_lut_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21120\,
            in2 => \N__9838\,
            in3 => \N__18298\,
            lcout => \transmit_module.n2093\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.old_VGA_HS_40_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10547\,
            lcout => \transmit_module.old_VGA_HS\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22961\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1_3_lut_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__21118\,
            in1 => \N__17933\,
            in2 => \_gnd_net_\,
            in3 => \N__18989\,
            lcout => \transmit_module.n2061\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i246_2_lut_4_lut_rep_30_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110011001100"
        )
    port map (
            in0 => \N__10546\,
            in1 => \N__21119\,
            in2 => \N__10615\,
            in3 => \N__10584\,
            lcout => \transmit_module.n3797\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.Y_DELTA_PATTERN_i7_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11533\,
            lcout => \transmit_module.Y_DELTA_PATTERN_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22938\,
            ce => \N__21449\,
            sr => \N__21195\
        );

    \transmit_module.Y_DELTA_PATTERN_i5_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9829\,
            lcout => \transmit_module.Y_DELTA_PATTERN_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22938\,
            ce => \N__21449\,
            sr => \N__21195\
        );

    \transmit_module.Y_DELTA_PATTERN_i6_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9835\,
            lcout => \transmit_module.Y_DELTA_PATTERN_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22938\,
            ce => \N__21449\,
            sr => \N__21195\
        );

    \transmit_module.Y_DELTA_PATTERN_i4_LC_12_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9823\,
            lcout => \transmit_module.Y_DELTA_PATTERN_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22938\,
            ce => \N__21449\,
            sr => \N__21195\
        );

    \transmit_module.Y_DELTA_PATTERN_i2_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9919\,
            lcout => \transmit_module.Y_DELTA_PATTERN_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22938\,
            ce => \N__21449\,
            sr => \N__21195\
        );

    \transmit_module.Y_DELTA_PATTERN_i3_LC_12_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9925\,
            lcout => \transmit_module.Y_DELTA_PATTERN_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22938\,
            ce => \N__21449\,
            sr => \N__21195\
        );

    \transmit_module.ADDR_Y_COMPONENT__i11_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23601\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23087\,
            ce => \N__17743\,
            sr => \N__21300\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__23630\,
            in1 => \N__9913\,
            in2 => \N__22233\,
            in3 => \N__9901\,
            lcout => \line_buffer.n3764\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2321_3_lut_LC_12_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__23639\,
            in1 => \N__9889\,
            in2 => \_gnd_net_\,
            in3 => \N__9877\,
            lcout => \line_buffer.n3647\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.Y__i0_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11178\,
            in2 => \_gnd_net_\,
            in3 => \N__9865\,
            lcout => \receive_module.rx_counter.Y_0\,
            ltout => OPEN,
            carryin => \bfn_13_10_0_\,
            carryout => \receive_module.rx_counter.n3271\,
            clk => \N__20141\,
            ce => \N__13092\,
            sr => \N__21947\
        );

    \receive_module.rx_counter.Y__i1_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11247\,
            in2 => \_gnd_net_\,
            in3 => \N__9862\,
            lcout => \receive_module.rx_counter.Y_1\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3271\,
            carryout => \receive_module.rx_counter.n3272\,
            clk => \N__20141\,
            ce => \N__13092\,
            sr => \N__21947\
        );

    \receive_module.rx_counter.Y__i2_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11266\,
            in2 => \_gnd_net_\,
            in3 => \N__9859\,
            lcout => \receive_module.rx_counter.Y_2\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3272\,
            carryout => \receive_module.rx_counter.n3273\,
            clk => \N__20141\,
            ce => \N__13092\,
            sr => \N__21947\
        );

    \receive_module.rx_counter.Y__i3_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11284\,
            in2 => \_gnd_net_\,
            in3 => \N__9856\,
            lcout => \receive_module.rx_counter.Y_3\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3273\,
            carryout => \receive_module.rx_counter.n3274\,
            clk => \N__20141\,
            ce => \N__13092\,
            sr => \N__21947\
        );

    \receive_module.rx_counter.Y__i4_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13122\,
            in2 => \_gnd_net_\,
            in3 => \N__9853\,
            lcout => \receive_module.rx_counter.Y_4\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3274\,
            carryout => \receive_module.rx_counter.n3275\,
            clk => \N__20141\,
            ce => \N__13092\,
            sr => \N__21947\
        );

    \receive_module.rx_counter.Y__i5_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11227\,
            in2 => \_gnd_net_\,
            in3 => \N__9940\,
            lcout => \receive_module.rx_counter.Y_5\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3275\,
            carryout => \receive_module.rx_counter.n3276\,
            clk => \N__20141\,
            ce => \N__13092\,
            sr => \N__21947\
        );

    \receive_module.rx_counter.Y__i6_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11212\,
            in2 => \_gnd_net_\,
            in3 => \N__9937\,
            lcout => \receive_module.rx_counter.Y_6\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3276\,
            carryout => \receive_module.rx_counter.n3277\,
            clk => \N__20141\,
            ce => \N__13092\,
            sr => \N__21947\
        );

    \receive_module.rx_counter.Y__i7_LC_13_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13164\,
            in2 => \_gnd_net_\,
            in3 => \N__9934\,
            lcout => \receive_module.rx_counter.Y_7\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3277\,
            carryout => \receive_module.rx_counter.n3278\,
            clk => \N__20141\,
            ce => \N__13092\,
            sr => \N__21947\
        );

    \receive_module.rx_counter.Y__i8_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16862\,
            in2 => \_gnd_net_\,
            in3 => \N__9931\,
            lcout => \receive_module.rx_counter.Y_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20145\,
            ce => \N__13096\,
            sr => \N__21956\
        );

    \transmit_module.ADDR_Y_COMPONENT__i7_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13543\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23274\,
            ce => \N__17774\,
            sr => \N__21261\
        );

    \transmit_module.video_signal_controller.i1_2_lut_rep_18_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__10118\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10988\,
            lcout => \transmit_module.video_signal_controller.n3785\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i2_2_lut_3_lut_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__10179\,
            in1 => \N__10981\,
            in2 => \_gnd_net_\,
            in3 => \N__10117\,
            lcout => \transmit_module.video_signal_controller.n8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_2_lut_rep_19_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11344\,
            in2 => \_gnd_net_\,
            in3 => \N__10072\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n3786_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_4_lut_adj_24_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101000"
        )
    port map (
            in0 => \N__11011\,
            in1 => \N__11379\,
            in2 => \N__9928\,
            in3 => \N__10188\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n7_adj_615_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i5_4_lut_LC_13_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__10094\,
            in1 => \N__10210\,
            in2 => \N__10204\,
            in3 => \N__10154\,
            lcout => \transmit_module.video_signal_controller.VGA_VISIBLE_N_578\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_2_lut_3_lut_adj_27_LC_13_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__10073\,
            in1 => \_gnd_net_\,
            in2 => \N__11352\,
            in3 => \N__11378\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i2_4_lut_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__10093\,
            in1 => \N__10153\,
            in2 => \N__10201\,
            in3 => \N__11012\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n3577_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_4_lut_LC_13_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101000"
        )
    port map (
            in0 => \N__10180\,
            in1 => \N__10198\,
            in2 => \N__10192\,
            in3 => \N__10189\,
            lcout => \transmit_module.video_signal_controller.n3486\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.VGA_VISIBLE_Y_64_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10521\,
            in2 => \_gnd_net_\,
            in3 => \N__10455\,
            lcout => \transmit_module.VGA_VISIBLE_Y\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23273\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_2_lut_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10133\,
            in2 => \_gnd_net_\,
            in3 => \N__11414\,
            lcout => \transmit_module.video_signal_controller.n3485\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i2288_2_lut_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10177\,
            in2 => \_gnd_net_\,
            in3 => \N__10156\,
            lcout => \transmit_module.video_signal_controller.n3614\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i2306_4_lut_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__10134\,
            in1 => \N__10120\,
            in2 => \N__10099\,
            in3 => \N__10075\,
            lcout => \transmit_module.video_signal_controller.n3632\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i246_2_lut_4_lut_rep_31_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110011001100"
        )
    port map (
            in0 => \N__10557\,
            in1 => \N__21059\,
            in2 => \N__10594\,
            in3 => \N__10614\,
            lcout => \transmit_module.n3798\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i5_3_lut_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__17905\,
            in1 => \N__10963\,
            in2 => \_gnd_net_\,
            in3 => \N__13338\,
            lcout => \transmit_module.n112\,
            ltout => \transmit_module.n112_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1603_4_lut_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001000100"
        )
    port map (
            in0 => \N__21004\,
            in1 => \N__11317\,
            in2 => \N__10837\,
            in3 => \N__18988\,
            lcout => n24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i246_2_lut_4_lut_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__10613\,
            in1 => \N__10590\,
            in2 => \N__21167\,
            in3 => \N__10556\,
            lcout => \transmit_module.n2147\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.VGA_VISIBLE_65_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__10525\,
            in1 => \N__10510\,
            in2 => \N__10498\,
            in3 => \N__10459\,
            lcout => \transmit_module.VGA_VISIBLE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23203\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i6_3_lut_LC_13_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__17906\,
            in1 => \N__10957\,
            in2 => \_gnd_net_\,
            in3 => \N__13305\,
            lcout => \transmit_module.n111\,
            ltout => \transmit_module.n111_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1604_4_lut_LC_13_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__18987\,
            in1 => \N__21005\,
            in2 => \N__10444\,
            in3 => \N__11295\,
            lcout => n23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.ADDR_Y_COMPONENT__i12_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22172\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23130\,
            ce => \N__17762\,
            sr => \N__21050\
        );

    \transmit_module.ADDR_Y_COMPONENT__i1_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13390\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23130\,
            ce => \N__17762\,
            sr => \N__21050\
        );

    \transmit_module.ADDR_Y_COMPONENT__i10_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13498\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23130\,
            ce => \N__17762\,
            sr => \N__21050\
        );

    \transmit_module.ADDR_Y_COMPONENT__i4_LC_13_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13342\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23130\,
            ce => \N__17762\,
            sr => \N__21050\
        );

    \transmit_module.ADDR_Y_COMPONENT__i5_LC_13_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13306\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23130\,
            ce => \N__17762\,
            sr => \N__21050\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_2422_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__23574\,
            in1 => \N__10951\,
            in2 => \N__22232\,
            in3 => \N__10936\,
            lcout => \line_buffer.n3752\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n3764_bdd_4_lut_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__10921\,
            in1 => \N__22215\,
            in2 => \N__10906\,
            in3 => \N__10885\,
            lcout => \line_buffer.n3767\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2320_3_lut_LC_13_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__23640\,
            in1 => \N__10879\,
            in2 => \_gnd_net_\,
            in3 => \N__10864\,
            lcout => OPEN,
            ltout => \line_buffer.n3646_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_12__bdd_4_lut_2397_LC_13_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001100100"
        )
    port map (
            in0 => \N__21683\,
            in1 => \N__22234\,
            in2 => \N__10846\,
            in3 => \N__10843\,
            lcout => \line_buffer.n3722\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i2_2_lut_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__13121\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13160\,
            lcout => \receive_module.rx_counter.n10_adj_610\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1_2_lut_adj_20_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__11282\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13120\,
            lcout => \receive_module.rx_counter.n4_adj_604\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i6_4_lut_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__11246\,
            in1 => \N__11283\,
            in2 => \N__16863\,
            in3 => \N__11265\,
            lcout => \receive_module.rx_counter.n14_adj_611\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i592_2_lut_rep_24_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11210\,
            in2 => \_gnd_net_\,
            in3 => \N__11225\,
            lcout => \receive_module.rx_counter.n3791\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i2_4_lut_adj_21_LC_14_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__11176\,
            in1 => \N__11281\,
            in2 => \N__11248\,
            in3 => \N__11263\,
            lcout => \receive_module.rx_counter.n3551\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i2_3_lut_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__11264\,
            in1 => \N__11177\,
            in2 => \_gnd_net_\,
            in3 => \N__11245\,
            lcout => \receive_module.rx_counter.n3548\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1_2_lut_3_lut_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__11226\,
            in1 => \N__13159\,
            in2 => \_gnd_net_\,
            in3 => \N__11211\,
            lcout => OPEN,
            ltout => \receive_module.rx_counter.n5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i3_4_lut_LC_14_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__16858\,
            in1 => \N__11194\,
            in2 => \N__11188\,
            in3 => \N__11185\,
            lcout => \receive_module.rx_counter.n3575\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.SYNC_46_LC_14_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__11179\,
            in1 => \N__11158\,
            in2 => \N__11152\,
            in3 => \N__13141\,
            lcout => \RX_TX_SYNC\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20142\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i8_3_lut_LC_14_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__17927\,
            in1 => \N__11143\,
            in2 => \_gnd_net_\,
            in3 => \N__13545\,
            lcout => \transmit_module.n109\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.X_DELTA_PATTERN_i0_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11137\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.X_DELTA_PATTERN_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23143\,
            ce => \N__11123\,
            sr => \N__11064\
        );

    \transmit_module.video_signal_controller.i2300_2_lut_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__11017\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10993\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n3626_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i7_4_lut_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000010"
        )
    port map (
            in0 => \N__11398\,
            in1 => \N__11380\,
            in2 => \N__11356\,
            in3 => \N__11353\,
            lcout => \transmit_module.video_signal_controller.n18_adj_616\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i0_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__19081\,
            in1 => \N__12078\,
            in2 => \N__21233\,
            in3 => \N__12051\,
            lcout => \transmit_module.TX_ADDR_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23100\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i7_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__19082\,
            in1 => \N__12801\,
            in2 => \N__21234\,
            in3 => \N__12777\,
            lcout => \transmit_module.TX_ADDR_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23100\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i5_LC_14_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001100100000"
        )
    port map (
            in0 => \N__11326\,
            in1 => \N__21131\,
            in2 => \N__19099\,
            in3 => \N__11296\,
            lcout => \transmit_module.TX_ADDR_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23100\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i2_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__19078\,
            in1 => \N__18577\,
            in2 => \N__21259\,
            in3 => \N__18556\,
            lcout => \transmit_module.TX_ADDR_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22989\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_14_i5_3_lut_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__13337\,
            in1 => \N__18273\,
            in2 => \_gnd_net_\,
            in3 => \N__13315\,
            lcout => \transmit_module.n143\,
            ltout => \transmit_module.n143_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i4_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__19079\,
            in1 => \N__21051\,
            in2 => \N__11305\,
            in3 => \N__11302\,
            lcout => \transmit_module.TX_ADDR_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22989\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_14_i6_3_lut_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__13297\,
            in1 => \N__18274\,
            in2 => \_gnd_net_\,
            in3 => \N__13276\,
            lcout => \transmit_module.n142\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i1_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__19077\,
            in1 => \N__11802\,
            in2 => \N__21258\,
            in3 => \N__11812\,
            lcout => \transmit_module.TX_ADDR_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22989\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_14_i7_3_lut_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__18300\,
            in1 => \N__13258\,
            in2 => \_gnd_net_\,
            in3 => \N__13234\,
            lcout => \transmit_module.n141\,
            ltout => \transmit_module.n141_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i6_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__19080\,
            in1 => \N__21052\,
            in2 => \N__11470\,
            in3 => \N__13053\,
            lcout => \transmit_module.TX_ADDR_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22989\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_14_i8_3_lut_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__18301\,
            in1 => \_gnd_net_\,
            in2 => \N__13546\,
            in3 => \N__13513\,
            lcout => \transmit_module.n140\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_14_i11_3_lut_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__18269\,
            in1 => \N__13496\,
            in2 => \_gnd_net_\,
            in3 => \N__13477\,
            lcout => \transmit_module.n137\,
            ltout => \transmit_module.n137_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i10_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__19023\,
            in1 => \N__21003\,
            in2 => \N__11467\,
            in3 => \N__12495\,
            lcout => \transmit_module.TX_ADDR_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23107\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i2_3_lut_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__13385\,
            in1 => \_gnd_net_\,
            in2 => \N__11464\,
            in3 => \N__17882\,
            lcout => \transmit_module.n115\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i11_3_lut_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100010111000"
        )
    port map (
            in0 => \N__13497\,
            in1 => \N__17881\,
            in2 => \N__11455\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.n106\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_14_i1_3_lut_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__13399\,
            in1 => \_gnd_net_\,
            in2 => \N__18299\,
            in3 => \N__13454\,
            lcout => \transmit_module.n147\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.VGA_VS_67_LC_14_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__11446\,
            in1 => \N__11440\,
            in2 => \N__11431\,
            in3 => \N__11422\,
            lcout => \ADV_VSYNC_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23107\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_14_i2_3_lut_LC_14_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__13384\,
            in1 => \_gnd_net_\,
            in2 => \N__13363\,
            in3 => \N__18294\,
            lcout => \transmit_module.n146\,
            ltout => \transmit_module.n146_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1600_4_lut_LC_14_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__19022\,
            in1 => \N__21002\,
            in2 => \N__11806\,
            in3 => \N__11803\,
            lcout => n27,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.Y_DELTA_PATTERN_i0_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11545\,
            lcout => \transmit_module.Y_DELTA_PATTERN_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22932\,
            ce => \N__21459\,
            sr => \N__21048\
        );

    \transmit_module.Y_DELTA_PATTERN_i9_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11524\,
            lcout => \transmit_module.Y_DELTA_PATTERN_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22932\,
            ce => \N__21459\,
            sr => \N__21048\
        );

    \transmit_module.Y_DELTA_PATTERN_i1_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11554\,
            lcout => \transmit_module.Y_DELTA_PATTERN_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22932\,
            ce => \N__21459\,
            sr => \N__21048\
        );

    \transmit_module.Y_DELTA_PATTERN_i8_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11539\,
            lcout => \transmit_module.Y_DELTA_PATTERN_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22932\,
            ce => \N__21459\,
            sr => \N__21048\
        );

    \transmit_module.Y_DELTA_PATTERN_i10_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19471\,
            lcout => \transmit_module.Y_DELTA_PATTERN_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22932\,
            ce => \N__21459\,
            sr => \N__21048\
        );

    \transmit_module.mux_12_i7_3_lut_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__17883\,
            in1 => \N__12505\,
            in2 => \_gnd_net_\,
            in3 => \N__13266\,
            lcout => \transmit_module.n110\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n3752_bdd_4_lut_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__11518\,
            in1 => \N__22125\,
            in2 => \N__11497\,
            in3 => \N__11476\,
            lcout => \line_buffer.n3755\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.ADDR_Y_COMPONENT__i6_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13267\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22979\,
            ce => \N__17770\,
            sr => \N__21117\
        );

    \transmit_module.ADDR_Y_COMPONENT__i0_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13456\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22979\,
            ce => \N__17770\,
            sr => \N__21117\
        );

    \transmit_module.i1609_4_lut_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__19093\,
            in1 => \N__12496\,
            in2 => \N__21205\,
            in3 => \N__12481\,
            lcout => n18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i1_3_lut_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__17908\,
            in1 => \N__12244\,
            in2 => \_gnd_net_\,
            in3 => \N__13455\,
            lcout => \transmit_module.n116\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i6_LC_14_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000001010"
        )
    port map (
            in0 => \N__12088\,
            in1 => \N__15679\,
            in2 => \N__21694\,
            in3 => \N__12238\,
            lcout => \TX_DATA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22747\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.VGA_R__i7_LC_14_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12232\,
            lcout => n1792,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22557\,
            ce => 'H',
            sr => \N__22319\
        );

    \transmit_module.VGA_R__i1_LC_14_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13807\,
            lcout => n1798,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22650\,
            ce => 'H',
            sr => \N__22321\
        );

    \line_buffer.i2353_3_lut_LC_14_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__12121\,
            in1 => \N__12103\,
            in2 => \_gnd_net_\,
            in3 => \N__23668\,
            lcout => \line_buffer.n3679\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1595_4_lut_LC_14_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__19109\,
            in1 => \N__12079\,
            in2 => \N__21280\,
            in3 => \N__12052\,
            lcout => n28,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1605_4_lut_LC_14_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__19113\,
            in1 => \N__13057\,
            in2 => \N__21281\,
            in3 => \N__13033\,
            lcout => n22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1606_4_lut_LC_14_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__19114\,
            in1 => \N__12805\,
            in2 => \N__21282\,
            in3 => \N__12781\,
            lcout => n21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.PULSE_1HZ_49_LC_15_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12543\,
            in2 => \_gnd_net_\,
            in3 => \N__12523\,
            lcout => \LED_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20128\,
            ce => \N__16266\,
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1_2_lut_LC_15_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16296\,
            in2 => \_gnd_net_\,
            in3 => \N__16326\,
            lcout => \receive_module.rx_counter.n7_adj_609\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i2302_2_lut_LC_15_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16278\,
            in2 => \_gnd_net_\,
            in3 => \N__16341\,
            lcout => OPEN,
            ltout => \receive_module.rx_counter.n3628_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i5_4_lut_LC_15_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__16356\,
            in1 => \N__16311\,
            in2 => \N__12532\,
            in3 => \N__12529\,
            lcout => \receive_module.rx_counter.n11\,
            ltout => \receive_module.rx_counter.n11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1286_2_lut_3_lut_LC_15_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__20462\,
            in1 => \_gnd_net_\,
            in2 => \N__12517\,
            in3 => \N__12513\,
            lcout => \receive_module.rx_counter.n2517\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.old_VS_52_LC_15_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20464\,
            lcout => \receive_module.rx_counter.old_VS\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20130\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i129_2_lut_rep_25_LC_15_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__12514\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20463\,
            lcout => \receive_module.rx_counter.n3792\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.O_VS_I_0_1_lut_rep_26_LC_15_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__20465\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \receive_module.n3793\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2315_3_lut_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__13198\,
            in1 => \N__13183\,
            in2 => \_gnd_net_\,
            in3 => \N__23659\,
            lcout => \line_buffer.n3641\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1_4_lut_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010001000"
        )
    port map (
            in0 => \N__13165\,
            in1 => \N__13140\,
            in2 => \N__13129\,
            in3 => \N__13102\,
            lcout => \receive_module.rx_counter.n4_adj_606\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i248_3_lut_3_lut_3_lut_LC_15_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101010101"
        )
    port map (
            in0 => \N__20483\,
            in1 => \N__18651\,
            in2 => \_gnd_net_\,
            in3 => \N__13075\,
            lcout => \receive_module.rx_counter.n2045\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.old_HS_51_LC_15_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__18652\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \receive_module.rx_counter.old_HS\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20137\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_2_lut_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16010\,
            in2 => \_gnd_net_\,
            in3 => \N__13069\,
            lcout => \receive_module.n136\,
            ltout => OPEN,
            carryin => \bfn_15_11_0_\,
            carryout => \receive_module.n3245\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_3_lut_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15758\,
            in2 => \_gnd_net_\,
            in3 => \N__13066\,
            lcout => \receive_module.n135\,
            ltout => OPEN,
            carryin => \receive_module.n3245\,
            carryout => \receive_module.n3246\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_4_lut_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13589\,
            in2 => \_gnd_net_\,
            in3 => \N__13063\,
            lcout => \receive_module.n134\,
            ltout => OPEN,
            carryin => \receive_module.n3246\,
            carryout => \receive_module.n3247\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_5_lut_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20240\,
            in3 => \N__13060\,
            lcout => \receive_module.n133\,
            ltout => OPEN,
            carryin => \receive_module.n3247\,
            carryout => \receive_module.n3248\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_6_lut_LC_15_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15218\,
            in2 => \_gnd_net_\,
            in3 => \N__13225\,
            lcout => \receive_module.n132\,
            ltout => OPEN,
            carryin => \receive_module.n3248\,
            carryout => \receive_module.n3249\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_7_lut_LC_15_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14990\,
            in2 => \_gnd_net_\,
            in3 => \N__13222\,
            lcout => \receive_module.n131\,
            ltout => OPEN,
            carryin => \receive_module.n3249\,
            carryout => \receive_module.n3250\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_8_lut_LC_15_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14714\,
            in3 => \N__13219\,
            lcout => \receive_module.n130\,
            ltout => OPEN,
            carryin => \receive_module.n3250\,
            carryout => \receive_module.n3251\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_9_lut_LC_15_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14462\,
            in2 => \_gnd_net_\,
            in3 => \N__13216\,
            lcout => \receive_module.n129\,
            ltout => OPEN,
            carryin => \receive_module.n3251\,
            carryout => \receive_module.n3252\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_10_lut_LC_15_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14210\,
            in2 => \_gnd_net_\,
            in3 => \N__13213\,
            lcout => \receive_module.n128\,
            ltout => OPEN,
            carryin => \bfn_15_12_0_\,
            carryout => \receive_module.n3253\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_11_lut_LC_15_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13976\,
            in2 => \_gnd_net_\,
            in3 => \N__13210\,
            lcout => \receive_module.n127\,
            ltout => OPEN,
            carryin => \receive_module.n3253\,
            carryout => \receive_module.n3254\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_12_lut_LC_15_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15479\,
            in2 => \_gnd_net_\,
            in3 => \N__13207\,
            lcout => \receive_module.n126\,
            ltout => OPEN,
            carryin => \receive_module.n3254\,
            carryout => \receive_module.n3255\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.BRAM_ADDR__i11_LC_15_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16685\,
            in2 => \_gnd_net_\,
            in3 => \N__13204\,
            lcout => \RX_ADDR_11\,
            ltout => OPEN,
            carryin => \receive_module.n3255\,
            carryout => \receive_module.n3256\,
            clk => \N__20143\,
            ce => \N__17053\,
            sr => \N__21946\
        );

    \receive_module.BRAM_ADDR__i12_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16784\,
            in2 => \_gnd_net_\,
            in3 => \N__13201\,
            lcout => \RX_ADDR_12\,
            ltout => OPEN,
            carryin => \receive_module.n3256\,
            carryout => \receive_module.n3257\,
            clk => \N__20143\,
            ce => \N__17053\,
            sr => \N__21946\
        );

    \receive_module.BRAM_ADDR__i13_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16737\,
            in2 => \_gnd_net_\,
            in3 => \N__13459\,
            lcout => \RX_ADDR_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20143\,
            ce => \N__17053\,
            sr => \N__21946\
        );

    \transmit_module.add_13_2_lut_LC_15_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13439\,
            in2 => \N__13422\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.n132\,
            ltout => OPEN,
            carryin => \bfn_15_13_0_\,
            carryout => \transmit_module.n3258\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_3_lut_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13389\,
            in3 => \N__13351\,
            lcout => \transmit_module.n131\,
            ltout => OPEN,
            carryin => \transmit_module.n3258\,
            carryout => \transmit_module.n3259\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_4_lut_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17955\,
            in2 => \_gnd_net_\,
            in3 => \N__13348\,
            lcout => \transmit_module.n130\,
            ltout => OPEN,
            carryin => \transmit_module.n3259\,
            carryout => \transmit_module.n3260\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_5_lut_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17796\,
            in2 => \_gnd_net_\,
            in3 => \N__13345\,
            lcout => \transmit_module.n129\,
            ltout => OPEN,
            carryin => \transmit_module.n3260\,
            carryout => \transmit_module.n3261\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_6_lut_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13336\,
            in2 => \_gnd_net_\,
            in3 => \N__13309\,
            lcout => \transmit_module.n128\,
            ltout => OPEN,
            carryin => \transmit_module.n3261\,
            carryout => \transmit_module.n3262\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_7_lut_LC_15_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13304\,
            in3 => \N__13270\,
            lcout => \transmit_module.n127\,
            ltout => OPEN,
            carryin => \transmit_module.n3262\,
            carryout => \transmit_module.n3263\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_8_lut_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13265\,
            in3 => \N__13228\,
            lcout => \transmit_module.n126\,
            ltout => OPEN,
            carryin => \transmit_module.n3263\,
            carryout => \transmit_module.n3264\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_9_lut_LC_15_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13544\,
            in3 => \N__13507\,
            lcout => \transmit_module.n125\,
            ltout => OPEN,
            carryin => \transmit_module.n3264\,
            carryout => \transmit_module.n3265\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_10_lut_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17353\,
            in3 => \N__13504\,
            lcout => \transmit_module.n124\,
            ltout => OPEN,
            carryin => \bfn_15_14_0_\,
            carryout => \transmit_module.n3266\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_11_lut_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17332\,
            in3 => \N__13501\,
            lcout => \transmit_module.n123\,
            ltout => OPEN,
            carryin => \transmit_module.n3266\,
            carryout => \transmit_module.n3267\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_12_lut_LC_15_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13495\,
            in2 => \_gnd_net_\,
            in3 => \N__13471\,
            lcout => \transmit_module.n122\,
            ltout => OPEN,
            carryin => \transmit_module.n3267\,
            carryout => \transmit_module.n3268\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_13_lut_LC_15_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23629\,
            in2 => \_gnd_net_\,
            in3 => \N__13468\,
            lcout => \transmit_module.n121\,
            ltout => OPEN,
            carryin => \transmit_module.n3268\,
            carryout => \transmit_module.n3269\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_14_lut_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22173\,
            in2 => \_gnd_net_\,
            in3 => \N__13465\,
            lcout => \transmit_module.n120\,
            ltout => OPEN,
            carryin => \transmit_module.n3269\,
            carryout => \transmit_module.n3270\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_15_lut_LC_15_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21645\,
            in2 => \_gnd_net_\,
            in3 => \N__13462\,
            lcout => \transmit_module.n119\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.ADDR_Y_COMPONENT__i9_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17329\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22982\,
            ce => \N__17766\,
            sr => \N__21053\
        );

    \transmit_module.ADDR_Y_COMPONENT__i8_LC_15_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17350\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22982\,
            ce => \N__17766\,
            sr => \N__21053\
        );

    \transmit_module.mux_12_i10_3_lut_LC_15_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__17884\,
            in1 => \N__13900\,
            in2 => \_gnd_net_\,
            in3 => \N__17331\,
            lcout => \transmit_module.n107\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1613_4_lut_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111110100"
        )
    port map (
            in0 => \N__17907\,
            in1 => \N__19024\,
            in2 => \N__21138\,
            in3 => \N__18307\,
            lcout => \transmit_module.n2039\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i12_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__13894\,
            in1 => \N__19097\,
            in2 => \_gnd_net_\,
            in3 => \N__13885\,
            lcout => \TX_ADDR_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22854\,
            ce => \N__13846\,
            sr => \N__21049\
        );

    \transmit_module.BRAM_ADDR__i13_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__17581\,
            in1 => \N__19098\,
            in2 => \_gnd_net_\,
            in3 => \N__13876\,
            lcout => \TX_ADDR_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22854\,
            ce => \N__13846\,
            sr => \N__21049\
        );

    \transmit_module.BRAM_ADDR__rep_1_i0_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__13867\,
            in1 => \N__19064\,
            in2 => \_gnd_net_\,
            in3 => \N__13855\,
            lcout => \TX_ADDR_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22872\,
            ce => \N__13842\,
            sr => \N__21235\
        );

    \transmit_module.mux_14_i3_3_lut_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__17979\,
            in1 => \N__18315\,
            in2 => \_gnd_net_\,
            in3 => \N__13822\,
            lcout => \transmit_module.n145\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i0_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__21652\,
            in1 => \N__13813\,
            in2 => \_gnd_net_\,
            in3 => \N__17521\,
            lcout => \TX_DATA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22833\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.BRAM_ADDR__i2_LC_15_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110010001100"
        )
    port map (
            in0 => \N__20672\,
            in1 => \N__13795\,
            in2 => \N__20503\,
            in3 => \N__13570\,
            lcout => \RX_ADDR_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20152\,
            ce => 'H',
            sr => \N__21979\
        );

    \transmit_module.video_signal_controller.i1120_1_lut_LC_15_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18316\,
            lcout => \transmit_module.n2354\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2354_3_lut_LC_15_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__15715\,
            in1 => \N__15700\,
            in2 => \_gnd_net_\,
            in3 => \N__23664\,
            lcout => \line_buffer.n3680\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.BRAM_ADDR__i10_LC_15_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111101000000"
        )
    port map (
            in0 => \N__20678\,
            in1 => \N__15442\,
            in2 => \N__20536\,
            in3 => \N__15673\,
            lcout => \RX_ADDR_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20158\,
            ce => 'H',
            sr => \N__21990\
        );

    \receive_module.BRAM_ADDR__i4_LC_15_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110010001100"
        )
    port map (
            in0 => \N__20693\,
            in1 => \N__15415\,
            in2 => \N__20567\,
            in3 => \N__15202\,
            lcout => \RX_ADDR_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20170\,
            ce => 'H',
            sr => \N__21997\
        );

    \receive_module.BRAM_ADDR__i5_LC_15_31_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011100010"
        )
    port map (
            in0 => \N__15178\,
            in1 => \N__20557\,
            in2 => \N__14956\,
            in3 => \N__20696\,
            lcout => \RX_ADDR_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20170\,
            ce => 'H',
            sr => \N__21997\
        );

    \receive_module.BRAM_ADDR__i6_LC_15_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111101000000"
        )
    port map (
            in0 => \N__20694\,
            in1 => \N__14686\,
            in2 => \N__20568\,
            in3 => \N__14914\,
            lcout => \RX_ADDR_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20170\,
            ce => 'H',
            sr => \N__21997\
        );

    \receive_module.BRAM_ADDR__i7_LC_15_31_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__20564\,
            in1 => \N__20697\,
            in2 => \N__14446\,
            in3 => \N__14662\,
            lcout => \RX_ADDR_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20170\,
            ce => 'H',
            sr => \N__21997\
        );

    \receive_module.BRAM_ADDR__i8_LC_15_31_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111101000000"
        )
    port map (
            in0 => \N__20695\,
            in1 => \N__14182\,
            in2 => \N__20569\,
            in3 => \N__14407\,
            lcout => \RX_ADDR_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20170\,
            ce => 'H',
            sr => \N__21997\
        );

    \receive_module.BRAM_ADDR__i9_LC_15_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__20565\,
            in1 => \N__20698\,
            in2 => \N__13942\,
            in3 => \N__14158\,
            lcout => \RX_ADDR_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20170\,
            ce => 'H',
            sr => \N__21997\
        );

    \receive_module.rx_counter.FRAME_COUNTER_243__i0_LC_16_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16357\,
            in2 => \_gnd_net_\,
            in3 => \N__16345\,
            lcout => \receive_module.rx_counter.FRAME_COUNTER_0\,
            ltout => OPEN,
            carryin => \bfn_16_5_0_\,
            carryout => \receive_module.rx_counter.n3310\,
            clk => \N__20129\,
            ce => \N__16267\,
            sr => \N__16243\
        );

    \receive_module.rx_counter.FRAME_COUNTER_243__i1_LC_16_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16342\,
            in2 => \_gnd_net_\,
            in3 => \N__16330\,
            lcout => \receive_module.rx_counter.FRAME_COUNTER_1\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3310\,
            carryout => \receive_module.rx_counter.n3311\,
            clk => \N__20129\,
            ce => \N__16267\,
            sr => \N__16243\
        );

    \receive_module.rx_counter.FRAME_COUNTER_243__i2_LC_16_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16327\,
            in2 => \_gnd_net_\,
            in3 => \N__16315\,
            lcout => \receive_module.rx_counter.FRAME_COUNTER_2\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3311\,
            carryout => \receive_module.rx_counter.n3312\,
            clk => \N__20129\,
            ce => \N__16267\,
            sr => \N__16243\
        );

    \receive_module.rx_counter.FRAME_COUNTER_243__i3_LC_16_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16312\,
            in2 => \_gnd_net_\,
            in3 => \N__16300\,
            lcout => \receive_module.rx_counter.FRAME_COUNTER_3\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3312\,
            carryout => \receive_module.rx_counter.n3313\,
            clk => \N__20129\,
            ce => \N__16267\,
            sr => \N__16243\
        );

    \receive_module.rx_counter.FRAME_COUNTER_243__i4_LC_16_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16297\,
            in2 => \_gnd_net_\,
            in3 => \N__16285\,
            lcout => \receive_module.rx_counter.FRAME_COUNTER_4\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3313\,
            carryout => \receive_module.rx_counter.n3314\,
            clk => \N__20129\,
            ce => \N__16267\,
            sr => \N__16243\
        );

    \receive_module.rx_counter.FRAME_COUNTER_243__i5_LC_16_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16279\,
            in2 => \_gnd_net_\,
            in3 => \N__16282\,
            lcout => \receive_module.rx_counter.FRAME_COUNTER_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20129\,
            ce => \N__16267\,
            sr => \N__16243\
        );

    \receive_module.BRAM_ADDR__i0_LC_16_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110010001100"
        )
    port map (
            in0 => \N__20673\,
            in1 => \N__16231\,
            in2 => \N__20535\,
            in3 => \N__15994\,
            lcout => \RX_ADDR_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20131\,
            ce => 'H',
            sr => \N__21933\
        );

    \receive_module.BRAM_ADDR__i1_LC_16_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010111000"
        )
    port map (
            in0 => \N__15751\,
            in1 => \N__20521\,
            in2 => \N__15973\,
            in3 => \N__20674\,
            lcout => \RX_ADDR_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20131\,
            ce => 'H',
            sr => \N__21933\
        );

    \line_buffer.i2308_3_lut_LC_16_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__23667\,
            in1 => \N__16573\,
            in2 => \_gnd_net_\,
            in3 => \N__16555\,
            lcout => \line_buffer.n3634\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2350_3_lut_LC_16_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__23655\,
            in1 => \N__16543\,
            in2 => \_gnd_net_\,
            in3 => \N__16525\,
            lcout => \line_buffer.n3676\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1_2_lut_adj_22_LC_16_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18593\,
            in2 => \_gnd_net_\,
            in3 => \N__19337\,
            lcout => OPEN,
            ltout => \receive_module.rx_counter.n4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i2_4_lut_LC_16_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__19320\,
            in1 => \N__19301\,
            in2 => \N__16510\,
            in3 => \N__19283\,
            lcout => \receive_module.rx_counter.n3581\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i2_2_lut_adj_19_LC_16_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19319\,
            in2 => \_gnd_net_\,
            in3 => \N__19338\,
            lcout => OPEN,
            ltout => \receive_module.rx_counter.n6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i2208_4_lut_LC_16_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__18594\,
            in1 => \N__19302\,
            in2 => \N__16507\,
            in3 => \N__19284\,
            lcout => \receive_module.rx_counter.n3534\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i59_4_lut_LC_16_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000110100001"
        )
    port map (
            in0 => \N__19266\,
            in1 => \N__16504\,
            in2 => \N__19249\,
            in3 => \N__16498\,
            lcout => \receive_module.rx_counter.n55_adj_607\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1_2_lut_3_lut_4_lut_adj_12_LC_16_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__16782\,
            in1 => \N__20635\,
            in2 => \N__16686\,
            in3 => \N__16735\,
            lcout => \line_buffer.n517\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1_2_lut_3_lut_4_lut_adj_17_LC_16_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__16678\,
            in1 => \N__16781\,
            in2 => \N__16741\,
            in3 => \N__20634\,
            lcout => \line_buffer.n452\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1_2_lut_3_lut_4_lut_adj_15_LC_16_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__16783\,
            in1 => \N__20636\,
            in2 => \N__16687\,
            in3 => \N__16736\,
            lcout => \line_buffer.n548\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.i245_2_lut_rep_28_LC_16_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__20631\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20534\,
            lcout => \receive_module.n3795\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1_2_lut_3_lut_4_lut_adj_14_LC_16_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__20629\,
            in1 => \N__16674\,
            in2 => \N__16785\,
            in3 => \N__16724\,
            lcout => \line_buffer.n451\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1_2_lut_3_lut_4_lut_adj_16_LC_16_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__20630\,
            in1 => \N__16675\,
            in2 => \N__16786\,
            in3 => \N__16725\,
            lcout => \line_buffer.n549\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1_2_lut_3_lut_4_lut_adj_13_LC_16_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__16673\,
            in1 => \N__16772\,
            in2 => \N__16738\,
            in3 => \N__20628\,
            lcout => \line_buffer.n516\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.O_VISIBLE_53_LC_16_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000101010"
        )
    port map (
            in0 => \N__16891\,
            in1 => \N__16879\,
            in2 => \N__16870\,
            in3 => \N__16834\,
            lcout => \RX_WE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20139\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1_2_lut_3_lut_4_lut_adj_11_LC_16_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__16677\,
            in1 => \N__16780\,
            in2 => \N__16740\,
            in3 => \N__20633\,
            lcout => \line_buffer.n581\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1_2_lut_3_lut_4_lut_LC_16_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__16779\,
            in1 => \N__20632\,
            in2 => \N__16739\,
            in3 => \N__16676\,
            lcout => \line_buffer.n580\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i3_LC_16_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__19068\,
            in1 => \N__17827\,
            in2 => \N__21268\,
            in3 => \N__18208\,
            lcout => \transmit_module.TX_ADDR_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22825\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sync_buffer.WIRE_OUT_8_LC_16_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17374\,
            lcout => \RX_TX_SYNC_BUFF\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVsync_buffer.WIRE_OUT_8C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sync_buffer.BUFFER_i0_LC_16_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17392\,
            lcout => \sync_buffer.BUFFER_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVsync_buffer.WIRE_OUT_8C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sync_buffer.BUFFER_i1_LC_16_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17380\,
            lcout => \sync_buffer.BUFFER_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVsync_buffer.WIRE_OUT_8C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_14_i9_3_lut_LC_16_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__18302\,
            in1 => \N__17351\,
            in2 => \_gnd_net_\,
            in3 => \N__17368\,
            lcout => \transmit_module.n139\,
            ltout => \transmit_module.n139_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i8_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__21055\,
            in1 => \N__19066\,
            in2 => \N__17362\,
            in3 => \N__18912\,
            lcout => \transmit_module.TX_ADDR_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22809\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i9_3_lut_LC_16_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__17928\,
            in1 => \N__17359\,
            in2 => \_gnd_net_\,
            in3 => \N__17352\,
            lcout => \transmit_module.n108\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i9_LC_16_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__19067\,
            in1 => \N__17293\,
            in2 => \N__21166\,
            in3 => \N__17302\,
            lcout => \transmit_module.TX_ADDR_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22809\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_14_i10_3_lut_LC_16_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__18303\,
            in1 => \N__17330\,
            in2 => \_gnd_net_\,
            in3 => \N__17308\,
            lcout => \transmit_module.n138\,
            ltout => \transmit_module.n138_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1608_4_lut_LC_16_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__21054\,
            in1 => \N__19065\,
            in2 => \N__17296\,
            in3 => \N__17292\,
            lcout => n19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.ADDR_Y_COMPONENT__i13_LC_16_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21644\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22853\,
            ce => \N__17779\,
            sr => \N__21266\
        );

    \line_buffer.TX_ADDR_12__bdd_4_lut_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__22124\,
            in1 => \N__19345\,
            in2 => \N__21675\,
            in3 => \N__17575\,
            lcout => \line_buffer.n3728\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n3746_bdd_4_lut_LC_16_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__17563\,
            in1 => \N__22123\,
            in2 => \N__17545\,
            in3 => \N__19414\,
            lcout => \line_buffer.n3749\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2348_3_lut_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__17515\,
            in1 => \N__17497\,
            in2 => \_gnd_net_\,
            in3 => \N__23543\,
            lcout => \line_buffer.n3674\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_12__bdd_4_lut_2392_LC_16_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011110010001100"
        )
    port map (
            in0 => \N__19378\,
            in1 => \N__22122\,
            in2 => \N__21674\,
            in3 => \N__17479\,
            lcout => \line_buffer.n3716\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i2_LC_16_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000001010"
        )
    port map (
            in0 => \N__19123\,
            in1 => \N__17467\,
            in2 => \N__21682\,
            in3 => \N__17461\,
            lcout => \TX_DATA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22883\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2314_3_lut_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__17455\,
            in1 => \N__17440\,
            in2 => \_gnd_net_\,
            in3 => \N__23544\,
            lcout => OPEN,
            ltout => \line_buffer.n3640_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i4_LC_16_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110010011000"
        )
    port map (
            in0 => \N__21661\,
            in1 => \N__17425\,
            in2 => \N__17419\,
            in3 => \N__17416\,
            lcout => \TX_DATA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22883\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i3_3_lut_LC_16_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__17929\,
            in1 => \N__17944\,
            in2 => \_gnd_net_\,
            in3 => \N__17972\,
            lcout => \transmit_module.n114\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1601_4_lut_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100001000"
        )
    port map (
            in0 => \N__18567\,
            in1 => \N__19059\,
            in2 => \N__21265\,
            in3 => \N__18549\,
            lcout => n26,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_14_i4_3_lut_LC_16_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__18314\,
            in1 => \N__17808\,
            in2 => \_gnd_net_\,
            in3 => \N__18220\,
            lcout => \transmit_module.n144\,
            ltout => \transmit_module.n144_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1602_4_lut_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__19060\,
            in1 => \N__21178\,
            in2 => \N__18196\,
            in3 => \N__17820\,
            lcout => n25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.ADDR_Y_COMPONENT__i2_LC_16_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17980\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22694\,
            ce => \N__17778\,
            sr => \N__21283\
        );

    \transmit_module.mux_12_i4_3_lut_LC_16_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__17807\,
            in1 => \N__17937\,
            in2 => \_gnd_net_\,
            in3 => \N__17785\,
            lcout => \transmit_module.n113\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.ADDR_Y_COMPONENT__i3_LC_16_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17809\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22694\,
            ce => \N__17778\,
            sr => \N__21283\
        );

    \transmit_module.VGA_R__i5_LC_16_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17707\,
            lcout => n1794,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22558\,
            ce => 'H',
            sr => \N__22315\
        );

    \transmit_module.VGA_R__i3_LC_16_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17638\,
            lcout => n1796,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22558\,
            ce => 'H',
            sr => \N__22315\
        );

    \line_buffer.i2347_3_lut_LC_16_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__19156\,
            in1 => \N__19141\,
            in2 => \_gnd_net_\,
            in3 => \N__23665\,
            lcout => \line_buffer.n3673\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1607_4_lut_LC_16_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__19086\,
            in1 => \N__18916\,
            in2 => \N__21318\,
            in3 => \N__18898\,
            lcout => n20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_TVP_CLK_c_THRU_LUT4_0_LC_16_32_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20182\,
            lcout => \GB_BUFFER_TVP_CLK_c_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i5_1_lut_rep_23_LC_17_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18645\,
            lcout => \receive_module.rx_counter.n3790\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.X_242__i0_LC_17_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18622\,
            in2 => \_gnd_net_\,
            in3 => \N__18616\,
            lcout => \receive_module.rx_counter.n10\,
            ltout => OPEN,
            carryin => \bfn_17_10_0_\,
            carryout => \receive_module.rx_counter.n3301\,
            clk => \N__20133\,
            ce => 'H',
            sr => \N__19234\
        );

    \receive_module.rx_counter.X_242__i1_LC_17_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18613\,
            in2 => \_gnd_net_\,
            in3 => \N__18607\,
            lcout => \receive_module.rx_counter.n9\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3301\,
            carryout => \receive_module.rx_counter.n3302\,
            clk => \N__20133\,
            ce => 'H',
            sr => \N__19234\
        );

    \receive_module.rx_counter.X_242__i2_LC_17_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18604\,
            in2 => \_gnd_net_\,
            in3 => \N__18598\,
            lcout => \receive_module.rx_counter.n8\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3302\,
            carryout => \receive_module.rx_counter.n3303\,
            clk => \N__20133\,
            ce => 'H',
            sr => \N__19234\
        );

    \receive_module.rx_counter.X_242__i3_LC_17_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18595\,
            in2 => \_gnd_net_\,
            in3 => \N__18580\,
            lcout => \receive_module.rx_counter.X_3\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3303\,
            carryout => \receive_module.rx_counter.n3304\,
            clk => \N__20133\,
            ce => 'H',
            sr => \N__19234\
        );

    \receive_module.rx_counter.X_242__i4_LC_17_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19339\,
            in2 => \_gnd_net_\,
            in3 => \N__19324\,
            lcout => \receive_module.rx_counter.X_4\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3304\,
            carryout => \receive_module.rx_counter.n3305\,
            clk => \N__20133\,
            ce => 'H',
            sr => \N__19234\
        );

    \receive_module.rx_counter.X_242__i5_LC_17_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19321\,
            in2 => \_gnd_net_\,
            in3 => \N__19306\,
            lcout => \receive_module.rx_counter.X_5\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3305\,
            carryout => \receive_module.rx_counter.n3306\,
            clk => \N__20133\,
            ce => 'H',
            sr => \N__19234\
        );

    \receive_module.rx_counter.X_242__i6_LC_17_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19303\,
            in2 => \_gnd_net_\,
            in3 => \N__19288\,
            lcout => \receive_module.rx_counter.X_6\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3306\,
            carryout => \receive_module.rx_counter.n3307\,
            clk => \N__20133\,
            ce => 'H',
            sr => \N__19234\
        );

    \receive_module.rx_counter.X_242__i7_LC_17_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19285\,
            in2 => \_gnd_net_\,
            in3 => \N__19270\,
            lcout => \receive_module.rx_counter.X_7\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3307\,
            carryout => \receive_module.rx_counter.n3308\,
            clk => \N__20133\,
            ce => 'H',
            sr => \N__19234\
        );

    \receive_module.rx_counter.X_242__i8_LC_17_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19267\,
            in2 => \_gnd_net_\,
            in3 => \N__19255\,
            lcout => \receive_module.rx_counter.X_8\,
            ltout => OPEN,
            carryin => \bfn_17_11_0_\,
            carryout => \receive_module.rx_counter.n3309\,
            clk => \N__20135\,
            ce => 'H',
            sr => \N__19233\
        );

    \receive_module.rx_counter.X_242__i9_LC_17_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19248\,
            in2 => \_gnd_net_\,
            in3 => \N__19252\,
            lcout => \receive_module.rx_counter.X_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20135\,
            ce => 'H',
            sr => \N__19233\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_2407_LC_17_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__23663\,
            in1 => \N__19213\,
            in2 => \N__22216\,
            in3 => \N__19204\,
            lcout => OPEN,
            ltout => \line_buffer.n3734_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n3734_bdd_4_lut_LC_17_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__19189\,
            in1 => \N__19174\,
            in2 => \N__19159\,
            in3 => \N__22178\,
            lcout => \line_buffer.n3737\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.Y_DELTA_PATTERN_i24_LC_17_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19459\,
            lcout => \transmit_module.Y_DELTA_PATTERN_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22994\,
            ce => \N__21482\,
            sr => \N__21303\
        );

    \transmit_module.Y_DELTA_PATTERN_i12_LC_17_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19447\,
            lcout => \transmit_module.Y_DELTA_PATTERN_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23073\,
            ce => \N__21461\,
            sr => \N__21171\
        );

    \transmit_module.Y_DELTA_PATTERN_i11_LC_17_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19477\,
            lcout => \transmit_module.Y_DELTA_PATTERN_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23073\,
            ce => \N__21461\,
            sr => \N__21171\
        );

    \transmit_module.Y_DELTA_PATTERN_i25_LC_17_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__19453\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.Y_DELTA_PATTERN_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23073\,
            ce => \N__21461\,
            sr => \N__21171\
        );

    \transmit_module.Y_DELTA_PATTERN_i26_LC_17_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__19504\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.Y_DELTA_PATTERN_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23073\,
            ce => \N__21461\,
            sr => \N__21171\
        );

    \transmit_module.Y_DELTA_PATTERN_i13_LC_17_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21565\,
            lcout => \transmit_module.Y_DELTA_PATTERN_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23073\,
            ce => \N__21461\,
            sr => \N__21171\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_2417_LC_17_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__23602\,
            in1 => \N__19441\,
            in2 => \N__22174\,
            in3 => \N__19429\,
            lcout => \line_buffer.n3746\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2351_3_lut_LC_17_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__23638\,
            in1 => \N__19408\,
            in2 => \_gnd_net_\,
            in3 => \N__19393\,
            lcout => \line_buffer.n3677\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2309_3_lut_LC_17_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__19372\,
            in1 => \N__23637\,
            in2 => \_gnd_net_\,
            in3 => \N__19360\,
            lcout => \line_buffer.n3635\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i5_LC_17_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__21684\,
            in1 => \N__19969\,
            in2 => \_gnd_net_\,
            in3 => \N__19924\,
            lcout => \TX_DATA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22843\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n3698_bdd_4_lut_LC_17_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__19960\,
            in1 => \N__22179\,
            in2 => \N__19945\,
            in3 => \N__20803\,
            lcout => \line_buffer.n3701\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.VGA_R__i6_LC_17_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19918\,
            lcout => n1793,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22690\,
            ce => 'H',
            sr => \N__22320\
        );

    \CONSTANT_ONE_LUT4_LC_17_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.Y_DELTA_PATTERN_i32_LC_18_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19519\,
            lcout => \transmit_module.Y_DELTA_PATTERN_32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23105\,
            ce => \N__21490\,
            sr => \N__21260\
        );

    \transmit_module.Y_DELTA_PATTERN_i27_LC_18_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19495\,
            lcout => \transmit_module.Y_DELTA_PATTERN_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23105\,
            ce => \N__21490\,
            sr => \N__21260\
        );

    \transmit_module.Y_DELTA_PATTERN_i28_LC_18_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19489\,
            lcout => \transmit_module.Y_DELTA_PATTERN_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23105\,
            ce => \N__21490\,
            sr => \N__21260\
        );

    \transmit_module.Y_DELTA_PATTERN_i29_LC_18_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19483\,
            lcout => \transmit_module.Y_DELTA_PATTERN_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23105\,
            ce => \N__21490\,
            sr => \N__21260\
        );

    \transmit_module.Y_DELTA_PATTERN_i30_LC_18_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20017\,
            lcout => \transmit_module.Y_DELTA_PATTERN_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23105\,
            ce => \N__21490\,
            sr => \N__21260\
        );

    \transmit_module.Y_DELTA_PATTERN_i31_LC_18_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20023\,
            lcout => \transmit_module.Y_DELTA_PATTERN_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23105\,
            ce => \N__21490\,
            sr => \N__21260\
        );

    \transmit_module.Y_DELTA_PATTERN_i22_LC_18_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19999\,
            lcout => \transmit_module.Y_DELTA_PATTERN_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22996\,
            ce => \N__21483\,
            sr => \N__21301\
        );

    \transmit_module.Y_DELTA_PATTERN_i21_LC_18_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20011\,
            lcout => \transmit_module.Y_DELTA_PATTERN_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22996\,
            ce => \N__21483\,
            sr => \N__21301\
        );

    \transmit_module.Y_DELTA_PATTERN_i23_LC_18_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20005\,
            lcout => \transmit_module.Y_DELTA_PATTERN_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22996\,
            ce => \N__21483\,
            sr => \N__21301\
        );

    \transmit_module.Y_DELTA_PATTERN_i15_LC_18_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19993\,
            lcout => \transmit_module.Y_DELTA_PATTERN_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22824\,
            ce => \N__21453\,
            sr => \N__21185\
        );

    \transmit_module.Y_DELTA_PATTERN_i19_LC_18_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__21496\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.Y_DELTA_PATTERN_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22824\,
            ce => \N__21453\,
            sr => \N__21185\
        );

    \transmit_module.Y_DELTA_PATTERN_i16_LC_18_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19987\,
            lcout => \transmit_module.Y_DELTA_PATTERN_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22824\,
            ce => \N__21453\,
            sr => \N__21185\
        );

    \transmit_module.Y_DELTA_PATTERN_i17_LC_18_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19975\,
            lcout => \transmit_module.Y_DELTA_PATTERN_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22824\,
            ce => \N__21453\,
            sr => \N__21185\
        );

    \transmit_module.Y_DELTA_PATTERN_i18_LC_18_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19981\,
            lcout => \transmit_module.Y_DELTA_PATTERN_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22824\,
            ce => \N__21453\,
            sr => \N__21185\
        );

    \transmit_module.Y_DELTA_PATTERN_i14_LC_18_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21571\,
            lcout => \transmit_module.Y_DELTA_PATTERN_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22947\,
            ce => \N__21484\,
            sr => \N__21302\
        );

    \transmit_module.VGA_R__i2_LC_18_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20752\,
            lcout => n1797,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22751\,
            ce => 'H',
            sr => \N__22322\
        );

    \transmit_module.Y_DELTA_PATTERN_i20_LC_19_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21502\,
            lcout => \transmit_module.Y_DELTA_PATTERN_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22995\,
            ce => \N__21489\,
            sr => \N__21267\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_2378_LC_19_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__23647\,
            in1 => \N__20833\,
            in2 => \N__22217\,
            in3 => \N__20818\,
            lcout => \line_buffer.n3698\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n3692_bdd_4_lut_LC_19_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__20791\,
            in1 => \N__22186\,
            in2 => \N__20776\,
            in3 => \N__20704\,
            lcout => OPEN,
            ltout => \line_buffer.n3695_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i1_LC_19_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21693\,
            in2 => \N__20755\,
            in3 => \N__21712\,
            lcout => \TX_DATA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22998\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_2373_LC_19_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__23653\,
            in1 => \N__20740\,
            in2 => \N__22218\,
            in3 => \N__20725\,
            lcout => \line_buffer.n3692\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.BRAM_ADDR__i3_LC_19_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110010001100"
        )
    port map (
            in0 => \N__20679\,
            in1 => \N__20584\,
            in2 => \N__20566\,
            in3 => \N__20209\,
            lcout => \RX_ADDR_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__20153\,
            ce => 'H',
            sr => \N__21989\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_2402_LC_20_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__23654\,
            in1 => \N__21904\,
            in2 => \N__22235\,
            in3 => \N__21892\,
            lcout => \line_buffer.n3710\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n3710_bdd_4_lut_LC_20_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__21883\,
            in1 => \N__22199\,
            in2 => \N__21868\,
            in3 => \N__21844\,
            lcout => \line_buffer.n3713\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_2427_LC_20_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100001011000"
        )
    port map (
            in0 => \N__22225\,
            in1 => \N__21838\,
            in2 => \N__23666\,
            in3 => \N__21820\,
            lcout => OPEN,
            ltout => \line_buffer.n3758_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n3758_bdd_4_lut_LC_20_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__21808\,
            in1 => \N__21790\,
            in2 => \N__21772\,
            in3 => \N__22227\,
            lcout => \line_buffer.n3761\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_2412_LC_20_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__23649\,
            in1 => \N__21769\,
            in2 => \N__22236\,
            in3 => \N__21757\,
            lcout => OPEN,
            ltout => \line_buffer.n3740_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n3740_bdd_4_lut_LC_20_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__21748\,
            in1 => \N__21730\,
            in2 => \N__21715\,
            in3 => \N__22226\,
            lcout => \line_buffer.n3743\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i3_LC_20_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__21691\,
            in1 => \N__21706\,
            in2 => \_gnd_net_\,
            in3 => \N__21700\,
            lcout => \TX_DATA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23096\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i7_LC_20_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__21692\,
            in1 => \N__21580\,
            in2 => \_gnd_net_\,
            in3 => \N__22003\,
            lcout => \TX_DATA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22981\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_2383_LC_20_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__23648\,
            in1 => \N__23473\,
            in2 => \N__22237\,
            in3 => \N__23458\,
            lcout => \line_buffer.n3704\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.VGA_R__i4_LC_20_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23443\,
            lcout => n1795,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22980\,
            ce => 'H',
            sr => \N__22326\
        );

    \transmit_module.VGA_R__i8_LC_20_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__23374\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ADV_B_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22832\,
            ce => 'H',
            sr => \N__22327\
        );

    \line_buffer.n3704_bdd_4_lut_LC_21_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__22252\,
            in1 => \N__22231\,
            in2 => \N__22030\,
            in3 => \N__22009\,
            lcout => \line_buffer.n3707\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
