// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     Sep 30 2018 19:20:56

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "main" view "INTERFACE"

module main (
    TVP_VIDEO,
    ADV_B,
    ADV_G,
    ADV_R,
    DEBUG,
    TVP_CLK,
    ADV_CLK,
    TVP_HSYNC,
    ADV_HSYNC,
    TVP_VSYNC,
    ADV_VSYNC,
    ADV_BLANK_N,
    LED,
    ADV_SYNC_N);

    input [9:0] TVP_VIDEO;
    output [7:0] ADV_B;
    output [7:0] ADV_G;
    output [7:0] ADV_R;
    inout [7:0] DEBUG;
    input TVP_CLK;
    output ADV_CLK;
    input TVP_HSYNC;
    output ADV_HSYNC;
    input TVP_VSYNC;
    output ADV_VSYNC;
    output ADV_BLANK_N;
    output LED;
    output ADV_SYNC_N;

    wire N__25256;
    wire N__25255;
    wire N__25254;
    wire N__25245;
    wire N__25244;
    wire N__25243;
    wire N__25236;
    wire N__25235;
    wire N__25234;
    wire N__25227;
    wire N__25226;
    wire N__25225;
    wire N__25218;
    wire N__25217;
    wire N__25216;
    wire N__25209;
    wire N__25208;
    wire N__25207;
    wire N__25200;
    wire N__25199;
    wire N__25198;
    wire N__25191;
    wire N__25190;
    wire N__25189;
    wire N__25182;
    wire N__25181;
    wire N__25180;
    wire N__25173;
    wire N__25172;
    wire N__25171;
    wire N__25164;
    wire N__25163;
    wire N__25162;
    wire N__25155;
    wire N__25154;
    wire N__25153;
    wire N__25146;
    wire N__25145;
    wire N__25144;
    wire N__25137;
    wire N__25136;
    wire N__25135;
    wire N__25128;
    wire N__25127;
    wire N__25126;
    wire N__25119;
    wire N__25118;
    wire N__25117;
    wire N__25110;
    wire N__25109;
    wire N__25108;
    wire N__25101;
    wire N__25100;
    wire N__25099;
    wire N__25092;
    wire N__25091;
    wire N__25090;
    wire N__25083;
    wire N__25082;
    wire N__25081;
    wire N__25074;
    wire N__25073;
    wire N__25072;
    wire N__25065;
    wire N__25064;
    wire N__25063;
    wire N__25056;
    wire N__25055;
    wire N__25054;
    wire N__25047;
    wire N__25046;
    wire N__25045;
    wire N__25038;
    wire N__25037;
    wire N__25036;
    wire N__25029;
    wire N__25028;
    wire N__25027;
    wire N__25020;
    wire N__25019;
    wire N__25018;
    wire N__25011;
    wire N__25010;
    wire N__25009;
    wire N__25002;
    wire N__25001;
    wire N__25000;
    wire N__24993;
    wire N__24992;
    wire N__24991;
    wire N__24984;
    wire N__24983;
    wire N__24982;
    wire N__24975;
    wire N__24974;
    wire N__24973;
    wire N__24966;
    wire N__24965;
    wire N__24964;
    wire N__24957;
    wire N__24956;
    wire N__24955;
    wire N__24948;
    wire N__24947;
    wire N__24946;
    wire N__24939;
    wire N__24938;
    wire N__24937;
    wire N__24930;
    wire N__24929;
    wire N__24928;
    wire N__24921;
    wire N__24920;
    wire N__24919;
    wire N__24912;
    wire N__24911;
    wire N__24910;
    wire N__24903;
    wire N__24902;
    wire N__24901;
    wire N__24894;
    wire N__24893;
    wire N__24892;
    wire N__24885;
    wire N__24884;
    wire N__24883;
    wire N__24876;
    wire N__24875;
    wire N__24874;
    wire N__24867;
    wire N__24866;
    wire N__24865;
    wire N__24858;
    wire N__24857;
    wire N__24856;
    wire N__24849;
    wire N__24848;
    wire N__24847;
    wire N__24840;
    wire N__24839;
    wire N__24838;
    wire N__24831;
    wire N__24830;
    wire N__24829;
    wire N__24822;
    wire N__24821;
    wire N__24820;
    wire N__24803;
    wire N__24800;
    wire N__24799;
    wire N__24798;
    wire N__24797;
    wire N__24796;
    wire N__24793;
    wire N__24792;
    wire N__24789;
    wire N__24786;
    wire N__24785;
    wire N__24784;
    wire N__24781;
    wire N__24778;
    wire N__24775;
    wire N__24772;
    wire N__24769;
    wire N__24766;
    wire N__24763;
    wire N__24760;
    wire N__24751;
    wire N__24748;
    wire N__24741;
    wire N__24738;
    wire N__24733;
    wire N__24728;
    wire N__24725;
    wire N__24722;
    wire N__24719;
    wire N__24716;
    wire N__24713;
    wire N__24710;
    wire N__24707;
    wire N__24704;
    wire N__24701;
    wire N__24698;
    wire N__24695;
    wire N__24692;
    wire N__24689;
    wire N__24686;
    wire N__24683;
    wire N__24680;
    wire N__24677;
    wire N__24674;
    wire N__24671;
    wire N__24668;
    wire N__24665;
    wire N__24664;
    wire N__24661;
    wire N__24658;
    wire N__24655;
    wire N__24652;
    wire N__24647;
    wire N__24644;
    wire N__24641;
    wire N__24638;
    wire N__24637;
    wire N__24636;
    wire N__24633;
    wire N__24632;
    wire N__24631;
    wire N__24630;
    wire N__24629;
    wire N__24628;
    wire N__24627;
    wire N__24626;
    wire N__24625;
    wire N__24624;
    wire N__24623;
    wire N__24622;
    wire N__24621;
    wire N__24620;
    wire N__24619;
    wire N__24618;
    wire N__24617;
    wire N__24616;
    wire N__24615;
    wire N__24614;
    wire N__24613;
    wire N__24612;
    wire N__24611;
    wire N__24610;
    wire N__24609;
    wire N__24608;
    wire N__24607;
    wire N__24606;
    wire N__24605;
    wire N__24604;
    wire N__24603;
    wire N__24602;
    wire N__24601;
    wire N__24600;
    wire N__24599;
    wire N__24598;
    wire N__24597;
    wire N__24596;
    wire N__24595;
    wire N__24594;
    wire N__24593;
    wire N__24592;
    wire N__24591;
    wire N__24590;
    wire N__24589;
    wire N__24588;
    wire N__24587;
    wire N__24586;
    wire N__24585;
    wire N__24584;
    wire N__24583;
    wire N__24582;
    wire N__24581;
    wire N__24580;
    wire N__24579;
    wire N__24578;
    wire N__24577;
    wire N__24576;
    wire N__24575;
    wire N__24574;
    wire N__24573;
    wire N__24572;
    wire N__24571;
    wire N__24570;
    wire N__24569;
    wire N__24568;
    wire N__24567;
    wire N__24566;
    wire N__24565;
    wire N__24564;
    wire N__24419;
    wire N__24416;
    wire N__24413;
    wire N__24410;
    wire N__24407;
    wire N__24404;
    wire N__24401;
    wire N__24398;
    wire N__24395;
    wire N__24392;
    wire N__24389;
    wire N__24386;
    wire N__24385;
    wire N__24384;
    wire N__24381;
    wire N__24380;
    wire N__24379;
    wire N__24378;
    wire N__24377;
    wire N__24374;
    wire N__24373;
    wire N__24370;
    wire N__24369;
    wire N__24368;
    wire N__24367;
    wire N__24364;
    wire N__24359;
    wire N__24358;
    wire N__24357;
    wire N__24354;
    wire N__24351;
    wire N__24348;
    wire N__24345;
    wire N__24344;
    wire N__24343;
    wire N__24342;
    wire N__24341;
    wire N__24340;
    wire N__24339;
    wire N__24338;
    wire N__24337;
    wire N__24336;
    wire N__24335;
    wire N__24332;
    wire N__24329;
    wire N__24326;
    wire N__24323;
    wire N__24320;
    wire N__24317;
    wire N__24314;
    wire N__24311;
    wire N__24310;
    wire N__24307;
    wire N__24304;
    wire N__24299;
    wire N__24296;
    wire N__24291;
    wire N__24290;
    wire N__24285;
    wire N__24282;
    wire N__24279;
    wire N__24276;
    wire N__24273;
    wire N__24270;
    wire N__24265;
    wire N__24262;
    wire N__24261;
    wire N__24254;
    wire N__24251;
    wire N__24248;
    wire N__24245;
    wire N__24242;
    wire N__24233;
    wire N__24230;
    wire N__24227;
    wire N__24224;
    wire N__24217;
    wire N__24210;
    wire N__24207;
    wire N__24202;
    wire N__24197;
    wire N__24194;
    wire N__24189;
    wire N__24184;
    wire N__24181;
    wire N__24178;
    wire N__24161;
    wire N__24158;
    wire N__24155;
    wire N__24152;
    wire N__24149;
    wire N__24146;
    wire N__24143;
    wire N__24140;
    wire N__24137;
    wire N__24136;
    wire N__24133;
    wire N__24130;
    wire N__24127;
    wire N__24126;
    wire N__24123;
    wire N__24120;
    wire N__24117;
    wire N__24114;
    wire N__24111;
    wire N__24108;
    wire N__24105;
    wire N__24100;
    wire N__24097;
    wire N__24094;
    wire N__24091;
    wire N__24086;
    wire N__24083;
    wire N__24080;
    wire N__24077;
    wire N__24074;
    wire N__24071;
    wire N__24068;
    wire N__24065;
    wire N__24062;
    wire N__24059;
    wire N__24056;
    wire N__24053;
    wire N__24050;
    wire N__24047;
    wire N__24044;
    wire N__24041;
    wire N__24038;
    wire N__24035;
    wire N__24032;
    wire N__24029;
    wire N__24026;
    wire N__24023;
    wire N__24020;
    wire N__24017;
    wire N__24016;
    wire N__24015;
    wire N__24012;
    wire N__24011;
    wire N__24010;
    wire N__24009;
    wire N__24008;
    wire N__24005;
    wire N__24002;
    wire N__23999;
    wire N__23998;
    wire N__23997;
    wire N__23996;
    wire N__23993;
    wire N__23990;
    wire N__23987;
    wire N__23986;
    wire N__23983;
    wire N__23980;
    wire N__23975;
    wire N__23974;
    wire N__23971;
    wire N__23968;
    wire N__23965;
    wire N__23960;
    wire N__23957;
    wire N__23954;
    wire N__23951;
    wire N__23950;
    wire N__23949;
    wire N__23946;
    wire N__23943;
    wire N__23940;
    wire N__23937;
    wire N__23928;
    wire N__23923;
    wire N__23920;
    wire N__23917;
    wire N__23914;
    wire N__23911;
    wire N__23902;
    wire N__23899;
    wire N__23888;
    wire N__23885;
    wire N__23882;
    wire N__23879;
    wire N__23876;
    wire N__23873;
    wire N__23870;
    wire N__23867;
    wire N__23864;
    wire N__23861;
    wire N__23858;
    wire N__23855;
    wire N__23852;
    wire N__23849;
    wire N__23848;
    wire N__23847;
    wire N__23846;
    wire N__23845;
    wire N__23844;
    wire N__23843;
    wire N__23842;
    wire N__23841;
    wire N__23840;
    wire N__23837;
    wire N__23834;
    wire N__23833;
    wire N__23832;
    wire N__23831;
    wire N__23828;
    wire N__23827;
    wire N__23826;
    wire N__23823;
    wire N__23820;
    wire N__23819;
    wire N__23818;
    wire N__23817;
    wire N__23816;
    wire N__23813;
    wire N__23810;
    wire N__23807;
    wire N__23806;
    wire N__23803;
    wire N__23798;
    wire N__23795;
    wire N__23792;
    wire N__23789;
    wire N__23784;
    wire N__23783;
    wire N__23780;
    wire N__23777;
    wire N__23774;
    wire N__23771;
    wire N__23768;
    wire N__23759;
    wire N__23756;
    wire N__23753;
    wire N__23750;
    wire N__23747;
    wire N__23742;
    wire N__23737;
    wire N__23734;
    wire N__23733;
    wire N__23730;
    wire N__23723;
    wire N__23712;
    wire N__23707;
    wire N__23704;
    wire N__23699;
    wire N__23696;
    wire N__23693;
    wire N__23686;
    wire N__23683;
    wire N__23680;
    wire N__23669;
    wire N__23666;
    wire N__23663;
    wire N__23660;
    wire N__23657;
    wire N__23654;
    wire N__23651;
    wire N__23648;
    wire N__23645;
    wire N__23642;
    wire N__23639;
    wire N__23636;
    wire N__23633;
    wire N__23630;
    wire N__23627;
    wire N__23624;
    wire N__23621;
    wire N__23618;
    wire N__23615;
    wire N__23612;
    wire N__23609;
    wire N__23606;
    wire N__23603;
    wire N__23602;
    wire N__23599;
    wire N__23596;
    wire N__23593;
    wire N__23592;
    wire N__23589;
    wire N__23586;
    wire N__23583;
    wire N__23580;
    wire N__23577;
    wire N__23574;
    wire N__23571;
    wire N__23568;
    wire N__23565;
    wire N__23562;
    wire N__23559;
    wire N__23556;
    wire N__23553;
    wire N__23546;
    wire N__23543;
    wire N__23542;
    wire N__23539;
    wire N__23536;
    wire N__23535;
    wire N__23530;
    wire N__23527;
    wire N__23526;
    wire N__23521;
    wire N__23518;
    wire N__23517;
    wire N__23516;
    wire N__23511;
    wire N__23508;
    wire N__23507;
    wire N__23506;
    wire N__23505;
    wire N__23502;
    wire N__23501;
    wire N__23500;
    wire N__23499;
    wire N__23498;
    wire N__23493;
    wire N__23490;
    wire N__23487;
    wire N__23486;
    wire N__23485;
    wire N__23484;
    wire N__23483;
    wire N__23482;
    wire N__23479;
    wire N__23476;
    wire N__23473;
    wire N__23472;
    wire N__23469;
    wire N__23468;
    wire N__23465;
    wire N__23464;
    wire N__23463;
    wire N__23460;
    wire N__23459;
    wire N__23458;
    wire N__23457;
    wire N__23456;
    wire N__23455;
    wire N__23450;
    wire N__23447;
    wire N__23444;
    wire N__23441;
    wire N__23440;
    wire N__23437;
    wire N__23436;
    wire N__23435;
    wire N__23434;
    wire N__23433;
    wire N__23430;
    wire N__23429;
    wire N__23428;
    wire N__23427;
    wire N__23426;
    wire N__23423;
    wire N__23422;
    wire N__23419;
    wire N__23414;
    wire N__23411;
    wire N__23408;
    wire N__23405;
    wire N__23404;
    wire N__23401;
    wire N__23398;
    wire N__23397;
    wire N__23394;
    wire N__23393;
    wire N__23392;
    wire N__23391;
    wire N__23390;
    wire N__23389;
    wire N__23386;
    wire N__23383;
    wire N__23380;
    wire N__23379;
    wire N__23378;
    wire N__23377;
    wire N__23376;
    wire N__23373;
    wire N__23372;
    wire N__23371;
    wire N__23368;
    wire N__23365;
    wire N__23364;
    wire N__23361;
    wire N__23354;
    wire N__23351;
    wire N__23348;
    wire N__23345;
    wire N__23342;
    wire N__23339;
    wire N__23336;
    wire N__23335;
    wire N__23332;
    wire N__23329;
    wire N__23328;
    wire N__23325;
    wire N__23322;
    wire N__23321;
    wire N__23320;
    wire N__23319;
    wire N__23318;
    wire N__23317;
    wire N__23316;
    wire N__23313;
    wire N__23312;
    wire N__23309;
    wire N__23306;
    wire N__23305;
    wire N__23304;
    wire N__23303;
    wire N__23302;
    wire N__23295;
    wire N__23290;
    wire N__23287;
    wire N__23282;
    wire N__23279;
    wire N__23276;
    wire N__23273;
    wire N__23270;
    wire N__23267;
    wire N__23264;
    wire N__23263;
    wire N__23262;
    wire N__23259;
    wire N__23254;
    wire N__23251;
    wire N__23248;
    wire N__23245;
    wire N__23242;
    wire N__23239;
    wire N__23236;
    wire N__23233;
    wire N__23230;
    wire N__23229;
    wire N__23228;
    wire N__23227;
    wire N__23222;
    wire N__23219;
    wire N__23218;
    wire N__23213;
    wire N__23206;
    wire N__23201;
    wire N__23198;
    wire N__23195;
    wire N__23194;
    wire N__23191;
    wire N__23188;
    wire N__23185;
    wire N__23184;
    wire N__23183;
    wire N__23182;
    wire N__23179;
    wire N__23176;
    wire N__23173;
    wire N__23170;
    wire N__23169;
    wire N__23166;
    wire N__23165;
    wire N__23162;
    wire N__23161;
    wire N__23158;
    wire N__23155;
    wire N__23154;
    wire N__23151;
    wire N__23148;
    wire N__23147;
    wire N__23142;
    wire N__23139;
    wire N__23136;
    wire N__23133;
    wire N__23132;
    wire N__23131;
    wire N__23130;
    wire N__23129;
    wire N__23126;
    wire N__23125;
    wire N__23124;
    wire N__23123;
    wire N__23112;
    wire N__23105;
    wire N__23102;
    wire N__23099;
    wire N__23096;
    wire N__23093;
    wire N__23092;
    wire N__23091;
    wire N__23088;
    wire N__23081;
    wire N__23078;
    wire N__23075;
    wire N__23072;
    wire N__23065;
    wire N__23062;
    wire N__23061;
    wire N__23058;
    wire N__23057;
    wire N__23054;
    wire N__23049;
    wire N__23046;
    wire N__23035;
    wire N__23032;
    wire N__23031;
    wire N__23026;
    wire N__23023;
    wire N__23020;
    wire N__23019;
    wire N__23016;
    wire N__23015;
    wire N__23012;
    wire N__23011;
    wire N__23004;
    wire N__23001;
    wire N__22998;
    wire N__22997;
    wire N__22994;
    wire N__22991;
    wire N__22988;
    wire N__22985;
    wire N__22980;
    wire N__22977;
    wire N__22976;
    wire N__22973;
    wire N__22970;
    wire N__22969;
    wire N__22966;
    wire N__22961;
    wire N__22956;
    wire N__22953;
    wire N__22950;
    wire N__22947;
    wire N__22944;
    wire N__22941;
    wire N__22938;
    wire N__22937;
    wire N__22936;
    wire N__22933;
    wire N__22932;
    wire N__22929;
    wire N__22922;
    wire N__22915;
    wire N__22912;
    wire N__22911;
    wire N__22910;
    wire N__22907;
    wire N__22900;
    wire N__22891;
    wire N__22888;
    wire N__22885;
    wire N__22882;
    wire N__22879;
    wire N__22870;
    wire N__22867;
    wire N__22860;
    wire N__22857;
    wire N__22854;
    wire N__22851;
    wire N__22848;
    wire N__22845;
    wire N__22844;
    wire N__22837;
    wire N__22834;
    wire N__22833;
    wire N__22824;
    wire N__22819;
    wire N__22816;
    wire N__22811;
    wire N__22808;
    wire N__22805;
    wire N__22796;
    wire N__22793;
    wire N__22786;
    wire N__22783;
    wire N__22780;
    wire N__22779;
    wire N__22776;
    wire N__22773;
    wire N__22772;
    wire N__22769;
    wire N__22764;
    wire N__22761;
    wire N__22758;
    wire N__22755;
    wire N__22752;
    wire N__22751;
    wire N__22748;
    wire N__22745;
    wire N__22742;
    wire N__22739;
    wire N__22736;
    wire N__22729;
    wire N__22724;
    wire N__22719;
    wire N__22714;
    wire N__22711;
    wire N__22710;
    wire N__22707;
    wire N__22704;
    wire N__22701;
    wire N__22700;
    wire N__22693;
    wire N__22688;
    wire N__22675;
    wire N__22672;
    wire N__22669;
    wire N__22666;
    wire N__22663;
    wire N__22654;
    wire N__22651;
    wire N__22648;
    wire N__22645;
    wire N__22644;
    wire N__22637;
    wire N__22632;
    wire N__22625;
    wire N__22620;
    wire N__22617;
    wire N__22612;
    wire N__22609;
    wire N__22606;
    wire N__22597;
    wire N__22590;
    wire N__22587;
    wire N__22584;
    wire N__22579;
    wire N__22576;
    wire N__22573;
    wire N__22570;
    wire N__22567;
    wire N__22564;
    wire N__22561;
    wire N__22554;
    wire N__22549;
    wire N__22546;
    wire N__22541;
    wire N__22538;
    wire N__22535;
    wire N__22528;
    wire N__22521;
    wire N__22518;
    wire N__22513;
    wire N__22502;
    wire N__22499;
    wire N__22496;
    wire N__22493;
    wire N__22490;
    wire N__22487;
    wire N__22484;
    wire N__22481;
    wire N__22478;
    wire N__22475;
    wire N__22472;
    wire N__22469;
    wire N__22466;
    wire N__22463;
    wire N__22460;
    wire N__22457;
    wire N__22454;
    wire N__22451;
    wire N__22448;
    wire N__22445;
    wire N__22442;
    wire N__22439;
    wire N__22436;
    wire N__22433;
    wire N__22430;
    wire N__22427;
    wire N__22424;
    wire N__22421;
    wire N__22418;
    wire N__22415;
    wire N__22412;
    wire N__22409;
    wire N__22406;
    wire N__22403;
    wire N__22400;
    wire N__22397;
    wire N__22394;
    wire N__22391;
    wire N__22388;
    wire N__22385;
    wire N__22382;
    wire N__22379;
    wire N__22376;
    wire N__22373;
    wire N__22370;
    wire N__22367;
    wire N__22364;
    wire N__22361;
    wire N__22358;
    wire N__22355;
    wire N__22352;
    wire N__22349;
    wire N__22346;
    wire N__22343;
    wire N__22340;
    wire N__22337;
    wire N__22334;
    wire N__22331;
    wire N__22328;
    wire N__22325;
    wire N__22322;
    wire N__22319;
    wire N__22316;
    wire N__22313;
    wire N__22310;
    wire N__22307;
    wire N__22304;
    wire N__22301;
    wire N__22298;
    wire N__22295;
    wire N__22292;
    wire N__22289;
    wire N__22286;
    wire N__22283;
    wire N__22280;
    wire N__22277;
    wire N__22274;
    wire N__22271;
    wire N__22268;
    wire N__22265;
    wire N__22262;
    wire N__22259;
    wire N__22258;
    wire N__22255;
    wire N__22252;
    wire N__22247;
    wire N__22244;
    wire N__22243;
    wire N__22240;
    wire N__22237;
    wire N__22234;
    wire N__22231;
    wire N__22228;
    wire N__22225;
    wire N__22220;
    wire N__22217;
    wire N__22214;
    wire N__22211;
    wire N__22208;
    wire N__22207;
    wire N__22204;
    wire N__22201;
    wire N__22198;
    wire N__22197;
    wire N__22194;
    wire N__22191;
    wire N__22188;
    wire N__22185;
    wire N__22182;
    wire N__22179;
    wire N__22176;
    wire N__22173;
    wire N__22170;
    wire N__22167;
    wire N__22162;
    wire N__22159;
    wire N__22154;
    wire N__22151;
    wire N__22150;
    wire N__22149;
    wire N__22148;
    wire N__22145;
    wire N__22142;
    wire N__22139;
    wire N__22136;
    wire N__22135;
    wire N__22134;
    wire N__22133;
    wire N__22132;
    wire N__22129;
    wire N__22122;
    wire N__22119;
    wire N__22116;
    wire N__22113;
    wire N__22110;
    wire N__22107;
    wire N__22100;
    wire N__22095;
    wire N__22092;
    wire N__22089;
    wire N__22086;
    wire N__22081;
    wire N__22078;
    wire N__22073;
    wire N__22070;
    wire N__22067;
    wire N__22064;
    wire N__22061;
    wire N__22058;
    wire N__22055;
    wire N__22052;
    wire N__22049;
    wire N__22046;
    wire N__22043;
    wire N__22040;
    wire N__22037;
    wire N__22034;
    wire N__22031;
    wire N__22028;
    wire N__22025;
    wire N__22022;
    wire N__22019;
    wire N__22016;
    wire N__22013;
    wire N__22010;
    wire N__22007;
    wire N__22004;
    wire N__22001;
    wire N__21998;
    wire N__21995;
    wire N__21992;
    wire N__21989;
    wire N__21986;
    wire N__21983;
    wire N__21980;
    wire N__21977;
    wire N__21974;
    wire N__21971;
    wire N__21968;
    wire N__21965;
    wire N__21962;
    wire N__21959;
    wire N__21956;
    wire N__21953;
    wire N__21950;
    wire N__21947;
    wire N__21944;
    wire N__21941;
    wire N__21938;
    wire N__21935;
    wire N__21932;
    wire N__21929;
    wire N__21926;
    wire N__21923;
    wire N__21920;
    wire N__21917;
    wire N__21914;
    wire N__21911;
    wire N__21908;
    wire N__21905;
    wire N__21902;
    wire N__21899;
    wire N__21896;
    wire N__21893;
    wire N__21890;
    wire N__21887;
    wire N__21884;
    wire N__21881;
    wire N__21878;
    wire N__21875;
    wire N__21872;
    wire N__21869;
    wire N__21866;
    wire N__21863;
    wire N__21862;
    wire N__21859;
    wire N__21856;
    wire N__21855;
    wire N__21852;
    wire N__21849;
    wire N__21846;
    wire N__21843;
    wire N__21840;
    wire N__21837;
    wire N__21832;
    wire N__21829;
    wire N__21826;
    wire N__21823;
    wire N__21820;
    wire N__21815;
    wire N__21812;
    wire N__21809;
    wire N__21806;
    wire N__21803;
    wire N__21800;
    wire N__21797;
    wire N__21794;
    wire N__21791;
    wire N__21788;
    wire N__21785;
    wire N__21782;
    wire N__21779;
    wire N__21776;
    wire N__21773;
    wire N__21770;
    wire N__21767;
    wire N__21764;
    wire N__21761;
    wire N__21758;
    wire N__21755;
    wire N__21752;
    wire N__21749;
    wire N__21746;
    wire N__21743;
    wire N__21740;
    wire N__21737;
    wire N__21734;
    wire N__21731;
    wire N__21728;
    wire N__21725;
    wire N__21722;
    wire N__21719;
    wire N__21716;
    wire N__21713;
    wire N__21710;
    wire N__21707;
    wire N__21704;
    wire N__21701;
    wire N__21698;
    wire N__21695;
    wire N__21692;
    wire N__21689;
    wire N__21686;
    wire N__21683;
    wire N__21680;
    wire N__21677;
    wire N__21674;
    wire N__21671;
    wire N__21668;
    wire N__21665;
    wire N__21662;
    wire N__21659;
    wire N__21656;
    wire N__21653;
    wire N__21650;
    wire N__21647;
    wire N__21644;
    wire N__21641;
    wire N__21638;
    wire N__21635;
    wire N__21632;
    wire N__21629;
    wire N__21626;
    wire N__21623;
    wire N__21622;
    wire N__21619;
    wire N__21618;
    wire N__21615;
    wire N__21614;
    wire N__21613;
    wire N__21612;
    wire N__21611;
    wire N__21608;
    wire N__21607;
    wire N__21606;
    wire N__21605;
    wire N__21604;
    wire N__21603;
    wire N__21602;
    wire N__21599;
    wire N__21596;
    wire N__21593;
    wire N__21586;
    wire N__21585;
    wire N__21582;
    wire N__21579;
    wire N__21572;
    wire N__21569;
    wire N__21566;
    wire N__21563;
    wire N__21558;
    wire N__21555;
    wire N__21552;
    wire N__21543;
    wire N__21530;
    wire N__21527;
    wire N__21524;
    wire N__21521;
    wire N__21518;
    wire N__21515;
    wire N__21512;
    wire N__21509;
    wire N__21506;
    wire N__21503;
    wire N__21500;
    wire N__21497;
    wire N__21494;
    wire N__21491;
    wire N__21488;
    wire N__21485;
    wire N__21482;
    wire N__21479;
    wire N__21476;
    wire N__21473;
    wire N__21470;
    wire N__21467;
    wire N__21464;
    wire N__21461;
    wire N__21458;
    wire N__21455;
    wire N__21452;
    wire N__21449;
    wire N__21446;
    wire N__21443;
    wire N__21440;
    wire N__21437;
    wire N__21434;
    wire N__21431;
    wire N__21430;
    wire N__21427;
    wire N__21424;
    wire N__21423;
    wire N__21420;
    wire N__21417;
    wire N__21414;
    wire N__21411;
    wire N__21408;
    wire N__21403;
    wire N__21400;
    wire N__21397;
    wire N__21394;
    wire N__21389;
    wire N__21386;
    wire N__21383;
    wire N__21380;
    wire N__21377;
    wire N__21374;
    wire N__21373;
    wire N__21370;
    wire N__21367;
    wire N__21364;
    wire N__21361;
    wire N__21356;
    wire N__21355;
    wire N__21352;
    wire N__21349;
    wire N__21346;
    wire N__21343;
    wire N__21340;
    wire N__21337;
    wire N__21334;
    wire N__21331;
    wire N__21326;
    wire N__21323;
    wire N__21320;
    wire N__21317;
    wire N__21314;
    wire N__21311;
    wire N__21310;
    wire N__21307;
    wire N__21304;
    wire N__21303;
    wire N__21300;
    wire N__21297;
    wire N__21294;
    wire N__21289;
    wire N__21286;
    wire N__21283;
    wire N__21280;
    wire N__21277;
    wire N__21272;
    wire N__21269;
    wire N__21266;
    wire N__21263;
    wire N__21260;
    wire N__21257;
    wire N__21254;
    wire N__21251;
    wire N__21248;
    wire N__21245;
    wire N__21242;
    wire N__21239;
    wire N__21236;
    wire N__21233;
    wire N__21230;
    wire N__21227;
    wire N__21224;
    wire N__21221;
    wire N__21218;
    wire N__21215;
    wire N__21212;
    wire N__21209;
    wire N__21206;
    wire N__21203;
    wire N__21200;
    wire N__21197;
    wire N__21194;
    wire N__21191;
    wire N__21188;
    wire N__21185;
    wire N__21182;
    wire N__21179;
    wire N__21176;
    wire N__21173;
    wire N__21170;
    wire N__21167;
    wire N__21164;
    wire N__21161;
    wire N__21158;
    wire N__21155;
    wire N__21152;
    wire N__21149;
    wire N__21146;
    wire N__21143;
    wire N__21140;
    wire N__21137;
    wire N__21134;
    wire N__21131;
    wire N__21130;
    wire N__21129;
    wire N__21126;
    wire N__21123;
    wire N__21120;
    wire N__21119;
    wire N__21118;
    wire N__21117;
    wire N__21112;
    wire N__21111;
    wire N__21108;
    wire N__21105;
    wire N__21102;
    wire N__21099;
    wire N__21096;
    wire N__21093;
    wire N__21086;
    wire N__21083;
    wire N__21080;
    wire N__21077;
    wire N__21074;
    wire N__21065;
    wire N__21064;
    wire N__21063;
    wire N__21062;
    wire N__21061;
    wire N__21058;
    wire N__21057;
    wire N__21056;
    wire N__21055;
    wire N__21054;
    wire N__21051;
    wire N__21048;
    wire N__21047;
    wire N__21046;
    wire N__21043;
    wire N__21040;
    wire N__21037;
    wire N__21034;
    wire N__21033;
    wire N__21032;
    wire N__21029;
    wire N__21026;
    wire N__21023;
    wire N__21022;
    wire N__21019;
    wire N__21016;
    wire N__21013;
    wire N__21010;
    wire N__21009;
    wire N__21006;
    wire N__21003;
    wire N__21000;
    wire N__20997;
    wire N__20994;
    wire N__20991;
    wire N__20990;
    wire N__20987;
    wire N__20984;
    wire N__20981;
    wire N__20978;
    wire N__20973;
    wire N__20968;
    wire N__20965;
    wire N__20956;
    wire N__20953;
    wire N__20950;
    wire N__20947;
    wire N__20940;
    wire N__20937;
    wire N__20934;
    wire N__20927;
    wire N__20918;
    wire N__20909;
    wire N__20906;
    wire N__20903;
    wire N__20900;
    wire N__20897;
    wire N__20894;
    wire N__20891;
    wire N__20888;
    wire N__20885;
    wire N__20882;
    wire N__20879;
    wire N__20878;
    wire N__20877;
    wire N__20876;
    wire N__20875;
    wire N__20872;
    wire N__20871;
    wire N__20870;
    wire N__20869;
    wire N__20868;
    wire N__20865;
    wire N__20862;
    wire N__20859;
    wire N__20856;
    wire N__20855;
    wire N__20850;
    wire N__20845;
    wire N__20842;
    wire N__20841;
    wire N__20840;
    wire N__20839;
    wire N__20836;
    wire N__20833;
    wire N__20830;
    wire N__20825;
    wire N__20824;
    wire N__20823;
    wire N__20822;
    wire N__20821;
    wire N__20820;
    wire N__20819;
    wire N__20818;
    wire N__20817;
    wire N__20812;
    wire N__20809;
    wire N__20806;
    wire N__20801;
    wire N__20798;
    wire N__20793;
    wire N__20790;
    wire N__20787;
    wire N__20782;
    wire N__20773;
    wire N__20772;
    wire N__20771;
    wire N__20770;
    wire N__20769;
    wire N__20766;
    wire N__20765;
    wire N__20764;
    wire N__20763;
    wire N__20756;
    wire N__20753;
    wire N__20748;
    wire N__20743;
    wire N__20738;
    wire N__20731;
    wire N__20728;
    wire N__20725;
    wire N__20720;
    wire N__20717;
    wire N__20712;
    wire N__20709;
    wire N__20704;
    wire N__20687;
    wire N__20684;
    wire N__20681;
    wire N__20678;
    wire N__20675;
    wire N__20672;
    wire N__20669;
    wire N__20666;
    wire N__20663;
    wire N__20660;
    wire N__20657;
    wire N__20656;
    wire N__20655;
    wire N__20654;
    wire N__20653;
    wire N__20652;
    wire N__20649;
    wire N__20646;
    wire N__20643;
    wire N__20636;
    wire N__20635;
    wire N__20634;
    wire N__20631;
    wire N__20628;
    wire N__20625;
    wire N__20622;
    wire N__20621;
    wire N__20620;
    wire N__20617;
    wire N__20614;
    wire N__20613;
    wire N__20612;
    wire N__20611;
    wire N__20610;
    wire N__20607;
    wire N__20604;
    wire N__20601;
    wire N__20598;
    wire N__20595;
    wire N__20592;
    wire N__20587;
    wire N__20584;
    wire N__20577;
    wire N__20558;
    wire N__20557;
    wire N__20554;
    wire N__20551;
    wire N__20548;
    wire N__20545;
    wire N__20542;
    wire N__20539;
    wire N__20536;
    wire N__20533;
    wire N__20528;
    wire N__20525;
    wire N__20524;
    wire N__20523;
    wire N__20520;
    wire N__20517;
    wire N__20516;
    wire N__20513;
    wire N__20508;
    wire N__20505;
    wire N__20502;
    wire N__20499;
    wire N__20496;
    wire N__20493;
    wire N__20486;
    wire N__20483;
    wire N__20480;
    wire N__20479;
    wire N__20476;
    wire N__20473;
    wire N__20472;
    wire N__20469;
    wire N__20466;
    wire N__20463;
    wire N__20456;
    wire N__20455;
    wire N__20454;
    wire N__20451;
    wire N__20448;
    wire N__20445;
    wire N__20444;
    wire N__20439;
    wire N__20436;
    wire N__20433;
    wire N__20430;
    wire N__20425;
    wire N__20420;
    wire N__20417;
    wire N__20416;
    wire N__20415;
    wire N__20414;
    wire N__20413;
    wire N__20410;
    wire N__20409;
    wire N__20408;
    wire N__20407;
    wire N__20404;
    wire N__20401;
    wire N__20398;
    wire N__20397;
    wire N__20394;
    wire N__20393;
    wire N__20392;
    wire N__20389;
    wire N__20386;
    wire N__20385;
    wire N__20384;
    wire N__20381;
    wire N__20378;
    wire N__20375;
    wire N__20372;
    wire N__20369;
    wire N__20366;
    wire N__20363;
    wire N__20360;
    wire N__20357;
    wire N__20356;
    wire N__20355;
    wire N__20354;
    wire N__20353;
    wire N__20352;
    wire N__20349;
    wire N__20346;
    wire N__20343;
    wire N__20340;
    wire N__20339;
    wire N__20338;
    wire N__20337;
    wire N__20336;
    wire N__20335;
    wire N__20332;
    wire N__20329;
    wire N__20328;
    wire N__20327;
    wire N__20326;
    wire N__20321;
    wire N__20316;
    wire N__20309;
    wire N__20306;
    wire N__20305;
    wire N__20302;
    wire N__20299;
    wire N__20298;
    wire N__20297;
    wire N__20296;
    wire N__20295;
    wire N__20294;
    wire N__20293;
    wire N__20292;
    wire N__20289;
    wire N__20288;
    wire N__20287;
    wire N__20286;
    wire N__20285;
    wire N__20284;
    wire N__20281;
    wire N__20272;
    wire N__20269;
    wire N__20268;
    wire N__20267;
    wire N__20264;
    wire N__20261;
    wire N__20260;
    wire N__20259;
    wire N__20258;
    wire N__20255;
    wire N__20252;
    wire N__20251;
    wire N__20250;
    wire N__20247;
    wire N__20244;
    wire N__20241;
    wire N__20240;
    wire N__20239;
    wire N__20238;
    wire N__20237;
    wire N__20236;
    wire N__20233;
    wire N__20230;
    wire N__20229;
    wire N__20220;
    wire N__20217;
    wire N__20214;
    wire N__20211;
    wire N__20208;
    wire N__20205;
    wire N__20202;
    wire N__20199;
    wire N__20196;
    wire N__20193;
    wire N__20190;
    wire N__20189;
    wire N__20188;
    wire N__20187;
    wire N__20186;
    wire N__20183;
    wire N__20180;
    wire N__20179;
    wire N__20176;
    wire N__20173;
    wire N__20172;
    wire N__20171;
    wire N__20170;
    wire N__20169;
    wire N__20168;
    wire N__20165;
    wire N__20164;
    wire N__20163;
    wire N__20160;
    wire N__20157;
    wire N__20152;
    wire N__20149;
    wire N__20146;
    wire N__20141;
    wire N__20138;
    wire N__20135;
    wire N__20132;
    wire N__20127;
    wire N__20124;
    wire N__20123;
    wire N__20122;
    wire N__20121;
    wire N__20118;
    wire N__20113;
    wire N__20110;
    wire N__20107;
    wire N__20104;
    wire N__20101;
    wire N__20096;
    wire N__20093;
    wire N__20090;
    wire N__20087;
    wire N__20080;
    wire N__20075;
    wire N__20070;
    wire N__20061;
    wire N__20058;
    wire N__20055;
    wire N__20052;
    wire N__20049;
    wire N__20046;
    wire N__20043;
    wire N__20038;
    wire N__20029;
    wire N__20026;
    wire N__20023;
    wire N__20020;
    wire N__20017;
    wire N__20016;
    wire N__20015;
    wire N__20012;
    wire N__20007;
    wire N__20002;
    wire N__19995;
    wire N__19992;
    wire N__19989;
    wire N__19984;
    wire N__19981;
    wire N__19978;
    wire N__19975;
    wire N__19972;
    wire N__19969;
    wire N__19966;
    wire N__19963;
    wire N__19956;
    wire N__19951;
    wire N__19946;
    wire N__19939;
    wire N__19936;
    wire N__19931;
    wire N__19920;
    wire N__19915;
    wire N__19910;
    wire N__19907;
    wire N__19902;
    wire N__19895;
    wire N__19890;
    wire N__19885;
    wire N__19882;
    wire N__19879;
    wire N__19872;
    wire N__19863;
    wire N__19854;
    wire N__19845;
    wire N__19826;
    wire N__19823;
    wire N__19820;
    wire N__19817;
    wire N__19814;
    wire N__19811;
    wire N__19808;
    wire N__19805;
    wire N__19802;
    wire N__19799;
    wire N__19796;
    wire N__19793;
    wire N__19790;
    wire N__19787;
    wire N__19784;
    wire N__19781;
    wire N__19778;
    wire N__19777;
    wire N__19774;
    wire N__19771;
    wire N__19770;
    wire N__19767;
    wire N__19766;
    wire N__19765;
    wire N__19762;
    wire N__19759;
    wire N__19756;
    wire N__19755;
    wire N__19752;
    wire N__19749;
    wire N__19748;
    wire N__19743;
    wire N__19742;
    wire N__19739;
    wire N__19736;
    wire N__19733;
    wire N__19730;
    wire N__19727;
    wire N__19724;
    wire N__19721;
    wire N__19718;
    wire N__19715;
    wire N__19712;
    wire N__19707;
    wire N__19702;
    wire N__19697;
    wire N__19692;
    wire N__19689;
    wire N__19686;
    wire N__19683;
    wire N__19680;
    wire N__19673;
    wire N__19672;
    wire N__19669;
    wire N__19666;
    wire N__19663;
    wire N__19658;
    wire N__19655;
    wire N__19652;
    wire N__19649;
    wire N__19646;
    wire N__19643;
    wire N__19640;
    wire N__19637;
    wire N__19634;
    wire N__19631;
    wire N__19628;
    wire N__19625;
    wire N__19622;
    wire N__19619;
    wire N__19616;
    wire N__19613;
    wire N__19610;
    wire N__19607;
    wire N__19604;
    wire N__19601;
    wire N__19598;
    wire N__19595;
    wire N__19592;
    wire N__19591;
    wire N__19588;
    wire N__19585;
    wire N__19580;
    wire N__19577;
    wire N__19576;
    wire N__19573;
    wire N__19570;
    wire N__19565;
    wire N__19564;
    wire N__19561;
    wire N__19558;
    wire N__19555;
    wire N__19552;
    wire N__19549;
    wire N__19546;
    wire N__19543;
    wire N__19540;
    wire N__19537;
    wire N__19534;
    wire N__19531;
    wire N__19528;
    wire N__19525;
    wire N__19522;
    wire N__19519;
    wire N__19516;
    wire N__19513;
    wire N__19510;
    wire N__19507;
    wire N__19504;
    wire N__19501;
    wire N__19498;
    wire N__19495;
    wire N__19492;
    wire N__19489;
    wire N__19486;
    wire N__19483;
    wire N__19480;
    wire N__19477;
    wire N__19474;
    wire N__19471;
    wire N__19468;
    wire N__19465;
    wire N__19462;
    wire N__19459;
    wire N__19456;
    wire N__19453;
    wire N__19450;
    wire N__19447;
    wire N__19444;
    wire N__19441;
    wire N__19438;
    wire N__19435;
    wire N__19432;
    wire N__19429;
    wire N__19426;
    wire N__19423;
    wire N__19420;
    wire N__19417;
    wire N__19414;
    wire N__19411;
    wire N__19408;
    wire N__19405;
    wire N__19402;
    wire N__19399;
    wire N__19396;
    wire N__19393;
    wire N__19390;
    wire N__19387;
    wire N__19384;
    wire N__19381;
    wire N__19378;
    wire N__19375;
    wire N__19372;
    wire N__19369;
    wire N__19366;
    wire N__19363;
    wire N__19360;
    wire N__19357;
    wire N__19354;
    wire N__19351;
    wire N__19346;
    wire N__19343;
    wire N__19340;
    wire N__19337;
    wire N__19334;
    wire N__19333;
    wire N__19332;
    wire N__19329;
    wire N__19328;
    wire N__19325;
    wire N__19322;
    wire N__19319;
    wire N__19316;
    wire N__19311;
    wire N__19308;
    wire N__19305;
    wire N__19298;
    wire N__19295;
    wire N__19294;
    wire N__19291;
    wire N__19288;
    wire N__19283;
    wire N__19280;
    wire N__19277;
    wire N__19274;
    wire N__19273;
    wire N__19272;
    wire N__19269;
    wire N__19266;
    wire N__19263;
    wire N__19262;
    wire N__19255;
    wire N__19252;
    wire N__19249;
    wire N__19246;
    wire N__19241;
    wire N__19238;
    wire N__19237;
    wire N__19234;
    wire N__19231;
    wire N__19226;
    wire N__19223;
    wire N__19220;
    wire N__19217;
    wire N__19216;
    wire N__19215;
    wire N__19212;
    wire N__19209;
    wire N__19208;
    wire N__19205;
    wire N__19200;
    wire N__19197;
    wire N__19194;
    wire N__19187;
    wire N__19184;
    wire N__19181;
    wire N__19178;
    wire N__19177;
    wire N__19174;
    wire N__19171;
    wire N__19170;
    wire N__19169;
    wire N__19164;
    wire N__19161;
    wire N__19158;
    wire N__19155;
    wire N__19152;
    wire N__19149;
    wire N__19142;
    wire N__19139;
    wire N__19136;
    wire N__19133;
    wire N__19130;
    wire N__19127;
    wire N__19124;
    wire N__19123;
    wire N__19120;
    wire N__19117;
    wire N__19112;
    wire N__19109;
    wire N__19108;
    wire N__19105;
    wire N__19102;
    wire N__19099;
    wire N__19096;
    wire N__19093;
    wire N__19090;
    wire N__19087;
    wire N__19084;
    wire N__19081;
    wire N__19078;
    wire N__19075;
    wire N__19072;
    wire N__19069;
    wire N__19066;
    wire N__19063;
    wire N__19060;
    wire N__19057;
    wire N__19054;
    wire N__19051;
    wire N__19048;
    wire N__19045;
    wire N__19042;
    wire N__19039;
    wire N__19036;
    wire N__19033;
    wire N__19030;
    wire N__19027;
    wire N__19024;
    wire N__19021;
    wire N__19018;
    wire N__19015;
    wire N__19012;
    wire N__19009;
    wire N__19006;
    wire N__19003;
    wire N__19000;
    wire N__18997;
    wire N__18994;
    wire N__18991;
    wire N__18988;
    wire N__18985;
    wire N__18982;
    wire N__18979;
    wire N__18976;
    wire N__18973;
    wire N__18970;
    wire N__18967;
    wire N__18964;
    wire N__18961;
    wire N__18958;
    wire N__18955;
    wire N__18952;
    wire N__18949;
    wire N__18946;
    wire N__18943;
    wire N__18940;
    wire N__18937;
    wire N__18934;
    wire N__18931;
    wire N__18928;
    wire N__18925;
    wire N__18922;
    wire N__18919;
    wire N__18916;
    wire N__18913;
    wire N__18910;
    wire N__18907;
    wire N__18904;
    wire N__18901;
    wire N__18898;
    wire N__18895;
    wire N__18890;
    wire N__18889;
    wire N__18886;
    wire N__18883;
    wire N__18880;
    wire N__18877;
    wire N__18874;
    wire N__18869;
    wire N__18866;
    wire N__18863;
    wire N__18860;
    wire N__18857;
    wire N__18854;
    wire N__18853;
    wire N__18850;
    wire N__18847;
    wire N__18844;
    wire N__18841;
    wire N__18838;
    wire N__18835;
    wire N__18832;
    wire N__18829;
    wire N__18826;
    wire N__18823;
    wire N__18820;
    wire N__18817;
    wire N__18814;
    wire N__18811;
    wire N__18808;
    wire N__18805;
    wire N__18802;
    wire N__18799;
    wire N__18796;
    wire N__18793;
    wire N__18790;
    wire N__18787;
    wire N__18784;
    wire N__18781;
    wire N__18778;
    wire N__18775;
    wire N__18772;
    wire N__18769;
    wire N__18766;
    wire N__18763;
    wire N__18760;
    wire N__18757;
    wire N__18754;
    wire N__18751;
    wire N__18748;
    wire N__18745;
    wire N__18742;
    wire N__18739;
    wire N__18736;
    wire N__18733;
    wire N__18730;
    wire N__18727;
    wire N__18724;
    wire N__18721;
    wire N__18718;
    wire N__18715;
    wire N__18712;
    wire N__18709;
    wire N__18706;
    wire N__18703;
    wire N__18700;
    wire N__18697;
    wire N__18694;
    wire N__18691;
    wire N__18688;
    wire N__18685;
    wire N__18682;
    wire N__18679;
    wire N__18676;
    wire N__18673;
    wire N__18670;
    wire N__18667;
    wire N__18664;
    wire N__18661;
    wire N__18658;
    wire N__18655;
    wire N__18652;
    wire N__18649;
    wire N__18644;
    wire N__18641;
    wire N__18638;
    wire N__18635;
    wire N__18632;
    wire N__18629;
    wire N__18626;
    wire N__18623;
    wire N__18620;
    wire N__18617;
    wire N__18614;
    wire N__18611;
    wire N__18608;
    wire N__18605;
    wire N__18602;
    wire N__18599;
    wire N__18596;
    wire N__18593;
    wire N__18590;
    wire N__18587;
    wire N__18584;
    wire N__18581;
    wire N__18578;
    wire N__18575;
    wire N__18572;
    wire N__18569;
    wire N__18568;
    wire N__18565;
    wire N__18562;
    wire N__18561;
    wire N__18560;
    wire N__18559;
    wire N__18558;
    wire N__18553;
    wire N__18550;
    wire N__18547;
    wire N__18544;
    wire N__18541;
    wire N__18540;
    wire N__18533;
    wire N__18532;
    wire N__18529;
    wire N__18526;
    wire N__18523;
    wire N__18520;
    wire N__18517;
    wire N__18514;
    wire N__18509;
    wire N__18504;
    wire N__18501;
    wire N__18498;
    wire N__18495;
    wire N__18492;
    wire N__18489;
    wire N__18486;
    wire N__18483;
    wire N__18480;
    wire N__18477;
    wire N__18470;
    wire N__18467;
    wire N__18464;
    wire N__18461;
    wire N__18458;
    wire N__18455;
    wire N__18454;
    wire N__18451;
    wire N__18448;
    wire N__18445;
    wire N__18442;
    wire N__18437;
    wire N__18434;
    wire N__18431;
    wire N__18428;
    wire N__18425;
    wire N__18422;
    wire N__18419;
    wire N__18418;
    wire N__18415;
    wire N__18412;
    wire N__18407;
    wire N__18406;
    wire N__18403;
    wire N__18402;
    wire N__18399;
    wire N__18396;
    wire N__18393;
    wire N__18392;
    wire N__18391;
    wire N__18388;
    wire N__18383;
    wire N__18382;
    wire N__18379;
    wire N__18376;
    wire N__18371;
    wire N__18368;
    wire N__18365;
    wire N__18362;
    wire N__18357;
    wire N__18354;
    wire N__18349;
    wire N__18346;
    wire N__18343;
    wire N__18338;
    wire N__18335;
    wire N__18332;
    wire N__18331;
    wire N__18328;
    wire N__18325;
    wire N__18320;
    wire N__18317;
    wire N__18314;
    wire N__18311;
    wire N__18308;
    wire N__18305;
    wire N__18302;
    wire N__18299;
    wire N__18296;
    wire N__18295;
    wire N__18292;
    wire N__18289;
    wire N__18288;
    wire N__18283;
    wire N__18282;
    wire N__18279;
    wire N__18276;
    wire N__18273;
    wire N__18270;
    wire N__18263;
    wire N__18260;
    wire N__18257;
    wire N__18254;
    wire N__18251;
    wire N__18248;
    wire N__18245;
    wire N__18242;
    wire N__18239;
    wire N__18238;
    wire N__18235;
    wire N__18232;
    wire N__18229;
    wire N__18226;
    wire N__18223;
    wire N__18218;
    wire N__18217;
    wire N__18214;
    wire N__18213;
    wire N__18212;
    wire N__18209;
    wire N__18208;
    wire N__18207;
    wire N__18204;
    wire N__18201;
    wire N__18198;
    wire N__18197;
    wire N__18196;
    wire N__18193;
    wire N__18190;
    wire N__18187;
    wire N__18186;
    wire N__18185;
    wire N__18178;
    wire N__18175;
    wire N__18172;
    wire N__18171;
    wire N__18170;
    wire N__18163;
    wire N__18160;
    wire N__18157;
    wire N__18156;
    wire N__18155;
    wire N__18148;
    wire N__18145;
    wire N__18142;
    wire N__18141;
    wire N__18140;
    wire N__18133;
    wire N__18130;
    wire N__18127;
    wire N__18126;
    wire N__18125;
    wire N__18124;
    wire N__18117;
    wire N__18114;
    wire N__18111;
    wire N__18110;
    wire N__18109;
    wire N__18102;
    wire N__18099;
    wire N__18096;
    wire N__18095;
    wire N__18094;
    wire N__18093;
    wire N__18090;
    wire N__18089;
    wire N__18088;
    wire N__18085;
    wire N__18080;
    wire N__18077;
    wire N__18074;
    wire N__18073;
    wire N__18072;
    wire N__18071;
    wire N__18070;
    wire N__18063;
    wire N__18060;
    wire N__18057;
    wire N__18054;
    wire N__18053;
    wire N__18052;
    wire N__18051;
    wire N__18050;
    wire N__18047;
    wire N__18044;
    wire N__18041;
    wire N__18038;
    wire N__18031;
    wire N__18028;
    wire N__18025;
    wire N__18022;
    wire N__18019;
    wire N__18012;
    wire N__18009;
    wire N__18006;
    wire N__18003;
    wire N__18000;
    wire N__17997;
    wire N__17990;
    wire N__17981;
    wire N__17976;
    wire N__17973;
    wire N__17966;
    wire N__17961;
    wire N__17956;
    wire N__17953;
    wire N__17950;
    wire N__17945;
    wire N__17942;
    wire N__17939;
    wire N__17934;
    wire N__17929;
    wire N__17924;
    wire N__17921;
    wire N__17920;
    wire N__17917;
    wire N__17914;
    wire N__17913;
    wire N__17912;
    wire N__17911;
    wire N__17908;
    wire N__17905;
    wire N__17902;
    wire N__17899;
    wire N__17896;
    wire N__17893;
    wire N__17892;
    wire N__17887;
    wire N__17886;
    wire N__17883;
    wire N__17882;
    wire N__17879;
    wire N__17876;
    wire N__17873;
    wire N__17870;
    wire N__17867;
    wire N__17864;
    wire N__17861;
    wire N__17858;
    wire N__17855;
    wire N__17852;
    wire N__17847;
    wire N__17842;
    wire N__17839;
    wire N__17834;
    wire N__17831;
    wire N__17828;
    wire N__17821;
    wire N__17818;
    wire N__17813;
    wire N__17810;
    wire N__17807;
    wire N__17804;
    wire N__17801;
    wire N__17798;
    wire N__17795;
    wire N__17792;
    wire N__17789;
    wire N__17788;
    wire N__17785;
    wire N__17782;
    wire N__17779;
    wire N__17776;
    wire N__17775;
    wire N__17774;
    wire N__17771;
    wire N__17770;
    wire N__17769;
    wire N__17766;
    wire N__17763;
    wire N__17762;
    wire N__17761;
    wire N__17758;
    wire N__17755;
    wire N__17752;
    wire N__17749;
    wire N__17744;
    wire N__17741;
    wire N__17738;
    wire N__17735;
    wire N__17732;
    wire N__17729;
    wire N__17726;
    wire N__17719;
    wire N__17716;
    wire N__17713;
    wire N__17708;
    wire N__17705;
    wire N__17702;
    wire N__17693;
    wire N__17690;
    wire N__17687;
    wire N__17684;
    wire N__17681;
    wire N__17678;
    wire N__17677;
    wire N__17674;
    wire N__17673;
    wire N__17672;
    wire N__17671;
    wire N__17668;
    wire N__17665;
    wire N__17662;
    wire N__17659;
    wire N__17658;
    wire N__17655;
    wire N__17654;
    wire N__17651;
    wire N__17646;
    wire N__17645;
    wire N__17642;
    wire N__17639;
    wire N__17636;
    wire N__17633;
    wire N__17630;
    wire N__17627;
    wire N__17624;
    wire N__17621;
    wire N__17618;
    wire N__17615;
    wire N__17612;
    wire N__17605;
    wire N__17600;
    wire N__17597;
    wire N__17594;
    wire N__17591;
    wire N__17584;
    wire N__17581;
    wire N__17576;
    wire N__17573;
    wire N__17570;
    wire N__17567;
    wire N__17564;
    wire N__17561;
    wire N__17558;
    wire N__17555;
    wire N__17552;
    wire N__17549;
    wire N__17546;
    wire N__17543;
    wire N__17540;
    wire N__17537;
    wire N__17534;
    wire N__17531;
    wire N__17528;
    wire N__17525;
    wire N__17522;
    wire N__17519;
    wire N__17516;
    wire N__17513;
    wire N__17510;
    wire N__17509;
    wire N__17506;
    wire N__17503;
    wire N__17500;
    wire N__17497;
    wire N__17494;
    wire N__17491;
    wire N__17488;
    wire N__17485;
    wire N__17482;
    wire N__17479;
    wire N__17476;
    wire N__17473;
    wire N__17470;
    wire N__17467;
    wire N__17464;
    wire N__17461;
    wire N__17458;
    wire N__17455;
    wire N__17452;
    wire N__17449;
    wire N__17446;
    wire N__17443;
    wire N__17440;
    wire N__17437;
    wire N__17434;
    wire N__17431;
    wire N__17428;
    wire N__17425;
    wire N__17422;
    wire N__17419;
    wire N__17416;
    wire N__17413;
    wire N__17410;
    wire N__17407;
    wire N__17404;
    wire N__17401;
    wire N__17398;
    wire N__17395;
    wire N__17392;
    wire N__17389;
    wire N__17386;
    wire N__17383;
    wire N__17380;
    wire N__17377;
    wire N__17374;
    wire N__17371;
    wire N__17368;
    wire N__17365;
    wire N__17362;
    wire N__17359;
    wire N__17356;
    wire N__17353;
    wire N__17350;
    wire N__17347;
    wire N__17344;
    wire N__17341;
    wire N__17338;
    wire N__17335;
    wire N__17332;
    wire N__17329;
    wire N__17326;
    wire N__17323;
    wire N__17320;
    wire N__17317;
    wire N__17314;
    wire N__17311;
    wire N__17308;
    wire N__17305;
    wire N__17302;
    wire N__17299;
    wire N__17296;
    wire N__17293;
    wire N__17288;
    wire N__17285;
    wire N__17282;
    wire N__17279;
    wire N__17276;
    wire N__17273;
    wire N__17272;
    wire N__17271;
    wire N__17268;
    wire N__17265;
    wire N__17264;
    wire N__17261;
    wire N__17256;
    wire N__17251;
    wire N__17246;
    wire N__17245;
    wire N__17242;
    wire N__17239;
    wire N__17236;
    wire N__17233;
    wire N__17230;
    wire N__17227;
    wire N__17224;
    wire N__17221;
    wire N__17218;
    wire N__17215;
    wire N__17212;
    wire N__17209;
    wire N__17206;
    wire N__17203;
    wire N__17200;
    wire N__17197;
    wire N__17194;
    wire N__17191;
    wire N__17188;
    wire N__17185;
    wire N__17182;
    wire N__17179;
    wire N__17176;
    wire N__17173;
    wire N__17170;
    wire N__17167;
    wire N__17164;
    wire N__17161;
    wire N__17158;
    wire N__17155;
    wire N__17152;
    wire N__17149;
    wire N__17146;
    wire N__17143;
    wire N__17140;
    wire N__17137;
    wire N__17134;
    wire N__17131;
    wire N__17128;
    wire N__17125;
    wire N__17122;
    wire N__17119;
    wire N__17116;
    wire N__17113;
    wire N__17110;
    wire N__17107;
    wire N__17104;
    wire N__17101;
    wire N__17098;
    wire N__17095;
    wire N__17092;
    wire N__17089;
    wire N__17086;
    wire N__17083;
    wire N__17080;
    wire N__17077;
    wire N__17074;
    wire N__17071;
    wire N__17068;
    wire N__17065;
    wire N__17062;
    wire N__17059;
    wire N__17056;
    wire N__17053;
    wire N__17050;
    wire N__17047;
    wire N__17044;
    wire N__17041;
    wire N__17038;
    wire N__17035;
    wire N__17030;
    wire N__17027;
    wire N__17024;
    wire N__17021;
    wire N__17020;
    wire N__17017;
    wire N__17016;
    wire N__17015;
    wire N__17012;
    wire N__17009;
    wire N__17006;
    wire N__17003;
    wire N__17000;
    wire N__16991;
    wire N__16988;
    wire N__16985;
    wire N__16982;
    wire N__16979;
    wire N__16976;
    wire N__16973;
    wire N__16972;
    wire N__16969;
    wire N__16966;
    wire N__16963;
    wire N__16960;
    wire N__16957;
    wire N__16954;
    wire N__16951;
    wire N__16948;
    wire N__16945;
    wire N__16942;
    wire N__16939;
    wire N__16936;
    wire N__16933;
    wire N__16930;
    wire N__16927;
    wire N__16924;
    wire N__16921;
    wire N__16918;
    wire N__16915;
    wire N__16912;
    wire N__16909;
    wire N__16906;
    wire N__16903;
    wire N__16900;
    wire N__16897;
    wire N__16894;
    wire N__16891;
    wire N__16888;
    wire N__16885;
    wire N__16882;
    wire N__16879;
    wire N__16876;
    wire N__16873;
    wire N__16870;
    wire N__16867;
    wire N__16864;
    wire N__16861;
    wire N__16858;
    wire N__16855;
    wire N__16852;
    wire N__16849;
    wire N__16846;
    wire N__16843;
    wire N__16840;
    wire N__16837;
    wire N__16834;
    wire N__16831;
    wire N__16828;
    wire N__16825;
    wire N__16822;
    wire N__16819;
    wire N__16816;
    wire N__16813;
    wire N__16810;
    wire N__16807;
    wire N__16804;
    wire N__16801;
    wire N__16798;
    wire N__16795;
    wire N__16792;
    wire N__16789;
    wire N__16786;
    wire N__16783;
    wire N__16780;
    wire N__16777;
    wire N__16774;
    wire N__16771;
    wire N__16768;
    wire N__16765;
    wire N__16762;
    wire N__16759;
    wire N__16756;
    wire N__16753;
    wire N__16750;
    wire N__16745;
    wire N__16742;
    wire N__16739;
    wire N__16736;
    wire N__16735;
    wire N__16732;
    wire N__16729;
    wire N__16726;
    wire N__16721;
    wire N__16718;
    wire N__16717;
    wire N__16716;
    wire N__16713;
    wire N__16712;
    wire N__16711;
    wire N__16708;
    wire N__16705;
    wire N__16702;
    wire N__16697;
    wire N__16694;
    wire N__16685;
    wire N__16682;
    wire N__16679;
    wire N__16676;
    wire N__16673;
    wire N__16670;
    wire N__16667;
    wire N__16666;
    wire N__16665;
    wire N__16664;
    wire N__16661;
    wire N__16658;
    wire N__16655;
    wire N__16652;
    wire N__16643;
    wire N__16642;
    wire N__16639;
    wire N__16636;
    wire N__16633;
    wire N__16628;
    wire N__16625;
    wire N__16622;
    wire N__16619;
    wire N__16616;
    wire N__16613;
    wire N__16610;
    wire N__16607;
    wire N__16604;
    wire N__16601;
    wire N__16598;
    wire N__16595;
    wire N__16592;
    wire N__16589;
    wire N__16586;
    wire N__16583;
    wire N__16580;
    wire N__16577;
    wire N__16576;
    wire N__16573;
    wire N__16570;
    wire N__16567;
    wire N__16564;
    wire N__16559;
    wire N__16556;
    wire N__16553;
    wire N__16552;
    wire N__16551;
    wire N__16548;
    wire N__16545;
    wire N__16544;
    wire N__16541;
    wire N__16536;
    wire N__16533;
    wire N__16526;
    wire N__16523;
    wire N__16520;
    wire N__16517;
    wire N__16514;
    wire N__16511;
    wire N__16508;
    wire N__16505;
    wire N__16502;
    wire N__16501;
    wire N__16498;
    wire N__16495;
    wire N__16494;
    wire N__16493;
    wire N__16488;
    wire N__16485;
    wire N__16482;
    wire N__16477;
    wire N__16474;
    wire N__16469;
    wire N__16466;
    wire N__16463;
    wire N__16460;
    wire N__16457;
    wire N__16454;
    wire N__16451;
    wire N__16448;
    wire N__16445;
    wire N__16442;
    wire N__16439;
    wire N__16436;
    wire N__16433;
    wire N__16430;
    wire N__16427;
    wire N__16424;
    wire N__16423;
    wire N__16422;
    wire N__16421;
    wire N__16418;
    wire N__16415;
    wire N__16410;
    wire N__16403;
    wire N__16400;
    wire N__16399;
    wire N__16398;
    wire N__16397;
    wire N__16394;
    wire N__16391;
    wire N__16386;
    wire N__16379;
    wire N__16376;
    wire N__16373;
    wire N__16370;
    wire N__16369;
    wire N__16366;
    wire N__16363;
    wire N__16362;
    wire N__16361;
    wire N__16360;
    wire N__16359;
    wire N__16356;
    wire N__16353;
    wire N__16348;
    wire N__16343;
    wire N__16334;
    wire N__16331;
    wire N__16328;
    wire N__16325;
    wire N__16322;
    wire N__16321;
    wire N__16318;
    wire N__16315;
    wire N__16312;
    wire N__16309;
    wire N__16306;
    wire N__16303;
    wire N__16300;
    wire N__16297;
    wire N__16294;
    wire N__16291;
    wire N__16288;
    wire N__16285;
    wire N__16282;
    wire N__16279;
    wire N__16276;
    wire N__16273;
    wire N__16270;
    wire N__16267;
    wire N__16264;
    wire N__16261;
    wire N__16258;
    wire N__16255;
    wire N__16252;
    wire N__16249;
    wire N__16246;
    wire N__16243;
    wire N__16240;
    wire N__16237;
    wire N__16234;
    wire N__16231;
    wire N__16228;
    wire N__16225;
    wire N__16222;
    wire N__16219;
    wire N__16216;
    wire N__16213;
    wire N__16210;
    wire N__16207;
    wire N__16204;
    wire N__16201;
    wire N__16198;
    wire N__16195;
    wire N__16192;
    wire N__16189;
    wire N__16186;
    wire N__16183;
    wire N__16180;
    wire N__16177;
    wire N__16174;
    wire N__16171;
    wire N__16168;
    wire N__16165;
    wire N__16162;
    wire N__16159;
    wire N__16156;
    wire N__16153;
    wire N__16150;
    wire N__16147;
    wire N__16144;
    wire N__16141;
    wire N__16138;
    wire N__16135;
    wire N__16132;
    wire N__16129;
    wire N__16126;
    wire N__16123;
    wire N__16120;
    wire N__16117;
    wire N__16114;
    wire N__16111;
    wire N__16108;
    wire N__16105;
    wire N__16100;
    wire N__16097;
    wire N__16094;
    wire N__16093;
    wire N__16090;
    wire N__16087;
    wire N__16082;
    wire N__16081;
    wire N__16078;
    wire N__16075;
    wire N__16072;
    wire N__16067;
    wire N__16066;
    wire N__16063;
    wire N__16060;
    wire N__16057;
    wire N__16054;
    wire N__16051;
    wire N__16048;
    wire N__16045;
    wire N__16042;
    wire N__16039;
    wire N__16036;
    wire N__16033;
    wire N__16030;
    wire N__16027;
    wire N__16024;
    wire N__16021;
    wire N__16018;
    wire N__16015;
    wire N__16012;
    wire N__16009;
    wire N__16006;
    wire N__16003;
    wire N__16000;
    wire N__15997;
    wire N__15994;
    wire N__15991;
    wire N__15988;
    wire N__15985;
    wire N__15982;
    wire N__15979;
    wire N__15976;
    wire N__15973;
    wire N__15970;
    wire N__15967;
    wire N__15964;
    wire N__15961;
    wire N__15958;
    wire N__15955;
    wire N__15952;
    wire N__15949;
    wire N__15946;
    wire N__15943;
    wire N__15940;
    wire N__15937;
    wire N__15934;
    wire N__15931;
    wire N__15928;
    wire N__15925;
    wire N__15922;
    wire N__15919;
    wire N__15916;
    wire N__15913;
    wire N__15910;
    wire N__15907;
    wire N__15904;
    wire N__15901;
    wire N__15898;
    wire N__15895;
    wire N__15892;
    wire N__15889;
    wire N__15886;
    wire N__15883;
    wire N__15880;
    wire N__15877;
    wire N__15874;
    wire N__15871;
    wire N__15868;
    wire N__15865;
    wire N__15862;
    wire N__15859;
    wire N__15854;
    wire N__15851;
    wire N__15850;
    wire N__15847;
    wire N__15844;
    wire N__15841;
    wire N__15838;
    wire N__15833;
    wire N__15830;
    wire N__15827;
    wire N__15826;
    wire N__15823;
    wire N__15820;
    wire N__15817;
    wire N__15812;
    wire N__15811;
    wire N__15808;
    wire N__15805;
    wire N__15802;
    wire N__15799;
    wire N__15796;
    wire N__15793;
    wire N__15790;
    wire N__15787;
    wire N__15784;
    wire N__15781;
    wire N__15778;
    wire N__15775;
    wire N__15772;
    wire N__15769;
    wire N__15766;
    wire N__15763;
    wire N__15760;
    wire N__15757;
    wire N__15754;
    wire N__15751;
    wire N__15748;
    wire N__15745;
    wire N__15742;
    wire N__15739;
    wire N__15736;
    wire N__15733;
    wire N__15730;
    wire N__15727;
    wire N__15724;
    wire N__15721;
    wire N__15718;
    wire N__15715;
    wire N__15712;
    wire N__15709;
    wire N__15706;
    wire N__15703;
    wire N__15700;
    wire N__15697;
    wire N__15694;
    wire N__15691;
    wire N__15688;
    wire N__15685;
    wire N__15682;
    wire N__15679;
    wire N__15676;
    wire N__15673;
    wire N__15670;
    wire N__15667;
    wire N__15664;
    wire N__15661;
    wire N__15658;
    wire N__15655;
    wire N__15652;
    wire N__15649;
    wire N__15646;
    wire N__15643;
    wire N__15640;
    wire N__15637;
    wire N__15634;
    wire N__15631;
    wire N__15628;
    wire N__15625;
    wire N__15622;
    wire N__15619;
    wire N__15616;
    wire N__15613;
    wire N__15610;
    wire N__15607;
    wire N__15602;
    wire N__15601;
    wire N__15598;
    wire N__15595;
    wire N__15592;
    wire N__15589;
    wire N__15586;
    wire N__15583;
    wire N__15580;
    wire N__15575;
    wire N__15572;
    wire N__15569;
    wire N__15566;
    wire N__15565;
    wire N__15562;
    wire N__15559;
    wire N__15556;
    wire N__15553;
    wire N__15550;
    wire N__15547;
    wire N__15544;
    wire N__15541;
    wire N__15536;
    wire N__15533;
    wire N__15532;
    wire N__15529;
    wire N__15528;
    wire N__15527;
    wire N__15524;
    wire N__15521;
    wire N__15518;
    wire N__15515;
    wire N__15510;
    wire N__15503;
    wire N__15500;
    wire N__15497;
    wire N__15496;
    wire N__15493;
    wire N__15492;
    wire N__15489;
    wire N__15488;
    wire N__15485;
    wire N__15482;
    wire N__15479;
    wire N__15476;
    wire N__15469;
    wire N__15464;
    wire N__15461;
    wire N__15460;
    wire N__15457;
    wire N__15454;
    wire N__15449;
    wire N__15446;
    wire N__15443;
    wire N__15440;
    wire N__15437;
    wire N__15434;
    wire N__15431;
    wire N__15430;
    wire N__15429;
    wire N__15426;
    wire N__15423;
    wire N__15420;
    wire N__15415;
    wire N__15410;
    wire N__15407;
    wire N__15404;
    wire N__15401;
    wire N__15398;
    wire N__15395;
    wire N__15392;
    wire N__15389;
    wire N__15386;
    wire N__15385;
    wire N__15382;
    wire N__15381;
    wire N__15378;
    wire N__15377;
    wire N__15374;
    wire N__15371;
    wire N__15368;
    wire N__15365;
    wire N__15356;
    wire N__15353;
    wire N__15352;
    wire N__15351;
    wire N__15350;
    wire N__15347;
    wire N__15342;
    wire N__15339;
    wire N__15334;
    wire N__15329;
    wire N__15326;
    wire N__15323;
    wire N__15320;
    wire N__15317;
    wire N__15314;
    wire N__15311;
    wire N__15308;
    wire N__15305;
    wire N__15304;
    wire N__15301;
    wire N__15300;
    wire N__15299;
    wire N__15296;
    wire N__15293;
    wire N__15290;
    wire N__15287;
    wire N__15284;
    wire N__15275;
    wire N__15272;
    wire N__15269;
    wire N__15268;
    wire N__15265;
    wire N__15262;
    wire N__15257;
    wire N__15256;
    wire N__15255;
    wire N__15254;
    wire N__15253;
    wire N__15252;
    wire N__15251;
    wire N__15250;
    wire N__15249;
    wire N__15248;
    wire N__15245;
    wire N__15244;
    wire N__15241;
    wire N__15240;
    wire N__15237;
    wire N__15234;
    wire N__15231;
    wire N__15228;
    wire N__15225;
    wire N__15222;
    wire N__15221;
    wire N__15220;
    wire N__15219;
    wire N__15216;
    wire N__15213;
    wire N__15212;
    wire N__15209;
    wire N__15206;
    wire N__15203;
    wire N__15200;
    wire N__15199;
    wire N__15196;
    wire N__15191;
    wire N__15188;
    wire N__15183;
    wire N__15180;
    wire N__15177;
    wire N__15174;
    wire N__15171;
    wire N__15168;
    wire N__15165;
    wire N__15164;
    wire N__15161;
    wire N__15158;
    wire N__15153;
    wire N__15150;
    wire N__15147;
    wire N__15142;
    wire N__15135;
    wire N__15132;
    wire N__15129;
    wire N__15124;
    wire N__15121;
    wire N__15112;
    wire N__15103;
    wire N__15098;
    wire N__15095;
    wire N__15092;
    wire N__15083;
    wire N__15080;
    wire N__15077;
    wire N__15074;
    wire N__15073;
    wire N__15072;
    wire N__15069;
    wire N__15066;
    wire N__15063;
    wire N__15060;
    wire N__15053;
    wire N__15052;
    wire N__15049;
    wire N__15048;
    wire N__15045;
    wire N__15042;
    wire N__15039;
    wire N__15036;
    wire N__15033;
    wire N__15026;
    wire N__15023;
    wire N__15020;
    wire N__15017;
    wire N__15016;
    wire N__15013;
    wire N__15012;
    wire N__15009;
    wire N__15006;
    wire N__15005;
    wire N__15002;
    wire N__14997;
    wire N__14994;
    wire N__14987;
    wire N__14984;
    wire N__14983;
    wire N__14982;
    wire N__14979;
    wire N__14976;
    wire N__14973;
    wire N__14970;
    wire N__14963;
    wire N__14960;
    wire N__14959;
    wire N__14956;
    wire N__14955;
    wire N__14954;
    wire N__14951;
    wire N__14948;
    wire N__14945;
    wire N__14942;
    wire N__14937;
    wire N__14930;
    wire N__14929;
    wire N__14926;
    wire N__14923;
    wire N__14922;
    wire N__14917;
    wire N__14916;
    wire N__14913;
    wire N__14910;
    wire N__14907;
    wire N__14900;
    wire N__14897;
    wire N__14896;
    wire N__14893;
    wire N__14892;
    wire N__14891;
    wire N__14888;
    wire N__14885;
    wire N__14880;
    wire N__14873;
    wire N__14872;
    wire N__14869;
    wire N__14866;
    wire N__14861;
    wire N__14858;
    wire N__14857;
    wire N__14854;
    wire N__14851;
    wire N__14848;
    wire N__14845;
    wire N__14840;
    wire N__14837;
    wire N__14834;
    wire N__14831;
    wire N__14828;
    wire N__14825;
    wire N__14822;
    wire N__14819;
    wire N__14816;
    wire N__14813;
    wire N__14812;
    wire N__14811;
    wire N__14810;
    wire N__14807;
    wire N__14804;
    wire N__14803;
    wire N__14800;
    wire N__14799;
    wire N__14796;
    wire N__14795;
    wire N__14794;
    wire N__14791;
    wire N__14788;
    wire N__14785;
    wire N__14782;
    wire N__14779;
    wire N__14778;
    wire N__14775;
    wire N__14772;
    wire N__14769;
    wire N__14764;
    wire N__14757;
    wire N__14754;
    wire N__14747;
    wire N__14738;
    wire N__14735;
    wire N__14734;
    wire N__14733;
    wire N__14732;
    wire N__14731;
    wire N__14730;
    wire N__14729;
    wire N__14726;
    wire N__14723;
    wire N__14722;
    wire N__14719;
    wire N__14718;
    wire N__14715;
    wire N__14714;
    wire N__14711;
    wire N__14708;
    wire N__14705;
    wire N__14702;
    wire N__14687;
    wire N__14684;
    wire N__14681;
    wire N__14676;
    wire N__14675;
    wire N__14670;
    wire N__14669;
    wire N__14668;
    wire N__14665;
    wire N__14662;
    wire N__14659;
    wire N__14656;
    wire N__14655;
    wire N__14654;
    wire N__14653;
    wire N__14650;
    wire N__14649;
    wire N__14644;
    wire N__14643;
    wire N__14640;
    wire N__14637;
    wire N__14634;
    wire N__14631;
    wire N__14628;
    wire N__14625;
    wire N__14622;
    wire N__14621;
    wire N__14620;
    wire N__14617;
    wire N__14614;
    wire N__14603;
    wire N__14600;
    wire N__14597;
    wire N__14594;
    wire N__14591;
    wire N__14576;
    wire N__14575;
    wire N__14574;
    wire N__14573;
    wire N__14570;
    wire N__14567;
    wire N__14566;
    wire N__14565;
    wire N__14562;
    wire N__14561;
    wire N__14560;
    wire N__14557;
    wire N__14554;
    wire N__14551;
    wire N__14548;
    wire N__14545;
    wire N__14542;
    wire N__14539;
    wire N__14536;
    wire N__14533;
    wire N__14532;
    wire N__14529;
    wire N__14526;
    wire N__14523;
    wire N__14520;
    wire N__14517;
    wire N__14514;
    wire N__14511;
    wire N__14508;
    wire N__14505;
    wire N__14500;
    wire N__14493;
    wire N__14490;
    wire N__14485;
    wire N__14474;
    wire N__14473;
    wire N__14472;
    wire N__14471;
    wire N__14468;
    wire N__14467;
    wire N__14464;
    wire N__14461;
    wire N__14460;
    wire N__14457;
    wire N__14456;
    wire N__14455;
    wire N__14452;
    wire N__14449;
    wire N__14446;
    wire N__14443;
    wire N__14440;
    wire N__14437;
    wire N__14434;
    wire N__14431;
    wire N__14430;
    wire N__14423;
    wire N__14414;
    wire N__14411;
    wire N__14408;
    wire N__14399;
    wire N__14396;
    wire N__14395;
    wire N__14394;
    wire N__14393;
    wire N__14390;
    wire N__14387;
    wire N__14384;
    wire N__14381;
    wire N__14376;
    wire N__14371;
    wire N__14366;
    wire N__14363;
    wire N__14360;
    wire N__14357;
    wire N__14354;
    wire N__14351;
    wire N__14348;
    wire N__14347;
    wire N__14346;
    wire N__14343;
    wire N__14340;
    wire N__14339;
    wire N__14336;
    wire N__14335;
    wire N__14334;
    wire N__14331;
    wire N__14328;
    wire N__14327;
    wire N__14324;
    wire N__14321;
    wire N__14318;
    wire N__14315;
    wire N__14312;
    wire N__14309;
    wire N__14306;
    wire N__14305;
    wire N__14302;
    wire N__14295;
    wire N__14290;
    wire N__14287;
    wire N__14284;
    wire N__14279;
    wire N__14272;
    wire N__14267;
    wire N__14264;
    wire N__14261;
    wire N__14258;
    wire N__14255;
    wire N__14252;
    wire N__14249;
    wire N__14248;
    wire N__14247;
    wire N__14246;
    wire N__14243;
    wire N__14240;
    wire N__14239;
    wire N__14236;
    wire N__14233;
    wire N__14228;
    wire N__14225;
    wire N__14222;
    wire N__14217;
    wire N__14214;
    wire N__14207;
    wire N__14204;
    wire N__14203;
    wire N__14200;
    wire N__14197;
    wire N__14194;
    wire N__14191;
    wire N__14186;
    wire N__14183;
    wire N__14182;
    wire N__14179;
    wire N__14176;
    wire N__14175;
    wire N__14174;
    wire N__14169;
    wire N__14166;
    wire N__14163;
    wire N__14156;
    wire N__14153;
    wire N__14150;
    wire N__14147;
    wire N__14144;
    wire N__14141;
    wire N__14138;
    wire N__14135;
    wire N__14132;
    wire N__14131;
    wire N__14128;
    wire N__14125;
    wire N__14122;
    wire N__14119;
    wire N__14116;
    wire N__14113;
    wire N__14110;
    wire N__14107;
    wire N__14104;
    wire N__14101;
    wire N__14098;
    wire N__14095;
    wire N__14092;
    wire N__14089;
    wire N__14086;
    wire N__14083;
    wire N__14080;
    wire N__14077;
    wire N__14074;
    wire N__14071;
    wire N__14068;
    wire N__14065;
    wire N__14062;
    wire N__14059;
    wire N__14056;
    wire N__14053;
    wire N__14050;
    wire N__14047;
    wire N__14044;
    wire N__14041;
    wire N__14038;
    wire N__14035;
    wire N__14032;
    wire N__14029;
    wire N__14026;
    wire N__14023;
    wire N__14020;
    wire N__14017;
    wire N__14014;
    wire N__14011;
    wire N__14008;
    wire N__14005;
    wire N__14002;
    wire N__13999;
    wire N__13996;
    wire N__13993;
    wire N__13990;
    wire N__13987;
    wire N__13984;
    wire N__13981;
    wire N__13978;
    wire N__13975;
    wire N__13972;
    wire N__13969;
    wire N__13966;
    wire N__13963;
    wire N__13960;
    wire N__13957;
    wire N__13954;
    wire N__13951;
    wire N__13948;
    wire N__13945;
    wire N__13942;
    wire N__13939;
    wire N__13936;
    wire N__13933;
    wire N__13930;
    wire N__13927;
    wire N__13922;
    wire N__13919;
    wire N__13916;
    wire N__13913;
    wire N__13910;
    wire N__13907;
    wire N__13904;
    wire N__13901;
    wire N__13898;
    wire N__13895;
    wire N__13892;
    wire N__13891;
    wire N__13890;
    wire N__13889;
    wire N__13886;
    wire N__13883;
    wire N__13880;
    wire N__13877;
    wire N__13868;
    wire N__13867;
    wire N__13864;
    wire N__13863;
    wire N__13862;
    wire N__13859;
    wire N__13856;
    wire N__13853;
    wire N__13850;
    wire N__13841;
    wire N__13840;
    wire N__13839;
    wire N__13838;
    wire N__13835;
    wire N__13832;
    wire N__13829;
    wire N__13826;
    wire N__13823;
    wire N__13814;
    wire N__13813;
    wire N__13812;
    wire N__13811;
    wire N__13808;
    wire N__13805;
    wire N__13800;
    wire N__13793;
    wire N__13790;
    wire N__13789;
    wire N__13788;
    wire N__13787;
    wire N__13784;
    wire N__13781;
    wire N__13776;
    wire N__13769;
    wire N__13768;
    wire N__13765;
    wire N__13764;
    wire N__13763;
    wire N__13758;
    wire N__13755;
    wire N__13752;
    wire N__13747;
    wire N__13742;
    wire N__13739;
    wire N__13736;
    wire N__13735;
    wire N__13734;
    wire N__13733;
    wire N__13728;
    wire N__13725;
    wire N__13722;
    wire N__13719;
    wire N__13712;
    wire N__13709;
    wire N__13708;
    wire N__13705;
    wire N__13702;
    wire N__13697;
    wire N__13694;
    wire N__13691;
    wire N__13688;
    wire N__13685;
    wire N__13682;
    wire N__13679;
    wire N__13676;
    wire N__13673;
    wire N__13670;
    wire N__13667;
    wire N__13664;
    wire N__13661;
    wire N__13658;
    wire N__13657;
    wire N__13656;
    wire N__13655;
    wire N__13652;
    wire N__13649;
    wire N__13646;
    wire N__13643;
    wire N__13634;
    wire N__13633;
    wire N__13632;
    wire N__13631;
    wire N__13628;
    wire N__13625;
    wire N__13622;
    wire N__13619;
    wire N__13610;
    wire N__13607;
    wire N__13604;
    wire N__13603;
    wire N__13602;
    wire N__13599;
    wire N__13596;
    wire N__13595;
    wire N__13592;
    wire N__13589;
    wire N__13584;
    wire N__13577;
    wire N__13574;
    wire N__13573;
    wire N__13572;
    wire N__13569;
    wire N__13568;
    wire N__13565;
    wire N__13562;
    wire N__13559;
    wire N__13556;
    wire N__13547;
    wire N__13544;
    wire N__13541;
    wire N__13540;
    wire N__13539;
    wire N__13538;
    wire N__13535;
    wire N__13532;
    wire N__13529;
    wire N__13526;
    wire N__13517;
    wire N__13514;
    wire N__13513;
    wire N__13512;
    wire N__13511;
    wire N__13508;
    wire N__13503;
    wire N__13500;
    wire N__13493;
    wire N__13490;
    wire N__13487;
    wire N__13486;
    wire N__13485;
    wire N__13484;
    wire N__13481;
    wire N__13478;
    wire N__13475;
    wire N__13472;
    wire N__13467;
    wire N__13464;
    wire N__13461;
    wire N__13456;
    wire N__13453;
    wire N__13448;
    wire N__13445;
    wire N__13442;
    wire N__13439;
    wire N__13436;
    wire N__13433;
    wire N__13430;
    wire N__13427;
    wire N__13424;
    wire N__13421;
    wire N__13418;
    wire N__13415;
    wire N__13412;
    wire N__13409;
    wire N__13406;
    wire N__13403;
    wire N__13400;
    wire N__13399;
    wire N__13396;
    wire N__13393;
    wire N__13392;
    wire N__13389;
    wire N__13386;
    wire N__13383;
    wire N__13380;
    wire N__13375;
    wire N__13374;
    wire N__13371;
    wire N__13368;
    wire N__13365;
    wire N__13358;
    wire N__13355;
    wire N__13352;
    wire N__13349;
    wire N__13346;
    wire N__13343;
    wire N__13342;
    wire N__13341;
    wire N__13340;
    wire N__13337;
    wire N__13334;
    wire N__13331;
    wire N__13328;
    wire N__13325;
    wire N__13322;
    wire N__13313;
    wire N__13312;
    wire N__13311;
    wire N__13310;
    wire N__13307;
    wire N__13304;
    wire N__13299;
    wire N__13292;
    wire N__13291;
    wire N__13290;
    wire N__13287;
    wire N__13284;
    wire N__13281;
    wire N__13274;
    wire N__13271;
    wire N__13270;
    wire N__13265;
    wire N__13262;
    wire N__13259;
    wire N__13256;
    wire N__13255;
    wire N__13250;
    wire N__13247;
    wire N__13244;
    wire N__13241;
    wire N__13238;
    wire N__13235;
    wire N__13232;
    wire N__13229;
    wire N__13226;
    wire N__13223;
    wire N__13220;
    wire N__13217;
    wire N__13214;
    wire N__13211;
    wire N__13210;
    wire N__13209;
    wire N__13206;
    wire N__13201;
    wire N__13196;
    wire N__13193;
    wire N__13192;
    wire N__13191;
    wire N__13188;
    wire N__13185;
    wire N__13182;
    wire N__13175;
    wire N__13172;
    wire N__13169;
    wire N__13166;
    wire N__13165;
    wire N__13162;
    wire N__13159;
    wire N__13156;
    wire N__13153;
    wire N__13148;
    wire N__13145;
    wire N__13142;
    wire N__13141;
    wire N__13138;
    wire N__13135;
    wire N__13130;
    wire N__13129;
    wire N__13126;
    wire N__13123;
    wire N__13122;
    wire N__13121;
    wire N__13120;
    wire N__13119;
    wire N__13118;
    wire N__13117;
    wire N__13116;
    wire N__13111;
    wire N__13096;
    wire N__13095;
    wire N__13090;
    wire N__13089;
    wire N__13088;
    wire N__13087;
    wire N__13086;
    wire N__13083;
    wire N__13080;
    wire N__13077;
    wire N__13074;
    wire N__13069;
    wire N__13068;
    wire N__13067;
    wire N__13064;
    wire N__13059;
    wire N__13054;
    wire N__13049;
    wire N__13040;
    wire N__13037;
    wire N__13036;
    wire N__13033;
    wire N__13030;
    wire N__13027;
    wire N__13024;
    wire N__13021;
    wire N__13018;
    wire N__13015;
    wire N__13012;
    wire N__13009;
    wire N__13006;
    wire N__13003;
    wire N__13000;
    wire N__12997;
    wire N__12994;
    wire N__12991;
    wire N__12988;
    wire N__12985;
    wire N__12982;
    wire N__12979;
    wire N__12976;
    wire N__12973;
    wire N__12970;
    wire N__12967;
    wire N__12964;
    wire N__12961;
    wire N__12958;
    wire N__12955;
    wire N__12952;
    wire N__12949;
    wire N__12946;
    wire N__12943;
    wire N__12940;
    wire N__12937;
    wire N__12934;
    wire N__12931;
    wire N__12928;
    wire N__12925;
    wire N__12922;
    wire N__12919;
    wire N__12916;
    wire N__12913;
    wire N__12910;
    wire N__12907;
    wire N__12904;
    wire N__12901;
    wire N__12898;
    wire N__12895;
    wire N__12892;
    wire N__12889;
    wire N__12886;
    wire N__12883;
    wire N__12880;
    wire N__12877;
    wire N__12874;
    wire N__12871;
    wire N__12868;
    wire N__12865;
    wire N__12862;
    wire N__12859;
    wire N__12856;
    wire N__12853;
    wire N__12850;
    wire N__12847;
    wire N__12844;
    wire N__12841;
    wire N__12838;
    wire N__12835;
    wire N__12832;
    wire N__12831;
    wire N__12830;
    wire N__12825;
    wire N__12822;
    wire N__12819;
    wire N__12816;
    wire N__12809;
    wire N__12808;
    wire N__12805;
    wire N__12802;
    wire N__12799;
    wire N__12796;
    wire N__12795;
    wire N__12790;
    wire N__12787;
    wire N__12786;
    wire N__12781;
    wire N__12778;
    wire N__12773;
    wire N__12772;
    wire N__12771;
    wire N__12768;
    wire N__12765;
    wire N__12762;
    wire N__12761;
    wire N__12760;
    wire N__12755;
    wire N__12752;
    wire N__12749;
    wire N__12746;
    wire N__12743;
    wire N__12736;
    wire N__12731;
    wire N__12728;
    wire N__12725;
    wire N__12722;
    wire N__12719;
    wire N__12716;
    wire N__12713;
    wire N__12710;
    wire N__12707;
    wire N__12704;
    wire N__12701;
    wire N__12698;
    wire N__12695;
    wire N__12692;
    wire N__12691;
    wire N__12690;
    wire N__12687;
    wire N__12684;
    wire N__12681;
    wire N__12680;
    wire N__12673;
    wire N__12670;
    wire N__12667;
    wire N__12664;
    wire N__12661;
    wire N__12658;
    wire N__12655;
    wire N__12652;
    wire N__12649;
    wire N__12646;
    wire N__12641;
    wire N__12638;
    wire N__12635;
    wire N__12632;
    wire N__12629;
    wire N__12626;
    wire N__12623;
    wire N__12622;
    wire N__12619;
    wire N__12616;
    wire N__12611;
    wire N__12610;
    wire N__12607;
    wire N__12604;
    wire N__12599;
    wire N__12598;
    wire N__12595;
    wire N__12592;
    wire N__12587;
    wire N__12586;
    wire N__12583;
    wire N__12580;
    wire N__12575;
    wire N__12574;
    wire N__12571;
    wire N__12568;
    wire N__12563;
    wire N__12562;
    wire N__12559;
    wire N__12556;
    wire N__12551;
    wire N__12550;
    wire N__12547;
    wire N__12544;
    wire N__12539;
    wire N__12536;
    wire N__12533;
    wire N__12530;
    wire N__12527;
    wire N__12524;
    wire N__12521;
    wire N__12520;
    wire N__12517;
    wire N__12514;
    wire N__12509;
    wire N__12506;
    wire N__12503;
    wire N__12500;
    wire N__12497;
    wire N__12494;
    wire N__12491;
    wire N__12488;
    wire N__12485;
    wire N__12482;
    wire N__12479;
    wire N__12476;
    wire N__12473;
    wire N__12472;
    wire N__12469;
    wire N__12466;
    wire N__12463;
    wire N__12460;
    wire N__12457;
    wire N__12454;
    wire N__12451;
    wire N__12448;
    wire N__12445;
    wire N__12442;
    wire N__12439;
    wire N__12436;
    wire N__12433;
    wire N__12430;
    wire N__12427;
    wire N__12424;
    wire N__12421;
    wire N__12418;
    wire N__12415;
    wire N__12412;
    wire N__12409;
    wire N__12406;
    wire N__12403;
    wire N__12400;
    wire N__12397;
    wire N__12394;
    wire N__12391;
    wire N__12388;
    wire N__12385;
    wire N__12382;
    wire N__12379;
    wire N__12376;
    wire N__12373;
    wire N__12370;
    wire N__12367;
    wire N__12364;
    wire N__12361;
    wire N__12358;
    wire N__12355;
    wire N__12352;
    wire N__12349;
    wire N__12346;
    wire N__12343;
    wire N__12340;
    wire N__12337;
    wire N__12334;
    wire N__12331;
    wire N__12328;
    wire N__12325;
    wire N__12322;
    wire N__12319;
    wire N__12316;
    wire N__12313;
    wire N__12310;
    wire N__12307;
    wire N__12304;
    wire N__12301;
    wire N__12298;
    wire N__12295;
    wire N__12294;
    wire N__12291;
    wire N__12288;
    wire N__12285;
    wire N__12282;
    wire N__12279;
    wire N__12276;
    wire N__12273;
    wire N__12270;
    wire N__12269;
    wire N__12266;
    wire N__12263;
    wire N__12260;
    wire N__12257;
    wire N__12254;
    wire N__12251;
    wire N__12248;
    wire N__12239;
    wire N__12236;
    wire N__12233;
    wire N__12230;
    wire N__12227;
    wire N__12224;
    wire N__12221;
    wire N__12220;
    wire N__12217;
    wire N__12214;
    wire N__12211;
    wire N__12208;
    wire N__12205;
    wire N__12202;
    wire N__12199;
    wire N__12196;
    wire N__12193;
    wire N__12190;
    wire N__12187;
    wire N__12184;
    wire N__12181;
    wire N__12178;
    wire N__12175;
    wire N__12172;
    wire N__12169;
    wire N__12166;
    wire N__12163;
    wire N__12160;
    wire N__12157;
    wire N__12154;
    wire N__12151;
    wire N__12148;
    wire N__12145;
    wire N__12142;
    wire N__12139;
    wire N__12136;
    wire N__12133;
    wire N__12130;
    wire N__12127;
    wire N__12124;
    wire N__12121;
    wire N__12118;
    wire N__12115;
    wire N__12112;
    wire N__12109;
    wire N__12106;
    wire N__12103;
    wire N__12100;
    wire N__12097;
    wire N__12094;
    wire N__12091;
    wire N__12088;
    wire N__12085;
    wire N__12082;
    wire N__12079;
    wire N__12076;
    wire N__12073;
    wire N__12070;
    wire N__12067;
    wire N__12064;
    wire N__12061;
    wire N__12058;
    wire N__12055;
    wire N__12052;
    wire N__12049;
    wire N__12046;
    wire N__12045;
    wire N__12042;
    wire N__12039;
    wire N__12036;
    wire N__12033;
    wire N__12030;
    wire N__12027;
    wire N__12024;
    wire N__12021;
    wire N__12018;
    wire N__12017;
    wire N__12014;
    wire N__12011;
    wire N__12008;
    wire N__12005;
    wire N__12002;
    wire N__11999;
    wire N__11990;
    wire N__11987;
    wire N__11984;
    wire N__11981;
    wire N__11978;
    wire N__11975;
    wire N__11972;
    wire N__11969;
    wire N__11966;
    wire N__11963;
    wire N__11962;
    wire N__11959;
    wire N__11956;
    wire N__11953;
    wire N__11950;
    wire N__11947;
    wire N__11944;
    wire N__11941;
    wire N__11938;
    wire N__11935;
    wire N__11932;
    wire N__11929;
    wire N__11926;
    wire N__11923;
    wire N__11920;
    wire N__11917;
    wire N__11914;
    wire N__11911;
    wire N__11908;
    wire N__11905;
    wire N__11902;
    wire N__11899;
    wire N__11896;
    wire N__11893;
    wire N__11890;
    wire N__11887;
    wire N__11884;
    wire N__11881;
    wire N__11878;
    wire N__11875;
    wire N__11872;
    wire N__11869;
    wire N__11866;
    wire N__11863;
    wire N__11860;
    wire N__11857;
    wire N__11854;
    wire N__11851;
    wire N__11848;
    wire N__11845;
    wire N__11842;
    wire N__11839;
    wire N__11836;
    wire N__11833;
    wire N__11830;
    wire N__11827;
    wire N__11824;
    wire N__11821;
    wire N__11818;
    wire N__11815;
    wire N__11812;
    wire N__11809;
    wire N__11806;
    wire N__11803;
    wire N__11800;
    wire N__11797;
    wire N__11794;
    wire N__11791;
    wire N__11788;
    wire N__11787;
    wire N__11784;
    wire N__11781;
    wire N__11778;
    wire N__11775;
    wire N__11772;
    wire N__11769;
    wire N__11766;
    wire N__11763;
    wire N__11760;
    wire N__11759;
    wire N__11756;
    wire N__11753;
    wire N__11750;
    wire N__11747;
    wire N__11744;
    wire N__11741;
    wire N__11732;
    wire N__11729;
    wire N__11726;
    wire N__11723;
    wire N__11722;
    wire N__11721;
    wire N__11718;
    wire N__11717;
    wire N__11716;
    wire N__11713;
    wire N__11712;
    wire N__11709;
    wire N__11706;
    wire N__11703;
    wire N__11700;
    wire N__11699;
    wire N__11698;
    wire N__11695;
    wire N__11692;
    wire N__11689;
    wire N__11682;
    wire N__11679;
    wire N__11676;
    wire N__11673;
    wire N__11670;
    wire N__11667;
    wire N__11660;
    wire N__11655;
    wire N__11652;
    wire N__11649;
    wire N__11646;
    wire N__11639;
    wire N__11636;
    wire N__11633;
    wire N__11630;
    wire N__11627;
    wire N__11624;
    wire N__11621;
    wire N__11618;
    wire N__11615;
    wire N__11612;
    wire N__11609;
    wire N__11606;
    wire N__11603;
    wire N__11600;
    wire N__11597;
    wire N__11596;
    wire N__11593;
    wire N__11590;
    wire N__11587;
    wire N__11584;
    wire N__11581;
    wire N__11578;
    wire N__11575;
    wire N__11572;
    wire N__11569;
    wire N__11566;
    wire N__11563;
    wire N__11560;
    wire N__11557;
    wire N__11554;
    wire N__11551;
    wire N__11548;
    wire N__11545;
    wire N__11542;
    wire N__11539;
    wire N__11536;
    wire N__11533;
    wire N__11530;
    wire N__11527;
    wire N__11524;
    wire N__11521;
    wire N__11518;
    wire N__11515;
    wire N__11512;
    wire N__11509;
    wire N__11506;
    wire N__11503;
    wire N__11500;
    wire N__11497;
    wire N__11494;
    wire N__11491;
    wire N__11488;
    wire N__11485;
    wire N__11482;
    wire N__11479;
    wire N__11476;
    wire N__11473;
    wire N__11470;
    wire N__11467;
    wire N__11464;
    wire N__11461;
    wire N__11458;
    wire N__11455;
    wire N__11452;
    wire N__11449;
    wire N__11446;
    wire N__11443;
    wire N__11440;
    wire N__11437;
    wire N__11434;
    wire N__11431;
    wire N__11428;
    wire N__11425;
    wire N__11422;
    wire N__11419;
    wire N__11416;
    wire N__11413;
    wire N__11410;
    wire N__11407;
    wire N__11404;
    wire N__11403;
    wire N__11400;
    wire N__11397;
    wire N__11394;
    wire N__11391;
    wire N__11388;
    wire N__11385;
    wire N__11382;
    wire N__11379;
    wire N__11378;
    wire N__11375;
    wire N__11372;
    wire N__11369;
    wire N__11366;
    wire N__11363;
    wire N__11358;
    wire N__11351;
    wire N__11348;
    wire N__11345;
    wire N__11342;
    wire N__11339;
    wire N__11336;
    wire N__11335;
    wire N__11332;
    wire N__11329;
    wire N__11326;
    wire N__11323;
    wire N__11320;
    wire N__11317;
    wire N__11314;
    wire N__11311;
    wire N__11308;
    wire N__11305;
    wire N__11302;
    wire N__11299;
    wire N__11296;
    wire N__11293;
    wire N__11290;
    wire N__11287;
    wire N__11284;
    wire N__11281;
    wire N__11278;
    wire N__11275;
    wire N__11272;
    wire N__11269;
    wire N__11266;
    wire N__11263;
    wire N__11260;
    wire N__11257;
    wire N__11254;
    wire N__11251;
    wire N__11248;
    wire N__11245;
    wire N__11242;
    wire N__11239;
    wire N__11236;
    wire N__11233;
    wire N__11230;
    wire N__11227;
    wire N__11224;
    wire N__11221;
    wire N__11218;
    wire N__11215;
    wire N__11212;
    wire N__11209;
    wire N__11206;
    wire N__11203;
    wire N__11200;
    wire N__11197;
    wire N__11194;
    wire N__11191;
    wire N__11188;
    wire N__11185;
    wire N__11182;
    wire N__11179;
    wire N__11176;
    wire N__11173;
    wire N__11170;
    wire N__11167;
    wire N__11164;
    wire N__11161;
    wire N__11158;
    wire N__11155;
    wire N__11152;
    wire N__11149;
    wire N__11146;
    wire N__11145;
    wire N__11142;
    wire N__11139;
    wire N__11136;
    wire N__11133;
    wire N__11130;
    wire N__11129;
    wire N__11126;
    wire N__11123;
    wire N__11120;
    wire N__11117;
    wire N__11114;
    wire N__11111;
    wire N__11108;
    wire N__11105;
    wire N__11102;
    wire N__11097;
    wire N__11090;
    wire N__11087;
    wire N__11084;
    wire N__11081;
    wire N__11078;
    wire N__11077;
    wire N__11074;
    wire N__11071;
    wire N__11068;
    wire N__11065;
    wire N__11062;
    wire N__11059;
    wire N__11056;
    wire N__11053;
    wire N__11050;
    wire N__11047;
    wire N__11044;
    wire N__11041;
    wire N__11038;
    wire N__11035;
    wire N__11032;
    wire N__11029;
    wire N__11026;
    wire N__11023;
    wire N__11020;
    wire N__11017;
    wire N__11014;
    wire N__11011;
    wire N__11008;
    wire N__11005;
    wire N__11002;
    wire N__10999;
    wire N__10996;
    wire N__10993;
    wire N__10990;
    wire N__10987;
    wire N__10984;
    wire N__10981;
    wire N__10978;
    wire N__10975;
    wire N__10972;
    wire N__10969;
    wire N__10966;
    wire N__10963;
    wire N__10960;
    wire N__10957;
    wire N__10954;
    wire N__10951;
    wire N__10948;
    wire N__10945;
    wire N__10942;
    wire N__10939;
    wire N__10936;
    wire N__10933;
    wire N__10930;
    wire N__10927;
    wire N__10924;
    wire N__10921;
    wire N__10918;
    wire N__10915;
    wire N__10912;
    wire N__10909;
    wire N__10906;
    wire N__10903;
    wire N__10900;
    wire N__10897;
    wire N__10894;
    wire N__10891;
    wire N__10888;
    wire N__10885;
    wire N__10882;
    wire N__10879;
    wire N__10876;
    wire N__10873;
    wire N__10872;
    wire N__10869;
    wire N__10866;
    wire N__10863;
    wire N__10862;
    wire N__10859;
    wire N__10856;
    wire N__10853;
    wire N__10850;
    wire N__10847;
    wire N__10844;
    wire N__10835;
    wire N__10832;
    wire N__10829;
    wire N__10826;
    wire N__10825;
    wire N__10822;
    wire N__10819;
    wire N__10816;
    wire N__10813;
    wire N__10810;
    wire N__10807;
    wire N__10804;
    wire N__10801;
    wire N__10798;
    wire N__10795;
    wire N__10792;
    wire N__10789;
    wire N__10786;
    wire N__10783;
    wire N__10780;
    wire N__10777;
    wire N__10774;
    wire N__10771;
    wire N__10768;
    wire N__10765;
    wire N__10762;
    wire N__10759;
    wire N__10756;
    wire N__10753;
    wire N__10750;
    wire N__10747;
    wire N__10744;
    wire N__10741;
    wire N__10738;
    wire N__10735;
    wire N__10732;
    wire N__10729;
    wire N__10726;
    wire N__10723;
    wire N__10720;
    wire N__10717;
    wire N__10714;
    wire N__10711;
    wire N__10708;
    wire N__10705;
    wire N__10702;
    wire N__10699;
    wire N__10696;
    wire N__10693;
    wire N__10690;
    wire N__10687;
    wire N__10684;
    wire N__10681;
    wire N__10678;
    wire N__10675;
    wire N__10672;
    wire N__10669;
    wire N__10666;
    wire N__10663;
    wire N__10660;
    wire N__10657;
    wire N__10654;
    wire N__10651;
    wire N__10648;
    wire N__10645;
    wire N__10642;
    wire N__10639;
    wire N__10636;
    wire N__10633;
    wire N__10632;
    wire N__10629;
    wire N__10626;
    wire N__10625;
    wire N__10622;
    wire N__10619;
    wire N__10616;
    wire N__10613;
    wire N__10610;
    wire N__10607;
    wire N__10604;
    wire N__10601;
    wire N__10598;
    wire N__10593;
    wire N__10586;
    wire N__10583;
    wire N__10580;
    wire N__10577;
    wire N__10574;
    wire N__10573;
    wire N__10570;
    wire N__10567;
    wire N__10564;
    wire N__10561;
    wire N__10558;
    wire N__10555;
    wire N__10552;
    wire N__10549;
    wire N__10546;
    wire N__10543;
    wire N__10540;
    wire N__10537;
    wire N__10534;
    wire N__10531;
    wire N__10528;
    wire N__10525;
    wire N__10522;
    wire N__10519;
    wire N__10516;
    wire N__10513;
    wire N__10510;
    wire N__10507;
    wire N__10504;
    wire N__10501;
    wire N__10498;
    wire N__10495;
    wire N__10492;
    wire N__10489;
    wire N__10486;
    wire N__10483;
    wire N__10480;
    wire N__10477;
    wire N__10474;
    wire N__10471;
    wire N__10468;
    wire N__10465;
    wire N__10462;
    wire N__10459;
    wire N__10456;
    wire N__10453;
    wire N__10450;
    wire N__10447;
    wire N__10444;
    wire N__10441;
    wire N__10438;
    wire N__10435;
    wire N__10432;
    wire N__10429;
    wire N__10426;
    wire N__10423;
    wire N__10420;
    wire N__10417;
    wire N__10414;
    wire N__10411;
    wire N__10408;
    wire N__10405;
    wire N__10402;
    wire N__10399;
    wire N__10396;
    wire N__10393;
    wire N__10390;
    wire N__10387;
    wire N__10384;
    wire N__10381;
    wire N__10378;
    wire N__10375;
    wire N__10372;
    wire N__10371;
    wire N__10368;
    wire N__10365;
    wire N__10362;
    wire N__10357;
    wire N__10356;
    wire N__10353;
    wire N__10350;
    wire N__10347;
    wire N__10344;
    wire N__10341;
    wire N__10334;
    wire N__10331;
    wire N__10328;
    wire N__10325;
    wire N__10324;
    wire N__10321;
    wire N__10318;
    wire N__10315;
    wire N__10312;
    wire N__10309;
    wire N__10306;
    wire N__10303;
    wire N__10300;
    wire N__10297;
    wire N__10294;
    wire N__10291;
    wire N__10288;
    wire N__10285;
    wire N__10282;
    wire N__10279;
    wire N__10276;
    wire N__10273;
    wire N__10270;
    wire N__10267;
    wire N__10264;
    wire N__10261;
    wire N__10258;
    wire N__10255;
    wire N__10252;
    wire N__10249;
    wire N__10246;
    wire N__10243;
    wire N__10240;
    wire N__10237;
    wire N__10234;
    wire N__10231;
    wire N__10228;
    wire N__10225;
    wire N__10222;
    wire N__10219;
    wire N__10216;
    wire N__10213;
    wire N__10210;
    wire N__10207;
    wire N__10204;
    wire N__10201;
    wire N__10198;
    wire N__10195;
    wire N__10192;
    wire N__10189;
    wire N__10186;
    wire N__10183;
    wire N__10180;
    wire N__10177;
    wire N__10174;
    wire N__10171;
    wire N__10168;
    wire N__10165;
    wire N__10162;
    wire N__10159;
    wire N__10156;
    wire N__10153;
    wire N__10150;
    wire N__10147;
    wire N__10144;
    wire N__10141;
    wire N__10138;
    wire N__10135;
    wire N__10132;
    wire N__10129;
    wire N__10128;
    wire N__10125;
    wire N__10122;
    wire N__10119;
    wire N__10116;
    wire N__10113;
    wire N__10110;
    wire N__10107;
    wire N__10106;
    wire N__10103;
    wire N__10100;
    wire N__10097;
    wire N__10094;
    wire N__10091;
    wire N__10086;
    wire N__10079;
    wire N__10076;
    wire N__10073;
    wire N__10070;
    wire N__10067;
    wire N__10066;
    wire N__10063;
    wire N__10060;
    wire N__10057;
    wire N__10054;
    wire N__10051;
    wire N__10048;
    wire N__10045;
    wire N__10042;
    wire N__10039;
    wire N__10036;
    wire N__10033;
    wire N__10030;
    wire N__10027;
    wire N__10024;
    wire N__10021;
    wire N__10018;
    wire N__10015;
    wire N__10012;
    wire N__10009;
    wire N__10006;
    wire N__10003;
    wire N__10000;
    wire N__9997;
    wire N__9994;
    wire N__9991;
    wire N__9988;
    wire N__9985;
    wire N__9982;
    wire N__9979;
    wire N__9976;
    wire N__9973;
    wire N__9970;
    wire N__9967;
    wire N__9964;
    wire N__9961;
    wire N__9958;
    wire N__9955;
    wire N__9952;
    wire N__9949;
    wire N__9946;
    wire N__9943;
    wire N__9940;
    wire N__9937;
    wire N__9934;
    wire N__9931;
    wire N__9928;
    wire N__9925;
    wire N__9922;
    wire N__9919;
    wire N__9916;
    wire N__9913;
    wire N__9910;
    wire N__9907;
    wire N__9904;
    wire N__9901;
    wire N__9898;
    wire N__9895;
    wire N__9892;
    wire N__9889;
    wire N__9886;
    wire N__9883;
    wire N__9880;
    wire N__9877;
    wire N__9874;
    wire N__9871;
    wire N__9870;
    wire N__9867;
    wire N__9864;
    wire N__9861;
    wire N__9858;
    wire N__9855;
    wire N__9852;
    wire N__9851;
    wire N__9848;
    wire N__9845;
    wire N__9842;
    wire N__9839;
    wire N__9836;
    wire N__9833;
    wire N__9824;
    wire N__9821;
    wire N__9818;
    wire N__9815;
    wire N__9812;
    wire N__9809;
    wire N__9806;
    wire N__9803;
    wire N__9800;
    wire N__9797;
    wire N__9794;
    wire N__9791;
    wire N__9788;
    wire N__9785;
    wire N__9782;
    wire N__9779;
    wire N__9776;
    wire N__9773;
    wire N__9770;
    wire N__9767;
    wire N__9764;
    wire N__9761;
    wire N__9758;
    wire N__9755;
    wire N__9752;
    wire N__9749;
    wire N__9746;
    wire N__9743;
    wire N__9740;
    wire N__9737;
    wire N__9734;
    wire N__9731;
    wire N__9728;
    wire N__9725;
    wire N__9722;
    wire N__9719;
    wire N__9716;
    wire N__9713;
    wire N__9710;
    wire N__9707;
    wire N__9704;
    wire N__9701;
    wire N__9698;
    wire N__9695;
    wire N__9692;
    wire N__9689;
    wire N__9686;
    wire N__9683;
    wire N__9680;
    wire N__9677;
    wire N__9674;
    wire N__9671;
    wire N__9668;
    wire N__9665;
    wire N__9662;
    wire N__9659;
    wire N__9656;
    wire N__9653;
    wire N__9650;
    wire N__9647;
    wire N__9644;
    wire N__9641;
    wire N__9640;
    wire N__9637;
    wire N__9636;
    wire N__9633;
    wire N__9630;
    wire N__9627;
    wire N__9624;
    wire N__9619;
    wire N__9618;
    wire N__9613;
    wire N__9610;
    wire N__9605;
    wire N__9602;
    wire N__9601;
    wire N__9600;
    wire N__9597;
    wire N__9592;
    wire N__9587;
    wire N__9586;
    wire N__9585;
    wire N__9582;
    wire N__9577;
    wire N__9572;
    wire N__9571;
    wire N__9570;
    wire N__9567;
    wire N__9562;
    wire N__9557;
    wire N__9556;
    wire N__9555;
    wire N__9552;
    wire N__9547;
    wire N__9542;
    wire N__9539;
    wire N__9538;
    wire N__9537;
    wire N__9534;
    wire N__9529;
    wire N__9524;
    wire N__9521;
    wire N__9518;
    wire N__9515;
    wire N__9512;
    wire N__9509;
    wire N__9508;
    wire N__9505;
    wire N__9504;
    wire N__9501;
    wire N__9498;
    wire N__9495;
    wire N__9488;
    wire N__9485;
    wire N__9482;
    wire N__9479;
    wire N__9476;
    wire N__9473;
    wire N__9470;
    wire N__9469;
    wire N__9466;
    wire N__9463;
    wire N__9458;
    wire N__9455;
    wire N__9452;
    wire N__9449;
    wire N__9446;
    wire N__9443;
    wire N__9442;
    wire N__9439;
    wire N__9436;
    wire N__9431;
    wire N__9430;
    wire N__9427;
    wire N__9424;
    wire N__9421;
    wire N__9416;
    wire N__9415;
    wire N__9412;
    wire N__9409;
    wire N__9406;
    wire N__9403;
    wire N__9400;
    wire N__9397;
    wire N__9392;
    wire N__9389;
    wire N__9386;
    wire N__9383;
    wire N__9382;
    wire N__9379;
    wire N__9376;
    wire N__9375;
    wire N__9370;
    wire N__9367;
    wire N__9362;
    wire N__9361;
    wire N__9358;
    wire N__9355;
    wire N__9352;
    wire N__9349;
    wire N__9346;
    wire N__9343;
    wire N__9340;
    wire N__9337;
    wire N__9334;
    wire N__9331;
    wire N__9326;
    wire N__9323;
    wire N__9320;
    wire N__9317;
    wire N__9314;
    wire N__9311;
    wire N__9308;
    wire N__9305;
    wire N__9302;
    wire N__9299;
    wire N__9296;
    wire N__9293;
    wire N__9290;
    wire N__9287;
    wire N__9284;
    wire N__9281;
    wire N__9278;
    wire N__9275;
    wire N__9272;
    wire N__9269;
    wire N__9266;
    wire N__9263;
    wire N__9260;
    wire N__9257;
    wire N__9256;
    wire N__9253;
    wire N__9250;
    wire N__9247;
    wire N__9244;
    wire N__9241;
    wire N__9238;
    wire N__9235;
    wire N__9232;
    wire N__9229;
    wire N__9226;
    wire N__9223;
    wire N__9220;
    wire N__9217;
    wire N__9214;
    wire N__9211;
    wire N__9208;
    wire N__9205;
    wire N__9202;
    wire N__9199;
    wire N__9196;
    wire N__9193;
    wire N__9190;
    wire N__9187;
    wire N__9184;
    wire N__9181;
    wire N__9178;
    wire N__9175;
    wire N__9172;
    wire N__9169;
    wire N__9166;
    wire N__9163;
    wire N__9160;
    wire N__9157;
    wire N__9154;
    wire N__9151;
    wire N__9148;
    wire N__9145;
    wire N__9142;
    wire N__9139;
    wire N__9136;
    wire N__9133;
    wire N__9130;
    wire N__9127;
    wire N__9124;
    wire N__9121;
    wire N__9118;
    wire N__9115;
    wire N__9112;
    wire N__9109;
    wire N__9106;
    wire N__9103;
    wire N__9100;
    wire N__9097;
    wire N__9094;
    wire N__9091;
    wire N__9088;
    wire N__9085;
    wire N__9082;
    wire N__9079;
    wire N__9076;
    wire N__9073;
    wire N__9070;
    wire N__9067;
    wire N__9064;
    wire N__9061;
    wire N__9058;
    wire N__9053;
    wire N__9050;
    wire N__9047;
    wire N__9044;
    wire N__9041;
    wire N__9038;
    wire N__9035;
    wire N__9032;
    wire N__9029;
    wire N__9026;
    wire N__9023;
    wire N__9020;
    wire N__9017;
    wire N__9014;
    wire N__9011;
    wire N__9008;
    wire N__9005;
    wire N__9002;
    wire N__8999;
    wire N__8996;
    wire N__8993;
    wire N__8990;
    wire N__8987;
    wire N__8984;
    wire N__8981;
    wire N__8978;
    wire N__8975;
    wire N__8972;
    wire N__8969;
    wire N__8966;
    wire N__8963;
    wire N__8960;
    wire N__8957;
    wire N__8954;
    wire N__8951;
    wire N__8948;
    wire N__8945;
    wire N__8942;
    wire N__8939;
    wire N__8936;
    wire N__8933;
    wire N__8930;
    wire N__8927;
    wire N__8924;
    wire N__8921;
    wire N__8918;
    wire N__8915;
    wire N__8912;
    wire N__8909;
    wire N__8906;
    wire N__8903;
    wire N__8900;
    wire N__8897;
    wire N__8894;
    wire N__8891;
    wire N__8888;
    wire N__8885;
    wire N__8882;
    wire N__8879;
    wire N__8876;
    wire N__8873;
    wire N__8870;
    wire N__8867;
    wire N__8864;
    wire N__8861;
    wire N__8858;
    wire N__8855;
    wire N__8852;
    wire N__8849;
    wire N__8846;
    wire N__8843;
    wire N__8840;
    wire N__8837;
    wire N__8834;
    wire N__8831;
    wire N__8828;
    wire N__8825;
    wire N__8822;
    wire N__8819;
    wire N__8816;
    wire N__8813;
    wire N__8810;
    wire N__8809;
    wire N__8806;
    wire N__8803;
    wire N__8798;
    wire N__8795;
    wire N__8792;
    wire N__8789;
    wire N__8788;
    wire N__8785;
    wire N__8782;
    wire N__8779;
    wire N__8776;
    wire N__8771;
    wire N__8768;
    wire N__8765;
    wire N__8762;
    wire N__8759;
    wire N__8756;
    wire N__8753;
    wire N__8750;
    wire N__8747;
    wire N__8744;
    wire N__8741;
    wire N__8738;
    wire N__8735;
    wire N__8732;
    wire N__8729;
    wire N__8726;
    wire N__8723;
    wire N__8720;
    wire N__8717;
    wire N__8714;
    wire N__8711;
    wire N__8708;
    wire N__8705;
    wire N__8702;
    wire N__8699;
    wire N__8696;
    wire N__8693;
    wire N__8690;
    wire N__8687;
    wire N__8684;
    wire N__8681;
    wire N__8678;
    wire N__8675;
    wire N__8672;
    wire N__8669;
    wire N__8666;
    wire N__8663;
    wire N__8660;
    wire N__8657;
    wire N__8654;
    wire N__8651;
    wire N__8648;
    wire N__8645;
    wire N__8642;
    wire N__8639;
    wire N__8636;
    wire N__8633;
    wire N__8630;
    wire N__8627;
    wire N__8624;
    wire N__8621;
    wire N__8618;
    wire N__8615;
    wire N__8614;
    wire N__8613;
    wire N__8610;
    wire N__8607;
    wire N__8604;
    wire N__8603;
    wire N__8600;
    wire N__8595;
    wire N__8592;
    wire N__8589;
    wire N__8584;
    wire N__8581;
    wire N__8578;
    wire N__8575;
    wire N__8572;
    wire N__8567;
    wire N__8564;
    wire N__8561;
    wire N__8558;
    wire N__8555;
    wire N__8552;
    wire N__8549;
    wire N__8546;
    wire N__8543;
    wire N__8540;
    wire N__8537;
    wire N__8534;
    wire N__8531;
    wire N__8528;
    wire N__8525;
    wire N__8522;
    wire N__8519;
    wire N__8516;
    wire N__8513;
    wire N__8510;
    wire N__8507;
    wire N__8504;
    wire N__8501;
    wire N__8498;
    wire N__8495;
    wire N__8492;
    wire N__8489;
    wire N__8486;
    wire N__8483;
    wire N__8480;
    wire N__8477;
    wire N__8474;
    wire N__8471;
    wire N__8468;
    wire N__8465;
    wire N__8462;
    wire N__8459;
    wire N__8456;
    wire N__8453;
    wire N__8450;
    wire N__8447;
    wire N__8444;
    wire N__8441;
    wire N__8438;
    wire N__8435;
    wire N__8432;
    wire N__8429;
    wire N__8426;
    wire N__8423;
    wire N__8420;
    wire N__8417;
    wire N__8414;
    wire N__8411;
    wire N__8408;
    wire N__8405;
    wire N__8402;
    wire N__8399;
    wire N__8396;
    wire N__8395;
    wire N__8392;
    wire N__8389;
    wire N__8386;
    wire N__8383;
    wire N__8380;
    wire N__8377;
    wire N__8374;
    wire N__8371;
    wire N__8366;
    wire N__8363;
    wire N__8360;
    wire N__8357;
    wire N__8354;
    wire N__8351;
    wire N__8348;
    wire N__8345;
    wire N__8342;
    wire N__8339;
    wire VCCG0;
    wire GNDG0;
    wire GB_BUFFER_DEBUG_c_2_c_THRU_CO;
    wire \transmit_module.Y_DELTA_PATTERN_70 ;
    wire TVP_VIDEO_c_3;
    wire \transmit_module.Y_DELTA_PATTERN_71 ;
    wire \transmit_module.Y_DELTA_PATTERN_35 ;
    wire \transmit_module.Y_DELTA_PATTERN_34 ;
    wire \transmit_module.Y_DELTA_PATTERN_72 ;
    wire \transmit_module.Y_DELTA_PATTERN_90 ;
    wire \transmit_module.Y_DELTA_PATTERN_89 ;
    wire \transmit_module.Y_DELTA_PATTERN_88 ;
    wire \transmit_module.Y_DELTA_PATTERN_36 ;
    wire \transmit_module.Y_DELTA_PATTERN_81 ;
    wire \transmit_module.Y_DELTA_PATTERN_80 ;
    wire \transmit_module.Y_DELTA_PATTERN_37 ;
    wire \transmit_module.Y_DELTA_PATTERN_79 ;
    wire \transmit_module.Y_DELTA_PATTERN_66 ;
    wire \transmit_module.Y_DELTA_PATTERN_69 ;
    wire \transmit_module.Y_DELTA_PATTERN_68 ;
    wire \transmit_module.Y_DELTA_PATTERN_67 ;
    wire \transmit_module.Y_DELTA_PATTERN_48 ;
    wire TVP_VIDEO_c_2;
    wire \line_buffer.n533 ;
    wire \tvp_video_buffer.BUFFER_0_3 ;
    wire \transmit_module.Y_DELTA_PATTERN_82 ;
    wire \transmit_module.Y_DELTA_PATTERN_49 ;
    wire \transmit_module.Y_DELTA_PATTERN_84 ;
    wire \transmit_module.Y_DELTA_PATTERN_83 ;
    wire \transmit_module.Y_DELTA_PATTERN_85 ;
    wire \transmit_module.Y_DELTA_PATTERN_87 ;
    wire \transmit_module.Y_DELTA_PATTERN_86 ;
    wire \transmit_module.Y_DELTA_PATTERN_91 ;
    wire \transmit_module.Y_DELTA_PATTERN_93 ;
    wire \transmit_module.Y_DELTA_PATTERN_92 ;
    wire \transmit_module.Y_DELTA_PATTERN_94 ;
    wire \transmit_module.Y_DELTA_PATTERN_97 ;
    wire \transmit_module.Y_DELTA_PATTERN_98 ;
    wire \transmit_module.Y_DELTA_PATTERN_96 ;
    wire \transmit_module.Y_DELTA_PATTERN_95 ;
    wire \transmit_module.Y_DELTA_PATTERN_33 ;
    wire \transmit_module.Y_DELTA_PATTERN_29 ;
    wire \transmit_module.Y_DELTA_PATTERN_32 ;
    wire \transmit_module.Y_DELTA_PATTERN_31 ;
    wire \transmit_module.Y_DELTA_PATTERN_30 ;
    wire \transmit_module.Y_DELTA_PATTERN_74 ;
    wire \transmit_module.Y_DELTA_PATTERN_73 ;
    wire \transmit_module.Y_DELTA_PATTERN_65 ;
    wire \transmit_module.Y_DELTA_PATTERN_64 ;
    wire \transmit_module.Y_DELTA_PATTERN_63 ;
    wire \transmit_module.Y_DELTA_PATTERN_75 ;
    wire \transmit_module.Y_DELTA_PATTERN_62 ;
    wire \transmit_module.Y_DELTA_PATTERN_78 ;
    wire \tvp_video_buffer.BUFFER_0_2 ;
    wire LED_c;
    wire DEBUG_c_1_c;
    wire \tvp_hs_buffer.BUFFER_0_0 ;
    wire \tvp_hs_buffer.BUFFER_1_0 ;
    wire \receive_module.rx_counter.n10 ;
    wire bfn_11_9_0_;
    wire \receive_module.rx_counter.n9_adj_612 ;
    wire \receive_module.rx_counter.n3147 ;
    wire \receive_module.rx_counter.n8_adj_611 ;
    wire \receive_module.rx_counter.n3148 ;
    wire \receive_module.rx_counter.n3149 ;
    wire \receive_module.rx_counter.n3150 ;
    wire \receive_module.rx_counter.n3151 ;
    wire \receive_module.rx_counter.n3152 ;
    wire \receive_module.rx_counter.n3153 ;
    wire \receive_module.rx_counter.n3154 ;
    wire bfn_11_10_0_;
    wire \receive_module.rx_counter.n3155 ;
    wire \transmit_module.Y_DELTA_PATTERN_50 ;
    wire \transmit_module.Y_DELTA_PATTERN_51 ;
    wire \transmit_module.Y_DELTA_PATTERN_58 ;
    wire \transmit_module.Y_DELTA_PATTERN_57 ;
    wire \transmit_module.Y_DELTA_PATTERN_22 ;
    wire \transmit_module.Y_DELTA_PATTERN_21 ;
    wire \transmit_module.Y_DELTA_PATTERN_24 ;
    wire \transmit_module.Y_DELTA_PATTERN_23 ;
    wire \transmit_module.Y_DELTA_PATTERN_28 ;
    wire \transmit_module.Y_DELTA_PATTERN_27 ;
    wire \transmit_module.Y_DELTA_PATTERN_13 ;
    wire \transmit_module.Y_DELTA_PATTERN_15 ;
    wire \transmit_module.Y_DELTA_PATTERN_14 ;
    wire \transmit_module.Y_DELTA_PATTERN_26 ;
    wire \transmit_module.Y_DELTA_PATTERN_25 ;
    wire \transmit_module.Y_DELTA_PATTERN_8 ;
    wire \transmit_module.Y_DELTA_PATTERN_99 ;
    wire \transmit_module.Y_DELTA_PATTERN_10 ;
    wire \transmit_module.Y_DELTA_PATTERN_9 ;
    wire \transmit_module.Y_DELTA_PATTERN_12 ;
    wire \transmit_module.Y_DELTA_PATTERN_11 ;
    wire \transmit_module.Y_DELTA_PATTERN_38 ;
    wire \transmit_module.Y_DELTA_PATTERN_40 ;
    wire \transmit_module.Y_DELTA_PATTERN_39 ;
    wire \transmit_module.Y_DELTA_PATTERN_41 ;
    wire \transmit_module.Y_DELTA_PATTERN_42 ;
    wire \transmit_module.Y_DELTA_PATTERN_43 ;
    wire \transmit_module.Y_DELTA_PATTERN_59 ;
    wire \transmit_module.Y_DELTA_PATTERN_45 ;
    wire \transmit_module.Y_DELTA_PATTERN_44 ;
    wire \transmit_module.Y_DELTA_PATTERN_47 ;
    wire \transmit_module.Y_DELTA_PATTERN_46 ;
    wire \transmit_module.Y_DELTA_PATTERN_61 ;
    wire \transmit_module.Y_DELTA_PATTERN_60 ;
    wire \transmit_module.Y_DELTA_PATTERN_77 ;
    wire \transmit_module.Y_DELTA_PATTERN_76 ;
    wire n24;
    wire TVP_VIDEO_c_4;
    wire DEBUG_c_0_c;
    wire \INVTVP_VSYNC_buff_I_0.BUFFER_0__i1C_net ;
    wire \TVP_VSYNC_buff_I_0.BUFFER_0_0 ;
    wire \INVTVP_VSYNC_buff_I_0.BUFFER_0__i2C_net ;
    wire \receive_module.rx_counter.X_8 ;
    wire \receive_module.rx_counter.X_9 ;
    wire \receive_module.rx_counter.n3630 ;
    wire \TVP_VSYNC_buff_I_0.BUFFER_1_0 ;
    wire \INVTVP_VSYNC_buff_I_0.WIRE_OUT_0__9C_net ;
    wire \line_buffer.n467 ;
    wire \receive_module.rx_counter.n4_cascade_ ;
    wire \receive_module.rx_counter.n3400 ;
    wire \line_buffer.n565 ;
    wire \receive_module.rx_counter.X_5 ;
    wire \receive_module.rx_counter.X_4 ;
    wire \receive_module.rx_counter.X_3 ;
    wire \receive_module.rx_counter.X_6 ;
    wire \receive_module.rx_counter.n6_cascade_ ;
    wire \receive_module.rx_counter.X_7 ;
    wire \receive_module.rx_counter.n3385 ;
    wire \receive_module.rx_counter.old_HS ;
    wire TVP_HSYNC_buff;
    wire bfn_12_11_0_;
    wire \receive_module.n3091 ;
    wire \receive_module.n3092 ;
    wire \receive_module.n3093 ;
    wire \receive_module.n3094 ;
    wire \receive_module.n3095 ;
    wire \receive_module.n3096 ;
    wire \receive_module.n3097 ;
    wire \receive_module.n3098 ;
    wire bfn_12_12_0_;
    wire \receive_module.n3099 ;
    wire \receive_module.n3100 ;
    wire \receive_module.n3101 ;
    wire \receive_module.n3102 ;
    wire \receive_module.n3103 ;
    wire \receive_module.n3632 ;
    wire \transmit_module.Y_DELTA_PATTERN_53 ;
    wire \transmit_module.Y_DELTA_PATTERN_52 ;
    wire \transmit_module.Y_DELTA_PATTERN_56 ;
    wire \transmit_module.Y_DELTA_PATTERN_55 ;
    wire \transmit_module.Y_DELTA_PATTERN_54 ;
    wire \transmit_module.video_signal_controller.n3629_cascade_ ;
    wire \transmit_module.video_signal_controller.n2901 ;
    wire bfn_12_15_0_;
    wire \transmit_module.video_signal_controller.n3125 ;
    wire \transmit_module.video_signal_controller.n3126 ;
    wire \transmit_module.video_signal_controller.n3127 ;
    wire \transmit_module.video_signal_controller.n3128 ;
    wire \transmit_module.video_signal_controller.n3129 ;
    wire \transmit_module.video_signal_controller.n3130 ;
    wire \transmit_module.video_signal_controller.n3131 ;
    wire \transmit_module.video_signal_controller.n3132 ;
    wire bfn_12_16_0_;
    wire \transmit_module.video_signal_controller.n3133 ;
    wire \transmit_module.video_signal_controller.n3134 ;
    wire \transmit_module.video_signal_controller.n3135 ;
    wire \transmit_module.Y_DELTA_PATTERN_2 ;
    wire \transmit_module.Y_DELTA_PATTERN_3 ;
    wire \transmit_module.Y_DELTA_PATTERN_5 ;
    wire \transmit_module.Y_DELTA_PATTERN_4 ;
    wire \transmit_module.Y_DELTA_PATTERN_7 ;
    wire \transmit_module.Y_DELTA_PATTERN_6 ;
    wire \receive_module.n131 ;
    wire RX_ADDR_5;
    wire \receive_module.n130 ;
    wire RX_ADDR_6;
    wire \receive_module.n129 ;
    wire RX_ADDR_7;
    wire \receive_module.n128 ;
    wire RX_ADDR_8;
    wire \receive_module.n127 ;
    wire RX_ADDR_9;
    wire \receive_module.n136 ;
    wire RX_ADDR_0;
    wire \receive_module.n135 ;
    wire RX_ADDR_1;
    wire \line_buffer.n593 ;
    wire \line_buffer.n585 ;
    wire \receive_module.n126 ;
    wire RX_ADDR_10;
    wire \receive_module.n133 ;
    wire RX_ADDR_3;
    wire \receive_module.n132 ;
    wire RX_ADDR_4;
    wire \tvp_video_buffer.BUFFER_1_2 ;
    wire RX_DATA_0;
    wire bfn_13_6_0_;
    wire \receive_module.rx_counter.n3156 ;
    wire \receive_module.rx_counter.n3157 ;
    wire \receive_module.rx_counter.n3158 ;
    wire \receive_module.rx_counter.n3159 ;
    wire \receive_module.rx_counter.n3160 ;
    wire \receive_module.rx_counter.n3623 ;
    wire \receive_module.rx_counter.FRAME_COUNTER_4 ;
    wire \receive_module.rx_counter.FRAME_COUNTER_2 ;
    wire \receive_module.rx_counter.FRAME_COUNTER_5 ;
    wire \receive_module.rx_counter.FRAME_COUNTER_1 ;
    wire \receive_module.rx_counter.FRAME_COUNTER_0 ;
    wire \receive_module.rx_counter.FRAME_COUNTER_3 ;
    wire \receive_module.rx_counter.n3473_cascade_ ;
    wire \receive_module.rx_counter.n7 ;
    wire \receive_module.rx_counter.n11 ;
    wire \receive_module.rx_counter.old_VS ;
    wire \receive_module.rx_counter.n11_cascade_ ;
    wire \receive_module.rx_counter.n2529 ;
    wire \receive_module.rx_counter.n4_adj_605 ;
    wire \receive_module.rx_counter.n3422_cascade_ ;
    wire \receive_module.rx_counter.n55_adj_606 ;
    wire \receive_module.rx_counter.n3394 ;
    wire \receive_module.rx_counter.n5 ;
    wire \receive_module.rx_counter.n3413 ;
    wire \line_buffer.n596 ;
    wire \receive_module.rx_counter.n4_adj_604 ;
    wire bfn_13_9_0_;
    wire \receive_module.rx_counter.n3117 ;
    wire \receive_module.rx_counter.n3118 ;
    wire \receive_module.rx_counter.n3119 ;
    wire \receive_module.rx_counter.n3120 ;
    wire \receive_module.rx_counter.Y_5 ;
    wire \receive_module.rx_counter.n3121 ;
    wire \receive_module.rx_counter.Y_6 ;
    wire \receive_module.rx_counter.n3122 ;
    wire \receive_module.rx_counter.n3123 ;
    wire \receive_module.rx_counter.n3124 ;
    wire bfn_13_10_0_;
    wire \receive_module.rx_counter.n2063 ;
    wire \receive_module.n134 ;
    wire TVP_VSYNC_buff;
    wire RX_ADDR_2;
    wire \receive_module.n3631 ;
    wire bfn_13_12_0_;
    wire \transmit_module.video_signal_controller.n3136 ;
    wire \transmit_module.video_signal_controller.n3137 ;
    wire \transmit_module.video_signal_controller.n3138 ;
    wire \transmit_module.video_signal_controller.n3139 ;
    wire \transmit_module.video_signal_controller.n3140 ;
    wire \transmit_module.video_signal_controller.n3141 ;
    wire \transmit_module.video_signal_controller.n3142 ;
    wire \transmit_module.video_signal_controller.n3143 ;
    wire bfn_13_13_0_;
    wire \transmit_module.video_signal_controller.n3144 ;
    wire \transmit_module.video_signal_controller.n3145 ;
    wire \transmit_module.video_signal_controller.n3146 ;
    wire \line_buffer.n564 ;
    wire \transmit_module.video_signal_controller.n3624 ;
    wire \transmit_module.video_signal_controller.VGA_X_2 ;
    wire \transmit_module.video_signal_controller.VGA_X_1 ;
    wire \transmit_module.video_signal_controller.VGA_X_0 ;
    wire \transmit_module.video_signal_controller.n2001 ;
    wire \transmit_module.video_signal_controller.n2917_cascade_ ;
    wire \transmit_module.video_signal_controller.n3313 ;
    wire \transmit_module.video_signal_controller.n2947_cascade_ ;
    wire \line_buffer.n522 ;
    wire \line_buffer.n530 ;
    wire \transmit_module.video_signal_controller.VGA_X_3 ;
    wire \transmit_module.video_signal_controller.VGA_X_5 ;
    wire \transmit_module.video_signal_controller.n18 ;
    wire \transmit_module.video_signal_controller.VGA_X_9 ;
    wire \transmit_module.video_signal_controller.VGA_X_10 ;
    wire \transmit_module.video_signal_controller.n4 ;
    wire \transmit_module.video_signal_controller.VGA_X_7 ;
    wire \transmit_module.video_signal_controller.n3625_cascade_ ;
    wire \transmit_module.video_signal_controller.VGA_X_4 ;
    wire \line_buffer.n597 ;
    wire \line_buffer.n594 ;
    wire \line_buffer.n586 ;
    wire \line_buffer.n3591 ;
    wire \line_buffer.n468 ;
    wire n25;
    wire \transmit_module.ADDR_Y_COMPONENT_3 ;
    wire \tvp_video_buffer.BUFFER_0_4 ;
    wire \receive_module.rx_counter.Y_4 ;
    wire \receive_module.rx_counter.Y_7 ;
    wire \receive_module.rx_counter.Y_1 ;
    wire \receive_module.rx_counter.Y_3 ;
    wire \receive_module.rx_counter.Y_2 ;
    wire \receive_module.rx_counter.Y_8 ;
    wire \receive_module.rx_counter.n10_adj_610 ;
    wire \receive_module.rx_counter.Y_0 ;
    wire \receive_module.rx_counter.n14_cascade_ ;
    wire \receive_module.rx_counter.n3633 ;
    wire RX_TX_SYNC;
    wire \sync_buffer.BUFFER_0_0 ;
    wire RX_ADDR_12;
    wire RX_WE;
    wire RX_ADDR_13;
    wire RX_ADDR_11;
    wire \line_buffer.n532 ;
    wire \tvp_video_buffer.BUFFER_1_3 ;
    wire RX_DATA_1;
    wire \sync_buffer.BUFFER_1_0 ;
    wire RX_TX_SYNC_BUFF;
    wire \transmit_module.video_signal_controller.n2036 ;
    wire \transmit_module.video_signal_controller.n2378 ;
    wire \transmit_module.video_signal_controller.n49_cascade_ ;
    wire \transmit_module.video_signal_controller.VGA_Y_1 ;
    wire \transmit_module.video_signal_controller.VGA_Y_0 ;
    wire \transmit_module.n113 ;
    wire \transmit_module.n142_cascade_ ;
    wire \transmit_module.video_signal_controller.n45 ;
    wire \transmit_module.video_signal_controller.n3412 ;
    wire \transmit_module.video_signal_controller.VGA_Y_8 ;
    wire \transmit_module.video_signal_controller.VGA_Y_7 ;
    wire \transmit_module.video_signal_controller.n3626 ;
    wire \transmit_module.video_signal_controller.VGA_Y_6 ;
    wire \transmit_module.video_signal_controller.n3626_cascade_ ;
    wire \transmit_module.video_signal_controller.VGA_Y_11 ;
    wire \transmit_module.n137_cascade_ ;
    wire \transmit_module.video_signal_controller.VGA_Y_5 ;
    wire \transmit_module.video_signal_controller.VGA_Y_3 ;
    wire \transmit_module.video_signal_controller.VGA_Y_4 ;
    wire \transmit_module.video_signal_controller.n3628 ;
    wire \transmit_module.video_signal_controller.VGA_Y_9 ;
    wire \transmit_module.video_signal_controller.n3331 ;
    wire \transmit_module.video_signal_controller.n7_adj_618_cascade_ ;
    wire \transmit_module.video_signal_controller.n3622 ;
    wire \transmit_module.video_signal_controller.VGA_VISIBLE_N_580_cascade_ ;
    wire \transmit_module.video_signal_controller.VGA_Y_10 ;
    wire \transmit_module.video_signal_controller.n3477 ;
    wire \transmit_module.video_signal_controller.n16 ;
    wire \transmit_module.video_signal_controller.VGA_Y_2 ;
    wire \transmit_module.video_signal_controller.VGA_X_8 ;
    wire \transmit_module.video_signal_controller.n3471 ;
    wire \transmit_module.video_signal_controller.n4_adj_617 ;
    wire \transmit_module.video_signal_controller.VGA_X_6 ;
    wire \transmit_module.n144 ;
    wire \transmit_module.n3636 ;
    wire \transmit_module.ADDR_Y_COMPONENT_0 ;
    wire \transmit_module.old_VGA_HS ;
    wire \transmit_module.VGA_VISIBLE_Y ;
    wire ADV_HSYNC_c;
    wire \transmit_module.n137 ;
    wire n18;
    wire \transmit_module.n116 ;
    wire \transmit_module.n147 ;
    wire n28;
    wire \transmit_module.n115 ;
    wire \transmit_module.n146 ;
    wire n27;
    wire DEBUG_c_3_c;
    wire DEBUG_c_4_c;
    wire DEBUG_c_5_c;
    wire \tvp_video_buffer.BUFFER_0_7 ;
    wire \transmit_module.TX_ADDR_0 ;
    wire \transmit_module.n132 ;
    wire bfn_15_13_0_;
    wire \transmit_module.n131 ;
    wire \transmit_module.n3104 ;
    wire \transmit_module.n3105 ;
    wire \transmit_module.TX_ADDR_3 ;
    wire \transmit_module.n129 ;
    wire \transmit_module.n3106 ;
    wire \transmit_module.n3107 ;
    wire \transmit_module.n127 ;
    wire \transmit_module.n3108 ;
    wire \transmit_module.n3109 ;
    wire \transmit_module.n3110 ;
    wire \transmit_module.n3111 ;
    wire bfn_15_14_0_;
    wire \transmit_module.n3112 ;
    wire \transmit_module.n122 ;
    wire \transmit_module.n3113 ;
    wire \transmit_module.n3114 ;
    wire \transmit_module.n3115 ;
    wire \transmit_module.n3116 ;
    wire \transmit_module.ADDR_Y_COMPONENT_5 ;
    wire \transmit_module.TX_ADDR_5 ;
    wire \transmit_module.n111 ;
    wire \transmit_module.n111_cascade_ ;
    wire \transmit_module.n142 ;
    wire n23;
    wire \transmit_module.video_signal_controller.VGA_VISIBLE_N_580 ;
    wire \transmit_module.video_signal_controller.n3333 ;
    wire \transmit_module.video_signal_controller.VGA_X_11 ;
    wire \transmit_module.video_signal_controller.n7 ;
    wire \transmit_module.ADDR_Y_COMPONENT_10 ;
    wire \transmit_module.TX_ADDR_10 ;
    wire \transmit_module.n106 ;
    wire \transmit_module.n120 ;
    wire \transmit_module.n121 ;
    wire \transmit_module.n119 ;
    wire \transmit_module.n2057 ;
    wire \transmit_module.n124 ;
    wire \transmit_module.n126 ;
    wire \transmit_module.n123 ;
    wire \transmit_module.n125 ;
    wire n22;
    wire \transmit_module.ADDR_Y_COMPONENT_8 ;
    wire \transmit_module.TX_ADDR_8 ;
    wire n21;
    wire \transmit_module.TX_ADDR_1 ;
    wire \transmit_module.ADDR_Y_COMPONENT_1 ;
    wire \transmit_module.n128 ;
    wire \transmit_module.n143 ;
    wire CONSTANT_ONE_NET;
    wire RX_DATA_3;
    wire \tvp_video_buffer.BUFFER_0_5 ;
    wire \tvp_video_buffer.BUFFER_1_5 ;
    wire \tvp_video_buffer.BUFFER_0_6 ;
    wire \tvp_video_buffer.BUFFER_1_6 ;
    wire RX_DATA_4;
    wire \tvp_video_buffer.BUFFER_1_7 ;
    wire RX_DATA_5;
    wire RX_DATA_6;
    wire DEBUG_c_6_c;
    wire \tvp_video_buffer.BUFFER_0_8 ;
    wire \tvp_video_buffer.BUFFER_1_8 ;
    wire \transmit_module.n141 ;
    wire \transmit_module.n2167 ;
    wire \transmit_module.n140 ;
    wire \transmit_module.n130 ;
    wire \transmit_module.n145_cascade_ ;
    wire \transmit_module.Y_DELTA_PATTERN_16 ;
    wire \transmit_module.Y_DELTA_PATTERN_17 ;
    wire \transmit_module.Y_DELTA_PATTERN_20 ;
    wire \transmit_module.Y_DELTA_PATTERN_19 ;
    wire \transmit_module.Y_DELTA_PATTERN_18 ;
    wire \transmit_module.ADDR_Y_COMPONENT_13 ;
    wire \transmit_module.ADDR_Y_COMPONENT_12 ;
    wire \transmit_module.ADDR_Y_COMPONENT_11 ;
    wire \transmit_module.Y_DELTA_PATTERN_1 ;
    wire \transmit_module.n108 ;
    wire \transmit_module.n139 ;
    wire n20;
    wire \transmit_module.ADDR_Y_COMPONENT_7 ;
    wire \transmit_module.TX_ADDR_7 ;
    wire \transmit_module.n109 ;
    wire \transmit_module.ADDR_Y_COMPONENT_6 ;
    wire \transmit_module.TX_ADDR_6 ;
    wire \transmit_module.n110 ;
    wire \transmit_module.ADDR_Y_COMPONENT_2 ;
    wire \transmit_module.TX_ADDR_2 ;
    wire \transmit_module.ADDR_Y_COMPONENT_9 ;
    wire \transmit_module.TX_ADDR_9 ;
    wire \transmit_module.n107 ;
    wire \transmit_module.n107_cascade_ ;
    wire \transmit_module.n138 ;
    wire n19;
    wire \transmit_module.n114 ;
    wire \transmit_module.n145 ;
    wire n26;
    wire \tvp_video_buffer.BUFFER_1_4 ;
    wire RX_DATA_2;
    wire \transmit_module.X_DELTA_PATTERN_0 ;
    wire \transmit_module.X_DELTA_PATTERN_10 ;
    wire \transmit_module.X_DELTA_PATTERN_15 ;
    wire \transmit_module.X_DELTA_PATTERN_14 ;
    wire \transmit_module.X_DELTA_PATTERN_13 ;
    wire \transmit_module.X_DELTA_PATTERN_12 ;
    wire \transmit_module.X_DELTA_PATTERN_11 ;
    wire \transmit_module.X_DELTA_PATTERN_9 ;
    wire \transmit_module.X_DELTA_PATTERN_8 ;
    wire \transmit_module.n3627 ;
    wire \line_buffer.n556 ;
    wire \line_buffer.n548 ;
    wire \transmit_module.Y_DELTA_PATTERN_0 ;
    wire \transmit_module.n112 ;
    wire \transmit_module.TX_ADDR_4 ;
    wire \transmit_module.ADDR_Y_COMPONENT_4 ;
    wire \transmit_module.n2069 ;
    wire ADV_VSYNC_c;
    wire \line_buffer.n529 ;
    wire \line_buffer.n521 ;
    wire \line_buffer.n3500_cascade_ ;
    wire \line_buffer.n3501 ;
    wire \line_buffer.n3537_cascade_ ;
    wire \line_buffer.n464 ;
    wire \line_buffer.n456 ;
    wire \line_buffer.n3497 ;
    wire \line_buffer.n524 ;
    wire \line_buffer.n516 ;
    wire \line_buffer.n560 ;
    wire \line_buffer.n552 ;
    wire \transmit_module.X_DELTA_PATTERN_1 ;
    wire \transmit_module.X_DELTA_PATTERN_2 ;
    wire \transmit_module.X_DELTA_PATTERN_3 ;
    wire \transmit_module.X_DELTA_PATTERN_5 ;
    wire \transmit_module.X_DELTA_PATTERN_4 ;
    wire \transmit_module.X_DELTA_PATTERN_7 ;
    wire \transmit_module.X_DELTA_PATTERN_6 ;
    wire \transmit_module.n2115 ;
    wire \transmit_module.n3635 ;
    wire \line_buffer.n463 ;
    wire \line_buffer.n455 ;
    wire \line_buffer.n3525 ;
    wire \line_buffer.n3524_cascade_ ;
    wire \line_buffer.n3521 ;
    wire \line_buffer.n3555_cascade_ ;
    wire \line_buffer.n3519 ;
    wire \line_buffer.n561 ;
    wire \line_buffer.n553 ;
    wire \line_buffer.n3498 ;
    wire \line_buffer.n587 ;
    wire \line_buffer.n579 ;
    wire n1814;
    wire TX_DATA_1;
    wire n1813;
    wire TX_DATA_5;
    wire n1809;
    wire TX_DATA_6;
    wire n1808;
    wire \line_buffer.n528 ;
    wire \line_buffer.n520 ;
    wire \line_buffer.n3594 ;
    wire \line_buffer.n592 ;
    wire \line_buffer.n584 ;
    wire \line_buffer.n3489 ;
    wire \line_buffer.n3488 ;
    wire \line_buffer.n3561 ;
    wire \line_buffer.n591 ;
    wire \line_buffer.n583 ;
    wire \line_buffer.n523 ;
    wire \line_buffer.n515 ;
    wire \line_buffer.n3597 ;
    wire \line_buffer.n3600_cascade_ ;
    wire TX_DATA_0;
    wire \transmit_module.VGA_VISIBLE ;
    wire TX_DATA_7;
    wire ADV_B_c;
    wire RX_DATA_7;
    wire \line_buffer.n465 ;
    wire \line_buffer.n457 ;
    wire \line_buffer.n3588 ;
    wire \line_buffer.n557 ;
    wire \line_buffer.n549 ;
    wire \line_buffer.n460 ;
    wire \line_buffer.n452 ;
    wire \line_buffer.n3549 ;
    wire \line_buffer.n3552_cascade_ ;
    wire \line_buffer.n527 ;
    wire \line_buffer.n519 ;
    wire \line_buffer.n3573 ;
    wire \line_buffer.n589 ;
    wire \line_buffer.n581 ;
    wire \line_buffer.n517 ;
    wire \line_buffer.n525 ;
    wire \line_buffer.n3603_cascade_ ;
    wire \line_buffer.n3606 ;
    wire \line_buffer.n462 ;
    wire \line_buffer.n454 ;
    wire \line_buffer.n3546_cascade_ ;
    wire \line_buffer.n3576 ;
    wire \line_buffer.n555 ;
    wire \line_buffer.n547 ;
    wire \line_buffer.n461 ;
    wire \line_buffer.n453 ;
    wire \line_buffer.n588 ;
    wire \line_buffer.n580 ;
    wire \line_buffer.n3522 ;
    wire \line_buffer.n458 ;
    wire \line_buffer.n450 ;
    wire \line_buffer.n3579 ;
    wire \line_buffer.n3582 ;
    wire TX_DATA_2;
    wire n1812;
    wire TX_DATA_4;
    wire n1810;
    wire \line_buffer.n554 ;
    wire \line_buffer.n562 ;
    wire \line_buffer.n3585 ;
    wire \line_buffer.n558 ;
    wire \line_buffer.n550 ;
    wire TX_ADDR_13;
    wire \line_buffer.n3482 ;
    wire \line_buffer.n3567_cascade_ ;
    wire \line_buffer.n3483 ;
    wire \line_buffer.n559 ;
    wire TX_ADDR_12;
    wire \line_buffer.n551 ;
    wire \line_buffer.n3543 ;
    wire \line_buffer.n582 ;
    wire \line_buffer.n590 ;
    wire \line_buffer.n3480 ;
    wire TX_DATA_3;
    wire n1811;
    wire ADV_CLK_c;
    wire \transmit_module.n2367 ;
    wire \tvp_video_buffer.BUFFER_1_9 ;
    wire \line_buffer.n526 ;
    wire \line_buffer.n518 ;
    wire \line_buffer.n3479 ;
    wire DEBUG_c_7_c;
    wire \tvp_video_buffer.BUFFER_0_9 ;
    wire DEBUG_c_2_c;
    wire \line_buffer.n459 ;
    wire \line_buffer.n451 ;
    wire TX_ADDR_11;
    wire \line_buffer.n3518 ;
    wire _gnd_net_;

    defparam \tx_pll.TX_PLL_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \tx_pll.TX_PLL_inst .TEST_MODE=1'b0;
    defparam \tx_pll.TX_PLL_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \tx_pll.TX_PLL_inst .PLLOUT_SELECT="GENCLK";
    defparam \tx_pll.TX_PLL_inst .FILTER_RANGE=3'b010;
    defparam \tx_pll.TX_PLL_inst .FEEDBACK_PATH="SIMPLE";
    defparam \tx_pll.TX_PLL_inst .FDA_RELATIVE=4'b0000;
    defparam \tx_pll.TX_PLL_inst .FDA_FEEDBACK=4'b0000;
    defparam \tx_pll.TX_PLL_inst .ENABLE_ICEGATE=1'b0;
    defparam \tx_pll.TX_PLL_inst .DIVR=4'b0000;
    defparam \tx_pll.TX_PLL_inst .DIVQ=3'b100;
    defparam \tx_pll.TX_PLL_inst .DIVF=7'b0100110;
    defparam \tx_pll.TX_PLL_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \tx_pll.TX_PLL_inst  (
            .EXTFEEDBACK(),
            .LATCHINPUTVALUE(),
            .SCLK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(ADV_CLK_c),
            .REFERENCECLK(N__8399),
            .RESETB(N__18070),
            .BYPASS(GNDG0),
            .SDI(),
            .DYNAMICDELAY({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7}),
            .PLLOUTGLOBAL());
    defparam \line_buffer.mem2_physical .WRITE_MODE=3;
    defparam \line_buffer.mem2_physical .READ_MODE=3;
    defparam \line_buffer.mem2_physical .INIT_F=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem2_physical .INIT_E=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem2_physical .INIT_D=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem2_physical .INIT_C=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem2_physical .INIT_B=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem2_physical .INIT_A=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem2_physical .INIT_9=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem2_physical .INIT_8=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem2_physical .INIT_7=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem2_physical .INIT_6=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem2_physical .INIT_5=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem2_physical .INIT_4=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem2_physical .INIT_3=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem2_physical .INIT_2=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem2_physical .INIT_1=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem2_physical .INIT_0=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    SB_RAM40_4K \line_buffer.mem2_physical  (
            .RDATA({dangling_wire_8,dangling_wire_9,dangling_wire_10,dangling_wire_11,\line_buffer.n465 ,dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,\line_buffer.n464 ,dangling_wire_19,dangling_wire_20,dangling_wire_21}),
            .RADDR({N__16186,N__18964,N__19420,N__17104,N__17374,N__16837,N__9121,N__14008,N__18712,N__15670,N__15922}),
            .WADDR({N__12349,N__10438,N__10681,N__10936,N__11194,N__11452,N__11833,N__12091,N__12892,N__9922,N__10183}),
            .MASK({dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29,dangling_wire_30,dangling_wire_31,dangling_wire_32,dangling_wire_33,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37}),
            .WDATA({dangling_wire_38,dangling_wire_39,dangling_wire_40,dangling_wire_41,N__22154,dangling_wire_42,dangling_wire_43,dangling_wire_44,dangling_wire_45,dangling_wire_46,dangling_wire_47,dangling_wire_48,N__18559,dangling_wire_49,dangling_wire_50,dangling_wire_51}),
            .RCLKE(),
            .RCLK(N__23228),
            .RE(N__18072),
            .WCLKE(),
            .WCLK(N__24625),
            .WE(N__14183));
    defparam \line_buffer.mem14_physical .WRITE_MODE=3;
    defparam \line_buffer.mem14_physical .READ_MODE=3;
    defparam \line_buffer.mem14_physical .INIT_F=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem14_physical .INIT_E=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem14_physical .INIT_D=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem14_physical .INIT_C=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem14_physical .INIT_B=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem14_physical .INIT_A=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem14_physical .INIT_9=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem14_physical .INIT_8=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem14_physical .INIT_7=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem14_physical .INIT_6=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem14_physical .INIT_5=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem14_physical .INIT_4=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem14_physical .INIT_3=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    defparam \line_buffer.mem14_physical .INIT_2=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    defparam \line_buffer.mem14_physical .INIT_1=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    defparam \line_buffer.mem14_physical .INIT_0=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    SB_RAM40_4K \line_buffer.mem14_physical  (
            .RDATA({dangling_wire_52,dangling_wire_53,dangling_wire_54,dangling_wire_55,\line_buffer.n552 ,dangling_wire_56,dangling_wire_57,dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,\line_buffer.n551 ,dangling_wire_63,dangling_wire_64,dangling_wire_65}),
            .RADDR({N__16258,N__19036,N__19492,N__17176,N__17446,N__16909,N__9193,N__14080,N__18784,N__15742,N__15994}),
            .WADDR({N__12421,N__10510,N__10753,N__11008,N__11266,N__11524,N__11905,N__12163,N__12964,N__9994,N__10255}),
            .MASK({dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73,dangling_wire_74,dangling_wire_75,dangling_wire_76,dangling_wire_77,dangling_wire_78,dangling_wire_79,dangling_wire_80,dangling_wire_81}),
            .WDATA({dangling_wire_82,dangling_wire_83,dangling_wire_84,dangling_wire_85,N__17671,dangling_wire_86,dangling_wire_87,dangling_wire_88,dangling_wire_89,dangling_wire_90,dangling_wire_91,dangling_wire_92,N__17762,dangling_wire_93,dangling_wire_94,dangling_wire_95}),
            .RCLKE(),
            .RCLK(N__23483),
            .RE(N__18170),
            .WCLKE(),
            .WCLK(N__24611),
            .WE(N__13374));
    defparam \line_buffer.mem5_physical .WRITE_MODE=3;
    defparam \line_buffer.mem5_physical .READ_MODE=3;
    defparam \line_buffer.mem5_physical .INIT_F=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem5_physical .INIT_E=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem5_physical .INIT_D=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem5_physical .INIT_C=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem5_physical .INIT_B=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem5_physical .INIT_A=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem5_physical .INIT_9=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem5_physical .INIT_8=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem5_physical .INIT_7=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem5_physical .INIT_6=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem5_physical .INIT_5=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem5_physical .INIT_4=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem5_physical .INIT_3=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    defparam \line_buffer.mem5_physical .INIT_2=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    defparam \line_buffer.mem5_physical .INIT_1=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    defparam \line_buffer.mem5_physical .INIT_0=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    SB_RAM40_4K \line_buffer.mem5_physical  (
            .RDATA({dangling_wire_96,dangling_wire_97,dangling_wire_98,dangling_wire_99,\line_buffer.n562 ,dangling_wire_100,dangling_wire_101,dangling_wire_102,dangling_wire_103,dangling_wire_104,dangling_wire_105,dangling_wire_106,\line_buffer.n561 ,dangling_wire_107,dangling_wire_108,dangling_wire_109}),
            .RADDR({N__16189,N__18985,N__19435,N__17113,N__17377,N__16840,N__9124,N__13999,N__18721,N__15679,N__15937}),
            .WADDR({N__12340,N__10441,N__10696,N__10945,N__11203,N__11467,N__11830,N__12088,N__12913,N__9937,N__10192}),
            .MASK({dangling_wire_110,dangling_wire_111,dangling_wire_112,dangling_wire_113,dangling_wire_114,dangling_wire_115,dangling_wire_116,dangling_wire_117,dangling_wire_118,dangling_wire_119,dangling_wire_120,dangling_wire_121,dangling_wire_122,dangling_wire_123,dangling_wire_124,dangling_wire_125}),
            .WDATA({dangling_wire_126,dangling_wire_127,dangling_wire_128,dangling_wire_129,N__22148,dangling_wire_130,dangling_wire_131,dangling_wire_132,dangling_wire_133,dangling_wire_134,dangling_wire_135,dangling_wire_136,N__18561,dangling_wire_137,dangling_wire_138,dangling_wire_139}),
            .RCLKE(),
            .RCLK(N__22710),
            .RE(N__18051),
            .WCLKE(),
            .WCLK(N__24624),
            .WE(N__9647));
    defparam \line_buffer.mem11_physical .WRITE_MODE=3;
    defparam \line_buffer.mem11_physical .READ_MODE=3;
    defparam \line_buffer.mem11_physical .INIT_F=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem11_physical .INIT_E=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem11_physical .INIT_D=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem11_physical .INIT_C=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem11_physical .INIT_B=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem11_physical .INIT_A=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem11_physical .INIT_9=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem11_physical .INIT_8=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem11_physical .INIT_7=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem11_physical .INIT_6=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem11_physical .INIT_5=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem11_physical .INIT_4=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem11_physical .INIT_3=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem11_physical .INIT_2=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem11_physical .INIT_1=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem11_physical .INIT_0=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    SB_RAM40_4K \line_buffer.mem11_physical  (
            .RDATA({dangling_wire_140,dangling_wire_141,dangling_wire_142,dangling_wire_143,\line_buffer.n520 ,dangling_wire_144,dangling_wire_145,dangling_wire_146,dangling_wire_147,dangling_wire_148,dangling_wire_149,dangling_wire_150,\line_buffer.n519 ,dangling_wire_151,dangling_wire_152,dangling_wire_153}),
            .RADDR({N__16294,N__19072,N__19528,N__17212,N__17482,N__16945,N__9229,N__14116,N__18820,N__15778,N__16030}),
            .WADDR({N__12457,N__10546,N__10789,N__11044,N__11302,N__11560,N__11941,N__12199,N__13000,N__10030,N__10291}),
            .MASK({dangling_wire_154,dangling_wire_155,dangling_wire_156,dangling_wire_157,dangling_wire_158,dangling_wire_159,dangling_wire_160,dangling_wire_161,dangling_wire_162,dangling_wire_163,dangling_wire_164,dangling_wire_165,dangling_wire_166,dangling_wire_167,dangling_wire_168,dangling_wire_169}),
            .WDATA({dangling_wire_170,dangling_wire_171,dangling_wire_172,dangling_wire_173,N__17654,dangling_wire_174,dangling_wire_175,dangling_wire_176,dangling_wire_177,dangling_wire_178,dangling_wire_179,dangling_wire_180,N__17761,dangling_wire_181,dangling_wire_182,dangling_wire_183}),
            .RCLKE(),
            .RCLK(N__23320),
            .RE(N__18197),
            .WCLKE(),
            .WCLK(N__24601),
            .WE(N__14395));
    defparam \line_buffer.mem21_physical .WRITE_MODE=3;
    defparam \line_buffer.mem21_physical .READ_MODE=3;
    defparam \line_buffer.mem21_physical .INIT_F=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem21_physical .INIT_E=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem21_physical .INIT_D=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem21_physical .INIT_C=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem21_physical .INIT_B=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem21_physical .INIT_A=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem21_physical .INIT_9=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem21_physical .INIT_8=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem21_physical .INIT_7=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem21_physical .INIT_6=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem21_physical .INIT_5=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem21_physical .INIT_4=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem21_physical .INIT_3=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem21_physical .INIT_2=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem21_physical .INIT_1=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem21_physical .INIT_0=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    SB_RAM40_4K \line_buffer.mem21_physical  (
            .RDATA({dangling_wire_184,dangling_wire_185,dangling_wire_186,dangling_wire_187,\line_buffer.n582 ,dangling_wire_188,dangling_wire_189,dangling_wire_190,dangling_wire_191,dangling_wire_192,dangling_wire_193,dangling_wire_194,\line_buffer.n581 ,dangling_wire_195,dangling_wire_196,dangling_wire_197}),
            .RADDR({N__16162,N__18940,N__19396,N__17080,N__17350,N__16813,N__9097,N__13984,N__18688,N__15646,N__15898}),
            .WADDR({N__12325,N__10414,N__10657,N__10912,N__11170,N__11428,N__11809,N__12067,N__12868,N__9898,N__10159}),
            .MASK({dangling_wire_198,dangling_wire_199,dangling_wire_200,dangling_wire_201,dangling_wire_202,dangling_wire_203,dangling_wire_204,dangling_wire_205,dangling_wire_206,dangling_wire_207,dangling_wire_208,dangling_wire_209,dangling_wire_210,dangling_wire_211,dangling_wire_212,dangling_wire_213}),
            .WDATA({dangling_wire_214,dangling_wire_215,dangling_wire_216,dangling_wire_217,N__17911,dangling_wire_218,dangling_wire_219,dangling_wire_220,dangling_wire_221,dangling_wire_222,dangling_wire_223,dangling_wire_224,N__19755,dangling_wire_225,dangling_wire_226,dangling_wire_227}),
            .RCLKE(),
            .RCLK(N__23057),
            .RE(N__18089),
            .WCLKE(),
            .WCLK(N__24631),
            .WE(N__12691));
    defparam \line_buffer.mem12_physical .WRITE_MODE=3;
    defparam \line_buffer.mem12_physical .READ_MODE=3;
    defparam \line_buffer.mem12_physical .INIT_F=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem12_physical .INIT_E=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem12_physical .INIT_D=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem12_physical .INIT_C=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem12_physical .INIT_B=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem12_physical .INIT_A=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem12_physical .INIT_9=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem12_physical .INIT_8=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem12_physical .INIT_7=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem12_physical .INIT_6=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem12_physical .INIT_5=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem12_physical .INIT_4=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem12_physical .INIT_3=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem12_physical .INIT_2=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem12_physical .INIT_1=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem12_physical .INIT_0=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    SB_RAM40_4K \line_buffer.mem12_physical  (
            .RDATA({dangling_wire_228,dangling_wire_229,dangling_wire_230,dangling_wire_231,\line_buffer.n518 ,dangling_wire_232,dangling_wire_233,dangling_wire_234,dangling_wire_235,dangling_wire_236,dangling_wire_237,dangling_wire_238,\line_buffer.n517 ,dangling_wire_239,dangling_wire_240,dangling_wire_241}),
            .RADDR({N__16282,N__19060,N__19516,N__17200,N__17470,N__16933,N__9217,N__14104,N__18808,N__15766,N__16018}),
            .WADDR({N__12445,N__10534,N__10777,N__11032,N__11290,N__11548,N__11929,N__12187,N__12988,N__10018,N__10279}),
            .MASK({dangling_wire_242,dangling_wire_243,dangling_wire_244,dangling_wire_245,dangling_wire_246,dangling_wire_247,dangling_wire_248,dangling_wire_249,dangling_wire_250,dangling_wire_251,dangling_wire_252,dangling_wire_253,dangling_wire_254,dangling_wire_255,dangling_wire_256,dangling_wire_257}),
            .WDATA({dangling_wire_258,dangling_wire_259,dangling_wire_260,dangling_wire_261,N__17886,dangling_wire_262,dangling_wire_263,dangling_wire_264,dangling_wire_265,dangling_wire_266,dangling_wire_267,dangling_wire_268,N__19742,dangling_wire_269,dangling_wire_270,dangling_wire_271}),
            .RCLKE(),
            .RCLK(N__23169),
            .RE(N__18196),
            .WCLKE(),
            .WCLK(N__24606),
            .WE(N__14393));
    defparam \line_buffer.mem24_physical .WRITE_MODE=3;
    defparam \line_buffer.mem24_physical .READ_MODE=3;
    defparam \line_buffer.mem24_physical .INIT_F=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem24_physical .INIT_E=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem24_physical .INIT_D=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem24_physical .INIT_C=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem24_physical .INIT_B=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem24_physical .INIT_A=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem24_physical .INIT_9=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem24_physical .INIT_8=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem24_physical .INIT_7=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem24_physical .INIT_6=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem24_physical .INIT_5=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem24_physical .INIT_4=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem24_physical .INIT_3=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem24_physical .INIT_2=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem24_physical .INIT_1=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem24_physical .INIT_0=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    SB_RAM40_4K \line_buffer.mem24_physical  (
            .RDATA({dangling_wire_272,dangling_wire_273,dangling_wire_274,dangling_wire_275,\line_buffer.n526 ,dangling_wire_276,dangling_wire_277,dangling_wire_278,dangling_wire_279,dangling_wire_280,dangling_wire_281,dangling_wire_282,\line_buffer.n525 ,dangling_wire_283,dangling_wire_284,dangling_wire_285}),
            .RADDR({N__16309,N__19105,N__19555,N__17233,N__17497,N__16960,N__9244,N__14119,N__18841,N__15799,N__16057}),
            .WADDR({N__12460,N__10561,N__10816,N__11065,N__11323,N__11587,N__11950,N__12208,N__13033,N__10057,N__10312}),
            .MASK({dangling_wire_286,dangling_wire_287,dangling_wire_288,dangling_wire_289,dangling_wire_290,dangling_wire_291,dangling_wire_292,dangling_wire_293,dangling_wire_294,dangling_wire_295,dangling_wire_296,dangling_wire_297,dangling_wire_298,dangling_wire_299,dangling_wire_300,dangling_wire_301}),
            .WDATA({dangling_wire_302,dangling_wire_303,dangling_wire_304,dangling_wire_305,N__17882,dangling_wire_306,dangling_wire_307,dangling_wire_308,dangling_wire_309,dangling_wire_310,dangling_wire_311,dangling_wire_312,N__19765,dangling_wire_313,dangling_wire_314,dangling_wire_315}),
            .RCLKE(),
            .RCLK(N__23542),
            .RE(N__18208),
            .WCLKE(),
            .WCLK(N__24589),
            .WE(N__8613));
    defparam \line_buffer.mem1_physical .WRITE_MODE=3;
    defparam \line_buffer.mem1_physical .READ_MODE=3;
    defparam \line_buffer.mem1_physical .INIT_F=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem1_physical .INIT_E=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem1_physical .INIT_D=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem1_physical .INIT_C=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem1_physical .INIT_B=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem1_physical .INIT_A=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem1_physical .INIT_9=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem1_physical .INIT_8=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem1_physical .INIT_7=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem1_physical .INIT_6=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem1_physical .INIT_5=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem1_physical .INIT_4=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem1_physical .INIT_3=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    defparam \line_buffer.mem1_physical .INIT_2=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    defparam \line_buffer.mem1_physical .INIT_1=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    defparam \line_buffer.mem1_physical .INIT_0=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    SB_RAM40_4K \line_buffer.mem1_physical  (
            .RDATA({dangling_wire_316,dangling_wire_317,dangling_wire_318,dangling_wire_319,\line_buffer.n554 ,dangling_wire_320,dangling_wire_321,dangling_wire_322,dangling_wire_323,dangling_wire_324,dangling_wire_325,dangling_wire_326,\line_buffer.n553 ,dangling_wire_327,dangling_wire_328,dangling_wire_329}),
            .RADDR({N__16318,N__19096,N__19552,N__17236,N__17506,N__16969,N__9253,N__14135,N__18844,N__15802,N__16054}),
            .WADDR({N__12476,N__10570,N__10813,N__11068,N__11326,N__11584,N__11963,N__12221,N__13024,N__10054,N__10315}),
            .MASK({dangling_wire_330,dangling_wire_331,dangling_wire_332,dangling_wire_333,dangling_wire_334,dangling_wire_335,dangling_wire_336,dangling_wire_337,dangling_wire_338,dangling_wire_339,dangling_wire_340,dangling_wire_341,dangling_wire_342,dangling_wire_343,dangling_wire_344,dangling_wire_345}),
            .WDATA({dangling_wire_346,dangling_wire_347,dangling_wire_348,dangling_wire_349,N__22132,dangling_wire_350,dangling_wire_351,dangling_wire_352,dangling_wire_353,dangling_wire_354,dangling_wire_355,dangling_wire_356,N__18540,dangling_wire_357,dangling_wire_358,dangling_wire_359}),
            .RCLKE(),
            .RCLK(N__23427),
            .RE(N__18213),
            .WCLKE(),
            .WCLK(N__24585),
            .WE(N__13400));
    defparam \line_buffer.mem15_physical .WRITE_MODE=3;
    defparam \line_buffer.mem15_physical .READ_MODE=3;
    defparam \line_buffer.mem15_physical .INIT_F=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem15_physical .INIT_E=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem15_physical .INIT_D=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem15_physical .INIT_C=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem15_physical .INIT_B=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem15_physical .INIT_A=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem15_physical .INIT_9=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem15_physical .INIT_8=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem15_physical .INIT_7=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem15_physical .INIT_6=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem15_physical .INIT_5=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem15_physical .INIT_4=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem15_physical .INIT_3=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    defparam \line_buffer.mem15_physical .INIT_2=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    defparam \line_buffer.mem15_physical .INIT_1=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    defparam \line_buffer.mem15_physical .INIT_0=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    SB_RAM40_4K \line_buffer.mem15_physical  (
            .RDATA({dangling_wire_360,dangling_wire_361,dangling_wire_362,dangling_wire_363,\line_buffer.n550 ,dangling_wire_364,dangling_wire_365,dangling_wire_366,dangling_wire_367,dangling_wire_368,dangling_wire_369,dangling_wire_370,\line_buffer.n549 ,dangling_wire_371,dangling_wire_372,dangling_wire_373}),
            .RADDR({N__16246,N__19024,N__19480,N__17164,N__17434,N__16897,N__9181,N__14068,N__18772,N__15730,N__15982}),
            .WADDR({N__12409,N__10498,N__10741,N__10996,N__11254,N__11512,N__11893,N__12151,N__12952,N__9982,N__10243}),
            .MASK({dangling_wire_374,dangling_wire_375,dangling_wire_376,dangling_wire_377,dangling_wire_378,dangling_wire_379,dangling_wire_380,dangling_wire_381,dangling_wire_382,dangling_wire_383,dangling_wire_384,dangling_wire_385,dangling_wire_386,dangling_wire_387,dangling_wire_388,dangling_wire_389}),
            .WDATA({dangling_wire_390,dangling_wire_391,dangling_wire_392,dangling_wire_393,N__17913,dangling_wire_394,dangling_wire_395,dangling_wire_396,dangling_wire_397,dangling_wire_398,dangling_wire_399,dangling_wire_400,N__19770,dangling_wire_401,dangling_wire_402,dangling_wire_403}),
            .RCLKE(),
            .RCLK(N__23426),
            .RE(N__18141),
            .WCLKE(),
            .WCLK(N__24613),
            .WE(N__13392));
    defparam \line_buffer.mem27_physical .WRITE_MODE=3;
    defparam \line_buffer.mem27_physical .READ_MODE=3;
    defparam \line_buffer.mem27_physical .INIT_F=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem27_physical .INIT_E=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem27_physical .INIT_D=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem27_physical .INIT_C=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem27_physical .INIT_B=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem27_physical .INIT_A=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem27_physical .INIT_9=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem27_physical .INIT_8=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem27_physical .INIT_7=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem27_physical .INIT_6=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem27_physical .INIT_5=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem27_physical .INIT_4=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem27_physical .INIT_3=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    defparam \line_buffer.mem27_physical .INIT_2=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    defparam \line_buffer.mem27_physical .INIT_1=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    defparam \line_buffer.mem27_physical .INIT_0=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    SB_RAM40_4K \line_buffer.mem27_physical  (
            .RDATA({dangling_wire_404,dangling_wire_405,dangling_wire_406,dangling_wire_407,\line_buffer.n558 ,dangling_wire_408,dangling_wire_409,dangling_wire_410,dangling_wire_411,dangling_wire_412,dangling_wire_413,dangling_wire_414,\line_buffer.n557 ,dangling_wire_415,dangling_wire_416,dangling_wire_417}),
            .RADDR({N__16273,N__19069,N__19519,N__17197,N__17461,N__16924,N__9208,N__14083,N__18805,N__15763,N__16021}),
            .WADDR({N__12424,N__10525,N__10780,N__11029,N__11287,N__11551,N__11914,N__12172,N__12997,N__10021,N__10276}),
            .MASK({dangling_wire_418,dangling_wire_419,dangling_wire_420,dangling_wire_421,dangling_wire_422,dangling_wire_423,dangling_wire_424,dangling_wire_425,dangling_wire_426,dangling_wire_427,dangling_wire_428,dangling_wire_429,dangling_wire_430,dangling_wire_431,dangling_wire_432,dangling_wire_433}),
            .WDATA({dangling_wire_434,dangling_wire_435,dangling_wire_436,dangling_wire_437,N__17912,dangling_wire_438,dangling_wire_439,dangling_wire_440,dangling_wire_441,dangling_wire_442,dangling_wire_443,dangling_wire_444,N__19748,dangling_wire_445,dangling_wire_446,dangling_wire_447}),
            .RCLKE(),
            .RCLK(N__23517),
            .RE(N__18185),
            .WCLKE(),
            .WCLK(N__24607),
            .WE(N__9618));
    defparam \line_buffer.mem4_physical .WRITE_MODE=3;
    defparam \line_buffer.mem4_physical .READ_MODE=3;
    defparam \line_buffer.mem4_physical .INIT_F=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem4_physical .INIT_E=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem4_physical .INIT_D=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem4_physical .INIT_C=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem4_physical .INIT_B=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem4_physical .INIT_A=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem4_physical .INIT_9=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem4_physical .INIT_8=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem4_physical .INIT_7=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem4_physical .INIT_6=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem4_physical .INIT_5=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem4_physical .INIT_4=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem4_physical .INIT_3=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem4_physical .INIT_2=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem4_physical .INIT_1=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem4_physical .INIT_0=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    SB_RAM40_4K \line_buffer.mem4_physical  (
            .RDATA({dangling_wire_448,dangling_wire_449,dangling_wire_450,dangling_wire_451,\line_buffer.n530 ,dangling_wire_452,dangling_wire_453,dangling_wire_454,dangling_wire_455,dangling_wire_456,dangling_wire_457,dangling_wire_458,\line_buffer.n529 ,dangling_wire_459,dangling_wire_460,dangling_wire_461}),
            .RADDR({N__16201,N__18997,N__19447,N__17125,N__17389,N__16852,N__9136,N__14011,N__18733,N__15691,N__15949}),
            .WADDR({N__12352,N__10453,N__10708,N__10957,N__11215,N__11479,N__11842,N__12100,N__12925,N__9949,N__10204}),
            .MASK({dangling_wire_462,dangling_wire_463,dangling_wire_464,dangling_wire_465,dangling_wire_466,dangling_wire_467,dangling_wire_468,dangling_wire_469,dangling_wire_470,dangling_wire_471,dangling_wire_472,dangling_wire_473,dangling_wire_474,dangling_wire_475,dangling_wire_476,dangling_wire_477}),
            .WDATA({dangling_wire_478,dangling_wire_479,dangling_wire_480,dangling_wire_481,N__22135,dangling_wire_482,dangling_wire_483,dangling_wire_484,dangling_wire_485,dangling_wire_486,dangling_wire_487,dangling_wire_488,N__18560,dangling_wire_489,dangling_wire_490,dangling_wire_491}),
            .RCLKE(),
            .RCLK(N__23318),
            .RE(N__18094),
            .WCLKE(),
            .WCLK(N__24622),
            .WE(N__8615));
    defparam \line_buffer.mem16_physical .WRITE_MODE=3;
    defparam \line_buffer.mem16_physical .READ_MODE=3;
    defparam \line_buffer.mem16_physical .INIT_F=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem16_physical .INIT_E=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem16_physical .INIT_D=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem16_physical .INIT_C=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem16_physical .INIT_B=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem16_physical .INIT_A=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem16_physical .INIT_9=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem16_physical .INIT_8=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem16_physical .INIT_7=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem16_physical .INIT_6=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem16_physical .INIT_5=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem16_physical .INIT_4=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem16_physical .INIT_3=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    defparam \line_buffer.mem16_physical .INIT_2=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    defparam \line_buffer.mem16_physical .INIT_1=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    defparam \line_buffer.mem16_physical .INIT_0=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    SB_RAM40_4K \line_buffer.mem16_physical  (
            .RDATA({dangling_wire_492,dangling_wire_493,dangling_wire_494,dangling_wire_495,\line_buffer.n548 ,dangling_wire_496,dangling_wire_497,dangling_wire_498,dangling_wire_499,dangling_wire_500,dangling_wire_501,dangling_wire_502,\line_buffer.n547 ,dangling_wire_503,dangling_wire_504,dangling_wire_505}),
            .RADDR({N__16234,N__19012,N__19468,N__17152,N__17422,N__16885,N__9169,N__14056,N__18760,N__15718,N__15970}),
            .WADDR({N__12397,N__10486,N__10729,N__10984,N__11242,N__11500,N__11881,N__12139,N__12940,N__9970,N__10231}),
            .MASK({dangling_wire_506,dangling_wire_507,dangling_wire_508,dangling_wire_509,dangling_wire_510,dangling_wire_511,dangling_wire_512,dangling_wire_513,dangling_wire_514,dangling_wire_515,dangling_wire_516,dangling_wire_517,dangling_wire_518,dangling_wire_519,dangling_wire_520,dangling_wire_521}),
            .WDATA({dangling_wire_522,dangling_wire_523,dangling_wire_524,dangling_wire_525,N__14334,dangling_wire_526,dangling_wire_527,dangling_wire_528,dangling_wire_529,dangling_wire_530,dangling_wire_531,dangling_wire_532,N__11716,dangling_wire_533,dangling_wire_534,dangling_wire_535}),
            .RCLKE(),
            .RCLK(N__23429),
            .RE(N__18140),
            .WCLKE(),
            .WCLK(N__24616),
            .WE(N__13399));
    defparam \line_buffer.mem30_physical .WRITE_MODE=3;
    defparam \line_buffer.mem30_physical .READ_MODE=3;
    defparam \line_buffer.mem30_physical .INIT_F=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem30_physical .INIT_E=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem30_physical .INIT_D=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem30_physical .INIT_C=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem30_physical .INIT_B=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem30_physical .INIT_A=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem30_physical .INIT_9=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem30_physical .INIT_8=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem30_physical .INIT_7=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem30_physical .INIT_6=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem30_physical .INIT_5=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem30_physical .INIT_4=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem30_physical .INIT_3=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    defparam \line_buffer.mem30_physical .INIT_2=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    defparam \line_buffer.mem30_physical .INIT_1=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    defparam \line_buffer.mem30_physical .INIT_0=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    SB_RAM40_4K \line_buffer.mem30_physical  (
            .RDATA({dangling_wire_536,dangling_wire_537,dangling_wire_538,dangling_wire_539,\line_buffer.n590 ,dangling_wire_540,dangling_wire_541,dangling_wire_542,dangling_wire_543,dangling_wire_544,dangling_wire_545,dangling_wire_546,\line_buffer.n589 ,dangling_wire_547,dangling_wire_548,dangling_wire_549}),
            .RADDR({N__16225,N__19021,N__19471,N__17149,N__17413,N__16876,N__9160,N__14035,N__18757,N__15715,N__15973}),
            .WADDR({N__12376,N__10477,N__10732,N__10981,N__11239,N__11503,N__11866,N__12124,N__12949,N__9973,N__10228}),
            .MASK({dangling_wire_550,dangling_wire_551,dangling_wire_552,dangling_wire_553,dangling_wire_554,dangling_wire_555,dangling_wire_556,dangling_wire_557,dangling_wire_558,dangling_wire_559,dangling_wire_560,dangling_wire_561,dangling_wire_562,dangling_wire_563,dangling_wire_564,dangling_wire_565}),
            .WDATA({dangling_wire_566,dangling_wire_567,dangling_wire_568,dangling_wire_569,N__17892,dangling_wire_570,dangling_wire_571,dangling_wire_572,dangling_wire_573,dangling_wire_574,dangling_wire_575,dangling_wire_576,N__19766,dangling_wire_577,dangling_wire_578,dangling_wire_579}),
            .RCLKE(),
            .RCLK(N__23440),
            .RE(N__18125),
            .WCLKE(),
            .WCLK(N__24617),
            .WE(N__13485));
    defparam \line_buffer.mem7_physical .WRITE_MODE=3;
    defparam \line_buffer.mem7_physical .READ_MODE=3;
    defparam \line_buffer.mem7_physical .INIT_F=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem7_physical .INIT_E=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem7_physical .INIT_D=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem7_physical .INIT_C=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem7_physical .INIT_B=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem7_physical .INIT_A=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem7_physical .INIT_9=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem7_physical .INIT_8=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem7_physical .INIT_7=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem7_physical .INIT_6=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem7_physical .INIT_5=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem7_physical .INIT_4=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem7_physical .INIT_3=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem7_physical .INIT_2=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem7_physical .INIT_1=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem7_physical .INIT_0=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    SB_RAM40_4K \line_buffer.mem7_physical  (
            .RDATA({dangling_wire_580,dangling_wire_581,dangling_wire_582,dangling_wire_583,\line_buffer.n457 ,dangling_wire_584,dangling_wire_585,dangling_wire_586,dangling_wire_587,dangling_wire_588,dangling_wire_589,dangling_wire_590,\line_buffer.n456 ,dangling_wire_591,dangling_wire_592,dangling_wire_593}),
            .RADDR({N__16165,N__18961,N__19411,N__17089,N__17353,N__16816,N__9100,N__13975,N__18697,N__15655,N__15913}),
            .WADDR({N__12316,N__10417,N__10672,N__10921,N__11179,N__11443,N__11806,N__12064,N__12889,N__9913,N__10168}),
            .MASK({dangling_wire_594,dangling_wire_595,dangling_wire_596,dangling_wire_597,dangling_wire_598,dangling_wire_599,dangling_wire_600,dangling_wire_601,dangling_wire_602,dangling_wire_603,dangling_wire_604,dangling_wire_605,dangling_wire_606,dangling_wire_607,dangling_wire_608,dangling_wire_609}),
            .WDATA({dangling_wire_610,dangling_wire_611,dangling_wire_612,dangling_wire_613,N__22150,dangling_wire_614,dangling_wire_615,dangling_wire_616,dangling_wire_617,dangling_wire_618,dangling_wire_619,dangling_wire_620,N__18569,dangling_wire_621,dangling_wire_622,dangling_wire_623}),
            .RCLKE(),
            .RCLK(N__23011),
            .RE(N__18052),
            .WCLKE(),
            .WCLK(N__24630),
            .WE(N__9375));
    defparam \line_buffer.mem20_physical .WRITE_MODE=3;
    defparam \line_buffer.mem20_physical .READ_MODE=3;
    defparam \line_buffer.mem20_physical .INIT_F=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem20_physical .INIT_E=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem20_physical .INIT_D=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem20_physical .INIT_C=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem20_physical .INIT_B=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem20_physical .INIT_A=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem20_physical .INIT_9=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem20_physical .INIT_8=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem20_physical .INIT_7=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem20_physical .INIT_6=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem20_physical .INIT_5=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem20_physical .INIT_4=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem20_physical .INIT_3=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem20_physical .INIT_2=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem20_physical .INIT_1=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem20_physical .INIT_0=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    SB_RAM40_4K \line_buffer.mem20_physical  (
            .RDATA({dangling_wire_624,dangling_wire_625,dangling_wire_626,dangling_wire_627,\line_buffer.n584 ,dangling_wire_628,dangling_wire_629,dangling_wire_630,dangling_wire_631,dangling_wire_632,dangling_wire_633,dangling_wire_634,\line_buffer.n583 ,dangling_wire_635,dangling_wire_636,dangling_wire_637}),
            .RADDR({N__16174,N__18952,N__19408,N__17092,N__17362,N__16825,N__9109,N__13996,N__18700,N__15658,N__15910}),
            .WADDR({N__12337,N__10426,N__10669,N__10924,N__11182,N__11440,N__11821,N__12079,N__12880,N__9910,N__10171}),
            .MASK({dangling_wire_638,dangling_wire_639,dangling_wire_640,dangling_wire_641,dangling_wire_642,dangling_wire_643,dangling_wire_644,dangling_wire_645,dangling_wire_646,dangling_wire_647,dangling_wire_648,dangling_wire_649,dangling_wire_650,dangling_wire_651,dangling_wire_652,dangling_wire_653}),
            .WDATA({dangling_wire_654,dangling_wire_655,dangling_wire_656,dangling_wire_657,N__17672,dangling_wire_658,dangling_wire_659,dangling_wire_660,dangling_wire_661,dangling_wire_662,dangling_wire_663,dangling_wire_664,N__17788,dangling_wire_665,dangling_wire_666,dangling_wire_667}),
            .RCLKE(),
            .RCLK(N__23091),
            .RE(N__18088),
            .WCLKE(),
            .WCLK(N__24629),
            .WE(N__12690));
    defparam \line_buffer.mem13_physical .WRITE_MODE=3;
    defparam \line_buffer.mem13_physical .READ_MODE=3;
    defparam \line_buffer.mem13_physical .INIT_F=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem13_physical .INIT_E=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem13_physical .INIT_D=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem13_physical .INIT_C=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem13_physical .INIT_B=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem13_physical .INIT_A=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem13_physical .INIT_9=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem13_physical .INIT_8=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem13_physical .INIT_7=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem13_physical .INIT_6=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem13_physical .INIT_5=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem13_physical .INIT_4=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem13_physical .INIT_3=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem13_physical .INIT_2=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem13_physical .INIT_1=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem13_physical .INIT_0=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    SB_RAM40_4K \line_buffer.mem13_physical  (
            .RDATA({dangling_wire_668,dangling_wire_669,dangling_wire_670,dangling_wire_671,\line_buffer.n516 ,dangling_wire_672,dangling_wire_673,dangling_wire_674,dangling_wire_675,dangling_wire_676,dangling_wire_677,dangling_wire_678,\line_buffer.n515 ,dangling_wire_679,dangling_wire_680,dangling_wire_681}),
            .RADDR({N__16270,N__19048,N__19504,N__17188,N__17458,N__16921,N__9205,N__14092,N__18796,N__15754,N__16006}),
            .WADDR({N__12433,N__10522,N__10765,N__11020,N__11278,N__11536,N__11917,N__12175,N__12976,N__10006,N__10267}),
            .MASK({dangling_wire_682,dangling_wire_683,dangling_wire_684,dangling_wire_685,dangling_wire_686,dangling_wire_687,dangling_wire_688,dangling_wire_689,dangling_wire_690,dangling_wire_691,dangling_wire_692,dangling_wire_693,dangling_wire_694,dangling_wire_695,dangling_wire_696,dangling_wire_697}),
            .WDATA({dangling_wire_698,dangling_wire_699,dangling_wire_700,dangling_wire_701,N__14327,dangling_wire_702,dangling_wire_703,dangling_wire_704,dangling_wire_705,dangling_wire_706,dangling_wire_707,dangling_wire_708,N__11699,dangling_wire_709,dangling_wire_710,dangling_wire_711}),
            .RCLKE(),
            .RCLK(N__22997),
            .RE(N__18171),
            .WCLKE(),
            .WCLK(N__24608),
            .WE(N__14394));
    defparam \line_buffer.mem19_physical .WRITE_MODE=3;
    defparam \line_buffer.mem19_physical .READ_MODE=3;
    defparam \line_buffer.mem19_physical .INIT_F=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem19_physical .INIT_E=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem19_physical .INIT_D=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem19_physical .INIT_C=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem19_physical .INIT_B=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem19_physical .INIT_A=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem19_physical .INIT_9=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem19_physical .INIT_8=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem19_physical .INIT_7=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem19_physical .INIT_6=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem19_physical .INIT_5=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem19_physical .INIT_4=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem19_physical .INIT_3=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem19_physical .INIT_2=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem19_physical .INIT_1=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem19_physical .INIT_0=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    SB_RAM40_4K \line_buffer.mem19_physical  (
            .RDATA({dangling_wire_712,dangling_wire_713,dangling_wire_714,dangling_wire_715,\line_buffer.n459 ,dangling_wire_716,dangling_wire_717,dangling_wire_718,dangling_wire_719,dangling_wire_720,dangling_wire_721,dangling_wire_722,\line_buffer.n458 ,dangling_wire_723,dangling_wire_724,dangling_wire_725}),
            .RADDR({N__16198,N__18976,N__19432,N__17116,N__17386,N__16849,N__9133,N__14020,N__18724,N__15682,N__15934}),
            .WADDR({N__12361,N__10450,N__10693,N__10948,N__11206,N__11464,N__11845,N__12103,N__12904,N__9934,N__10195}),
            .MASK({dangling_wire_726,dangling_wire_727,dangling_wire_728,dangling_wire_729,dangling_wire_730,dangling_wire_731,dangling_wire_732,dangling_wire_733,dangling_wire_734,dangling_wire_735,dangling_wire_736,dangling_wire_737,dangling_wire_738,dangling_wire_739,dangling_wire_740,dangling_wire_741}),
            .WDATA({dangling_wire_742,dangling_wire_743,dangling_wire_744,dangling_wire_745,N__14335,dangling_wire_746,dangling_wire_747,dangling_wire_748,dangling_wire_749,dangling_wire_750,dangling_wire_751,dangling_wire_752,N__11717,dangling_wire_753,dangling_wire_754,dangling_wire_755}),
            .RCLKE(),
            .RCLK(N__23124),
            .RE(N__18073),
            .WCLKE(),
            .WCLK(N__24623),
            .WE(N__14182));
    defparam \line_buffer.mem23_physical .WRITE_MODE=3;
    defparam \line_buffer.mem23_physical .READ_MODE=3;
    defparam \line_buffer.mem23_physical .INIT_F=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem23_physical .INIT_E=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem23_physical .INIT_D=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem23_physical .INIT_C=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem23_physical .INIT_B=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem23_physical .INIT_A=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem23_physical .INIT_9=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem23_physical .INIT_8=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem23_physical .INIT_7=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem23_physical .INIT_6=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem23_physical .INIT_5=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem23_physical .INIT_4=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem23_physical .INIT_3=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem23_physical .INIT_2=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem23_physical .INIT_1=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem23_physical .INIT_0=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    SB_RAM40_4K \line_buffer.mem23_physical  (
            .RDATA({dangling_wire_756,dangling_wire_757,dangling_wire_758,dangling_wire_759,\line_buffer.n528 ,dangling_wire_760,dangling_wire_761,dangling_wire_762,dangling_wire_763,dangling_wire_764,dangling_wire_765,dangling_wire_766,\line_buffer.n527 ,dangling_wire_767,dangling_wire_768,dangling_wire_769}),
            .RADDR({N__16321,N__19112,N__19565,N__17245,N__17509,N__16972,N__9256,N__14131,N__18853,N__15811,N__16067}),
            .WADDR({N__12472,N__10573,N__10826,N__11077,N__11335,N__11597,N__11962,N__12220,N__13040,N__10067,N__10324}),
            .MASK({dangling_wire_770,dangling_wire_771,dangling_wire_772,dangling_wire_773,dangling_wire_774,dangling_wire_775,dangling_wire_776,dangling_wire_777,dangling_wire_778,dangling_wire_779,dangling_wire_780,dangling_wire_781,dangling_wire_782,dangling_wire_783,dangling_wire_784,dangling_wire_785}),
            .WDATA({dangling_wire_786,dangling_wire_787,dangling_wire_788,dangling_wire_789,N__17677,dangling_wire_790,dangling_wire_791,dangling_wire_792,dangling_wire_793,dangling_wire_794,dangling_wire_795,dangling_wire_796,N__17770,dangling_wire_797,dangling_wire_798,dangling_wire_799}),
            .RCLKE(),
            .RCLK(N__23546),
            .RE(N__18217),
            .WCLKE(),
            .WCLK(N__24579),
            .WE(N__8614));
    defparam \line_buffer.mem0_physical .WRITE_MODE=3;
    defparam \line_buffer.mem0_physical .READ_MODE=3;
    defparam \line_buffer.mem0_physical .INIT_F=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem0_physical .INIT_E=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem0_physical .INIT_D=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem0_physical .INIT_C=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem0_physical .INIT_B=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem0_physical .INIT_A=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem0_physical .INIT_9=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem0_physical .INIT_8=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem0_physical .INIT_7=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem0_physical .INIT_6=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem0_physical .INIT_5=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem0_physical .INIT_4=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem0_physical .INIT_3=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem0_physical .INIT_2=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem0_physical .INIT_1=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem0_physical .INIT_0=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    SB_RAM40_4K \line_buffer.mem0_physical  (
            .RDATA({dangling_wire_800,dangling_wire_801,dangling_wire_802,dangling_wire_803,\line_buffer.n522 ,dangling_wire_804,dangling_wire_805,dangling_wire_806,dangling_wire_807,dangling_wire_808,dangling_wire_809,dangling_wire_810,\line_buffer.n521 ,dangling_wire_811,dangling_wire_812,dangling_wire_813}),
            .RADDR({N__16325,N__19108,N__19564,N__17246,N__17513,N__16976,N__9260,N__14141,N__18854,N__15812,N__16066}),
            .WADDR({N__12482,N__10577,N__10825,N__11078,N__11336,N__11596,N__11969,N__12227,N__13036,N__10066,N__10325}),
            .MASK({dangling_wire_814,dangling_wire_815,dangling_wire_816,dangling_wire_817,dangling_wire_818,dangling_wire_819,dangling_wire_820,dangling_wire_821,dangling_wire_822,dangling_wire_823,dangling_wire_824,dangling_wire_825,dangling_wire_826,dangling_wire_827,dangling_wire_828,dangling_wire_829}),
            .WDATA({dangling_wire_830,dangling_wire_831,dangling_wire_832,dangling_wire_833,N__22133,dangling_wire_834,dangling_wire_835,dangling_wire_836,dangling_wire_837,dangling_wire_838,dangling_wire_839,dangling_wire_840,N__18558,dangling_wire_841,dangling_wire_842,dangling_wire_843}),
            .RCLKE(),
            .RCLK(N__23428),
            .RE(N__18218),
            .WCLKE(),
            .WCLK(N__24574),
            .WE(N__14399));
    defparam \line_buffer.mem26_physical .WRITE_MODE=3;
    defparam \line_buffer.mem26_physical .READ_MODE=3;
    defparam \line_buffer.mem26_physical .INIT_F=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem26_physical .INIT_E=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem26_physical .INIT_D=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem26_physical .INIT_C=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem26_physical .INIT_B=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem26_physical .INIT_A=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem26_physical .INIT_9=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem26_physical .INIT_8=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem26_physical .INIT_7=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem26_physical .INIT_6=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem26_physical .INIT_5=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem26_physical .INIT_4=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem26_physical .INIT_3=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    defparam \line_buffer.mem26_physical .INIT_2=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    defparam \line_buffer.mem26_physical .INIT_1=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    defparam \line_buffer.mem26_physical .INIT_0=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    SB_RAM40_4K \line_buffer.mem26_physical  (
            .RDATA({dangling_wire_844,dangling_wire_845,dangling_wire_846,dangling_wire_847,\line_buffer.n560 ,dangling_wire_848,dangling_wire_849,dangling_wire_850,dangling_wire_851,dangling_wire_852,dangling_wire_853,dangling_wire_854,\line_buffer.n559 ,dangling_wire_855,dangling_wire_856,dangling_wire_857}),
            .RADDR({N__16285,N__19081,N__19531,N__17209,N__17473,N__16936,N__9220,N__14095,N__18817,N__15775,N__16033}),
            .WADDR({N__12436,N__10537,N__10792,N__11041,N__11299,N__11563,N__11926,N__12184,N__13009,N__10033,N__10288}),
            .MASK({dangling_wire_858,dangling_wire_859,dangling_wire_860,dangling_wire_861,dangling_wire_862,dangling_wire_863,dangling_wire_864,dangling_wire_865,dangling_wire_866,dangling_wire_867,dangling_wire_868,dangling_wire_869,dangling_wire_870,dangling_wire_871,dangling_wire_872,dangling_wire_873}),
            .WDATA({dangling_wire_874,dangling_wire_875,dangling_wire_876,dangling_wire_877,N__17645,dangling_wire_878,dangling_wire_879,dangling_wire_880,dangling_wire_881,dangling_wire_882,dangling_wire_883,dangling_wire_884,N__17774,dangling_wire_885,dangling_wire_886,dangling_wire_887}),
            .RCLKE(),
            .RCLK(N__23526),
            .RE(N__18186),
            .WCLKE(),
            .WCLK(N__24603),
            .WE(N__9640));
    defparam \line_buffer.mem3_physical .WRITE_MODE=3;
    defparam \line_buffer.mem3_physical .READ_MODE=3;
    defparam \line_buffer.mem3_physical .INIT_F=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem3_physical .INIT_E=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem3_physical .INIT_D=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem3_physical .INIT_C=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem3_physical .INIT_B=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem3_physical .INIT_A=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem3_physical .INIT_9=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem3_physical .INIT_8=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem3_physical .INIT_7=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem3_physical .INIT_6=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem3_physical .INIT_5=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem3_physical .INIT_4=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem3_physical .INIT_3=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem3_physical .INIT_2=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem3_physical .INIT_1=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem3_physical .INIT_0=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    SB_RAM40_4K \line_buffer.mem3_physical  (
            .RDATA({dangling_wire_888,dangling_wire_889,dangling_wire_890,dangling_wire_891,\line_buffer.n586 ,dangling_wire_892,dangling_wire_893,dangling_wire_894,dangling_wire_895,dangling_wire_896,dangling_wire_897,dangling_wire_898,\line_buffer.n585 ,dangling_wire_899,dangling_wire_900,dangling_wire_901}),
            .RADDR({N__16237,N__19033,N__19483,N__17161,N__17425,N__16888,N__9172,N__14047,N__18769,N__15727,N__15985}),
            .WADDR({N__12388,N__10489,N__10744,N__10993,N__11251,N__11515,N__11878,N__12136,N__12961,N__9985,N__10240}),
            .MASK({dangling_wire_902,dangling_wire_903,dangling_wire_904,dangling_wire_905,dangling_wire_906,dangling_wire_907,dangling_wire_908,dangling_wire_909,dangling_wire_910,dangling_wire_911,dangling_wire_912,dangling_wire_913,dangling_wire_914,dangling_wire_915,dangling_wire_916,dangling_wire_917}),
            .WDATA({dangling_wire_918,dangling_wire_919,dangling_wire_920,dangling_wire_921,N__22134,dangling_wire_922,dangling_wire_923,dangling_wire_924,dangling_wire_925,dangling_wire_926,dangling_wire_927,dangling_wire_928,N__18532,dangling_wire_929,dangling_wire_930,dangling_wire_931}),
            .RCLKE(),
            .RCLK(N__23304),
            .RE(N__18126),
            .WCLKE(),
            .WCLK(N__24615),
            .WE(N__12680));
    defparam \line_buffer.mem17_physical .WRITE_MODE=3;
    defparam \line_buffer.mem17_physical .READ_MODE=3;
    defparam \line_buffer.mem17_physical .INIT_F=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem17_physical .INIT_E=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem17_physical .INIT_D=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem17_physical .INIT_C=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem17_physical .INIT_B=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem17_physical .INIT_A=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem17_physical .INIT_9=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem17_physical .INIT_8=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem17_physical .INIT_7=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem17_physical .INIT_6=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem17_physical .INIT_5=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem17_physical .INIT_4=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem17_physical .INIT_3=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem17_physical .INIT_2=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem17_physical .INIT_1=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem17_physical .INIT_0=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    SB_RAM40_4K \line_buffer.mem17_physical  (
            .RDATA({dangling_wire_932,dangling_wire_933,dangling_wire_934,dangling_wire_935,\line_buffer.n463 ,dangling_wire_936,dangling_wire_937,dangling_wire_938,dangling_wire_939,dangling_wire_940,dangling_wire_941,dangling_wire_942,\line_buffer.n462 ,dangling_wire_943,dangling_wire_944,dangling_wire_945}),
            .RADDR({N__16222,N__19000,N__19456,N__17140,N__17410,N__16873,N__9157,N__14044,N__18748,N__15706,N__15958}),
            .WADDR({N__12385,N__10474,N__10717,N__10972,N__11230,N__11488,N__11869,N__12127,N__12928,N__9958,N__10219}),
            .MASK({dangling_wire_946,dangling_wire_947,dangling_wire_948,dangling_wire_949,dangling_wire_950,dangling_wire_951,dangling_wire_952,dangling_wire_953,dangling_wire_954,dangling_wire_955,dangling_wire_956,dangling_wire_957,dangling_wire_958,dangling_wire_959,dangling_wire_960,dangling_wire_961}),
            .WDATA({dangling_wire_962,dangling_wire_963,dangling_wire_964,dangling_wire_965,N__17658,dangling_wire_966,dangling_wire_967,dangling_wire_968,dangling_wire_969,dangling_wire_970,dangling_wire_971,dangling_wire_972,N__17775,dangling_wire_973,dangling_wire_974,dangling_wire_975}),
            .RCLKE(),
            .RCLK(N__23312),
            .RE(N__18110),
            .WCLKE(),
            .WCLK(N__24618),
            .WE(N__14174));
    defparam \line_buffer.mem31_physical .WRITE_MODE=3;
    defparam \line_buffer.mem31_physical .READ_MODE=3;
    defparam \line_buffer.mem31_physical .INIT_F=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem31_physical .INIT_E=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem31_physical .INIT_D=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem31_physical .INIT_C=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem31_physical .INIT_B=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem31_physical .INIT_A=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem31_physical .INIT_9=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem31_physical .INIT_8=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem31_physical .INIT_7=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem31_physical .INIT_6=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem31_physical .INIT_5=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem31_physical .INIT_4=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem31_physical .INIT_3=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    defparam \line_buffer.mem31_physical .INIT_2=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    defparam \line_buffer.mem31_physical .INIT_1=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    defparam \line_buffer.mem31_physical .INIT_0=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    SB_RAM40_4K \line_buffer.mem31_physical  (
            .RDATA({dangling_wire_976,dangling_wire_977,dangling_wire_978,dangling_wire_979,\line_buffer.n588 ,dangling_wire_980,dangling_wire_981,dangling_wire_982,dangling_wire_983,dangling_wire_984,dangling_wire_985,dangling_wire_986,\line_buffer.n587 ,dangling_wire_987,dangling_wire_988,dangling_wire_989}),
            .RADDR({N__16213,N__19009,N__19459,N__17137,N__17401,N__16864,N__9148,N__14023,N__18745,N__15703,N__15961}),
            .WADDR({N__12364,N__10465,N__10720,N__10969,N__11227,N__11491,N__11854,N__12112,N__12937,N__9961,N__10216}),
            .MASK({dangling_wire_990,dangling_wire_991,dangling_wire_992,dangling_wire_993,dangling_wire_994,dangling_wire_995,dangling_wire_996,dangling_wire_997,dangling_wire_998,dangling_wire_999,dangling_wire_1000,dangling_wire_1001,dangling_wire_1002,dangling_wire_1003,dangling_wire_1004,dangling_wire_1005}),
            .WDATA({dangling_wire_1006,dangling_wire_1007,dangling_wire_1008,dangling_wire_1009,N__14348,dangling_wire_1010,dangling_wire_1011,dangling_wire_1012,dangling_wire_1013,dangling_wire_1014,dangling_wire_1015,dangling_wire_1016,N__11721,dangling_wire_1017,dangling_wire_1018,dangling_wire_1019}),
            .RCLKE(),
            .RCLK(N__23165),
            .RE(N__18095),
            .WCLKE(),
            .WCLK(N__24620),
            .WE(N__13486));
    defparam \line_buffer.mem9_physical .INIT_0=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem9_physical .WRITE_MODE=3;
    defparam \line_buffer.mem9_physical .READ_MODE=3;
    defparam \line_buffer.mem9_physical .INIT_F=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem9_physical .INIT_E=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem9_physical .INIT_D=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem9_physical .INIT_C=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem9_physical .INIT_B=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem9_physical .INIT_A=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem9_physical .INIT_9=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem9_physical .INIT_8=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem9_physical .INIT_7=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem9_physical .INIT_6=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem9_physical .INIT_5=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem9_physical .INIT_4=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem9_physical .INIT_3=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem9_physical .INIT_2=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem9_physical .INIT_1=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    SB_RAM40_4K \line_buffer.mem9_physical  (
            .RDATA({dangling_wire_1020,dangling_wire_1021,dangling_wire_1022,dangling_wire_1023,\line_buffer.n453 ,dangling_wire_1024,dangling_wire_1025,dangling_wire_1026,dangling_wire_1027,dangling_wire_1028,dangling_wire_1029,dangling_wire_1030,\line_buffer.n452 ,dangling_wire_1031,dangling_wire_1032,dangling_wire_1033}),
            .RADDR({N__16141,N__18937,N__19387,N__17065,N__17329,N__16792,N__9076,N__13951,N__18673,N__15631,N__15889}),
            .WADDR({N__12291,N__10393,N__10648,N__10897,N__11155,N__11419,N__11781,N__12039,N__12865,N__9889,N__10144}),
            .MASK({dangling_wire_1034,dangling_wire_1035,dangling_wire_1036,dangling_wire_1037,dangling_wire_1038,dangling_wire_1039,dangling_wire_1040,dangling_wire_1041,dangling_wire_1042,dangling_wire_1043,dangling_wire_1044,dangling_wire_1045,dangling_wire_1046,dangling_wire_1047,dangling_wire_1048,dangling_wire_1049}),
            .WDATA({dangling_wire_1050,dangling_wire_1051,dangling_wire_1052,dangling_wire_1053,N__17924,dangling_wire_1054,dangling_wire_1055,dangling_wire_1056,dangling_wire_1057,dangling_wire_1058,dangling_wire_1059,dangling_wire_1060,N__19778,dangling_wire_1061,dangling_wire_1062,dangling_wire_1063}),
            .RCLKE(),
            .RCLK(N__22644),
            .RE(N__18093),
            .WCLKE(),
            .WCLK(N__24637),
            .WE(N__9383));
    defparam \line_buffer.mem29_physical .WRITE_MODE=3;
    defparam \line_buffer.mem29_physical .READ_MODE=3;
    defparam \line_buffer.mem29_physical .INIT_F=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem29_physical .INIT_E=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem29_physical .INIT_D=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem29_physical .INIT_C=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem29_physical .INIT_B=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem29_physical .INIT_A=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem29_physical .INIT_9=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem29_physical .INIT_8=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem29_physical .INIT_7=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem29_physical .INIT_6=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem29_physical .INIT_5=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem29_physical .INIT_4=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem29_physical .INIT_3=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    defparam \line_buffer.mem29_physical .INIT_2=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    defparam \line_buffer.mem29_physical .INIT_1=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    defparam \line_buffer.mem29_physical .INIT_0=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    SB_RAM40_4K \line_buffer.mem29_physical  (
            .RDATA({dangling_wire_1064,dangling_wire_1065,dangling_wire_1066,dangling_wire_1067,\line_buffer.n592 ,dangling_wire_1068,dangling_wire_1069,dangling_wire_1070,dangling_wire_1071,dangling_wire_1072,dangling_wire_1073,dangling_wire_1074,\line_buffer.n591 ,dangling_wire_1075,dangling_wire_1076,dangling_wire_1077}),
            .RADDR({N__16249,N__19045,N__19495,N__17173,N__17437,N__16900,N__9184,N__14059,N__18781,N__15739,N__15997}),
            .WADDR({N__12400,N__10501,N__10756,N__11005,N__11263,N__11527,N__11890,N__12148,N__12973,N__9997,N__10252}),
            .MASK({dangling_wire_1078,dangling_wire_1079,dangling_wire_1080,dangling_wire_1081,dangling_wire_1082,dangling_wire_1083,dangling_wire_1084,dangling_wire_1085,dangling_wire_1086,dangling_wire_1087,dangling_wire_1088,dangling_wire_1089,dangling_wire_1090,dangling_wire_1091,dangling_wire_1092,dangling_wire_1093}),
            .WDATA({dangling_wire_1094,dangling_wire_1095,dangling_wire_1096,dangling_wire_1097,N__17673,dangling_wire_1098,dangling_wire_1099,dangling_wire_1100,dangling_wire_1101,dangling_wire_1102,dangling_wire_1103,dangling_wire_1104,N__17769,dangling_wire_1105,dangling_wire_1106,dangling_wire_1107}),
            .RCLKE(),
            .RCLK(N__23456),
            .RE(N__18155),
            .WCLKE(),
            .WCLK(N__24612),
            .WE(N__13484));
    defparam \line_buffer.mem6_physical .WRITE_MODE=3;
    defparam \line_buffer.mem6_physical .READ_MODE=3;
    defparam \line_buffer.mem6_physical .INIT_F=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem6_physical .INIT_E=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem6_physical .INIT_D=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem6_physical .INIT_C=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem6_physical .INIT_B=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem6_physical .INIT_A=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem6_physical .INIT_9=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem6_physical .INIT_8=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem6_physical .INIT_7=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem6_physical .INIT_6=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem6_physical .INIT_5=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem6_physical .INIT_4=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem6_physical .INIT_3=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    defparam \line_buffer.mem6_physical .INIT_2=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    defparam \line_buffer.mem6_physical .INIT_1=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    defparam \line_buffer.mem6_physical .INIT_0=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    SB_RAM40_4K \line_buffer.mem6_physical  (
            .RDATA({dangling_wire_1108,dangling_wire_1109,dangling_wire_1110,dangling_wire_1111,\line_buffer.n594 ,dangling_wire_1112,dangling_wire_1113,dangling_wire_1114,dangling_wire_1115,dangling_wire_1116,dangling_wire_1117,dangling_wire_1118,\line_buffer.n593 ,dangling_wire_1119,dangling_wire_1120,dangling_wire_1121}),
            .RADDR({N__16177,N__18973,N__19423,N__17101,N__17365,N__16828,N__9112,N__13987,N__18709,N__15667,N__15925}),
            .WADDR({N__12328,N__10429,N__10684,N__10933,N__11191,N__11455,N__11818,N__12076,N__12901,N__9925,N__10180}),
            .MASK({dangling_wire_1122,dangling_wire_1123,dangling_wire_1124,dangling_wire_1125,dangling_wire_1126,dangling_wire_1127,dangling_wire_1128,dangling_wire_1129,dangling_wire_1130,dangling_wire_1131,dangling_wire_1132,dangling_wire_1133,dangling_wire_1134,dangling_wire_1135,dangling_wire_1136,dangling_wire_1137}),
            .WDATA({dangling_wire_1138,dangling_wire_1139,dangling_wire_1140,dangling_wire_1141,N__22149,dangling_wire_1142,dangling_wire_1143,dangling_wire_1144,dangling_wire_1145,dangling_wire_1146,dangling_wire_1147,dangling_wire_1148,N__18568,dangling_wire_1149,dangling_wire_1150,dangling_wire_1151}),
            .RCLKE(),
            .RCLK(N__23182),
            .RE(N__18050),
            .WCLKE(),
            .WCLK(N__24627),
            .WE(N__13493));
    defparam \line_buffer.mem10_physical .WRITE_MODE=3;
    defparam \line_buffer.mem10_physical .READ_MODE=3;
    defparam \line_buffer.mem10_physical .INIT_F=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem10_physical .INIT_E=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem10_physical .INIT_D=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem10_physical .INIT_C=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem10_physical .INIT_B=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem10_physical .INIT_A=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem10_physical .INIT_9=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem10_physical .INIT_8=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem10_physical .INIT_7=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem10_physical .INIT_6=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem10_physical .INIT_5=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem10_physical .INIT_4=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem10_physical .INIT_3=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem10_physical .INIT_2=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem10_physical .INIT_1=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem10_physical .INIT_0=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    SB_RAM40_4K \line_buffer.mem10_physical  (
            .RDATA({dangling_wire_1152,dangling_wire_1153,dangling_wire_1154,dangling_wire_1155,\line_buffer.n451 ,dangling_wire_1156,dangling_wire_1157,dangling_wire_1158,dangling_wire_1159,dangling_wire_1160,dangling_wire_1161,dangling_wire_1162,\line_buffer.n450 ,dangling_wire_1163,dangling_wire_1164,dangling_wire_1165}),
            .RADDR({N__16306,N__19084,N__19540,N__17224,N__17494,N__16957,N__9241,N__14128,N__18832,N__15790,N__16042}),
            .WADDR({N__12469,N__10558,N__10801,N__11056,N__11314,N__11572,N__11953,N__12211,N__13012,N__10042,N__10303}),
            .MASK({dangling_wire_1166,dangling_wire_1167,dangling_wire_1168,dangling_wire_1169,dangling_wire_1170,dangling_wire_1171,dangling_wire_1172,dangling_wire_1173,dangling_wire_1174,dangling_wire_1175,dangling_wire_1176,dangling_wire_1177,dangling_wire_1178,dangling_wire_1179,dangling_wire_1180,dangling_wire_1181}),
            .WDATA({dangling_wire_1182,dangling_wire_1183,dangling_wire_1184,dangling_wire_1185,N__14339,dangling_wire_1186,dangling_wire_1187,dangling_wire_1188,dangling_wire_1189,dangling_wire_1190,dangling_wire_1191,dangling_wire_1192,N__11698,dangling_wire_1193,dangling_wire_1194,dangling_wire_1195}),
            .RCLKE(),
            .RCLK(N__23321),
            .RE(N__18212),
            .WCLKE(),
            .WCLK(N__24593),
            .WE(N__9361));
    defparam \line_buffer.mem22_physical .INIT_0=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem22_physical .WRITE_MODE=3;
    defparam \line_buffer.mem22_physical .READ_MODE=3;
    defparam \line_buffer.mem22_physical .INIT_F=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem22_physical .INIT_E=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem22_physical .INIT_D=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem22_physical .INIT_C=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem22_physical .INIT_B=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem22_physical .INIT_A=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem22_physical .INIT_9=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem22_physical .INIT_8=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem22_physical .INIT_7=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem22_physical .INIT_6=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem22_physical .INIT_5=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem22_physical .INIT_4=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem22_physical .INIT_3=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem22_physical .INIT_2=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem22_physical .INIT_1=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    SB_RAM40_4K \line_buffer.mem22_physical  (
            .RDATA({dangling_wire_1196,dangling_wire_1197,dangling_wire_1198,dangling_wire_1199,\line_buffer.n580 ,dangling_wire_1200,dangling_wire_1201,dangling_wire_1202,dangling_wire_1203,dangling_wire_1204,dangling_wire_1205,dangling_wire_1206,\line_buffer.n579 ,dangling_wire_1207,dangling_wire_1208,dangling_wire_1209}),
            .RADDR({N__16150,N__18928,N__19384,N__17068,N__17338,N__16801,N__9085,N__13972,N__18676,N__15634,N__15886}),
            .WADDR({N__12313,N__10402,N__10645,N__10900,N__11158,N__11416,N__11797,N__12055,N__12856,N__9886,N__10147}),
            .MASK({dangling_wire_1210,dangling_wire_1211,dangling_wire_1212,dangling_wire_1213,dangling_wire_1214,dangling_wire_1215,dangling_wire_1216,dangling_wire_1217,dangling_wire_1218,dangling_wire_1219,dangling_wire_1220,dangling_wire_1221,dangling_wire_1222,dangling_wire_1223,dangling_wire_1224,dangling_wire_1225}),
            .WDATA({dangling_wire_1226,dangling_wire_1227,dangling_wire_1228,dangling_wire_1229,N__14346,dangling_wire_1230,dangling_wire_1231,dangling_wire_1232,dangling_wire_1233,dangling_wire_1234,dangling_wire_1235,dangling_wire_1236,N__11723,dangling_wire_1237,dangling_wire_1238,dangling_wire_1239}),
            .RCLKE(),
            .RCLK(N__22751),
            .RE(N__18124),
            .WCLKE(),
            .WCLK(N__24636),
            .WE(N__12695));
    defparam \line_buffer.mem25_physical .WRITE_MODE=3;
    defparam \line_buffer.mem25_physical .READ_MODE=3;
    defparam \line_buffer.mem25_physical .INIT_F=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem25_physical .INIT_E=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem25_physical .INIT_D=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem25_physical .INIT_C=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem25_physical .INIT_B=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem25_physical .INIT_A=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem25_physical .INIT_9=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem25_physical .INIT_8=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem25_physical .INIT_7=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem25_physical .INIT_6=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem25_physical .INIT_5=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem25_physical .INIT_4=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem25_physical .INIT_3=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem25_physical .INIT_2=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem25_physical .INIT_1=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem25_physical .INIT_0=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    SB_RAM40_4K \line_buffer.mem25_physical  (
            .RDATA({dangling_wire_1240,dangling_wire_1241,dangling_wire_1242,dangling_wire_1243,\line_buffer.n524 ,dangling_wire_1244,dangling_wire_1245,dangling_wire_1246,dangling_wire_1247,dangling_wire_1248,dangling_wire_1249,dangling_wire_1250,\line_buffer.n523 ,dangling_wire_1251,dangling_wire_1252,dangling_wire_1253}),
            .RADDR({N__16297,N__19093,N__19543,N__17221,N__17485,N__16948,N__9232,N__14107,N__18829,N__15787,N__16045}),
            .WADDR({N__12448,N__10549,N__10804,N__11053,N__11311,N__11575,N__11938,N__12196,N__13021,N__10045,N__10300}),
            .MASK({dangling_wire_1254,dangling_wire_1255,dangling_wire_1256,dangling_wire_1257,dangling_wire_1258,dangling_wire_1259,dangling_wire_1260,dangling_wire_1261,dangling_wire_1262,dangling_wire_1263,dangling_wire_1264,dangling_wire_1265,dangling_wire_1266,dangling_wire_1267,dangling_wire_1268,dangling_wire_1269}),
            .WDATA({dangling_wire_1270,dangling_wire_1271,dangling_wire_1272,dangling_wire_1273,N__14347,dangling_wire_1274,dangling_wire_1275,dangling_wire_1276,dangling_wire_1277,dangling_wire_1278,dangling_wire_1279,dangling_wire_1280,N__11712,dangling_wire_1281,dangling_wire_1282,dangling_wire_1283}),
            .RCLKE(),
            .RCLK(N__23535),
            .RE(N__18207),
            .WCLKE(),
            .WCLK(N__24598),
            .WE(N__8603));
    defparam \line_buffer.mem8_physical .WRITE_MODE=3;
    defparam \line_buffer.mem8_physical .READ_MODE=3;
    defparam \line_buffer.mem8_physical .INIT_F=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem8_physical .INIT_E=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem8_physical .INIT_D=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem8_physical .INIT_C=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem8_physical .INIT_B=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem8_physical .INIT_A=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem8_physical .INIT_9=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem8_physical .INIT_8=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem8_physical .INIT_7=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem8_physical .INIT_6=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem8_physical .INIT_5=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem8_physical .INIT_4=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem8_physical .INIT_3=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem8_physical .INIT_2=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem8_physical .INIT_1=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem8_physical .INIT_0=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    SB_RAM40_4K \line_buffer.mem8_physical  (
            .RDATA({dangling_wire_1284,dangling_wire_1285,dangling_wire_1286,dangling_wire_1287,\line_buffer.n455 ,dangling_wire_1288,dangling_wire_1289,dangling_wire_1290,dangling_wire_1291,dangling_wire_1292,dangling_wire_1293,dangling_wire_1294,\line_buffer.n454 ,dangling_wire_1295,dangling_wire_1296,dangling_wire_1297}),
            .RADDR({N__16153,N__18949,N__19399,N__17077,N__17341,N__16804,N__9088,N__13963,N__18685,N__15643,N__15901}),
            .WADDR({N__12304,N__10405,N__10660,N__10909,N__11167,N__11431,N__11794,N__12052,N__12877,N__9901,N__10156}),
            .MASK({dangling_wire_1298,dangling_wire_1299,dangling_wire_1300,dangling_wire_1301,dangling_wire_1302,dangling_wire_1303,dangling_wire_1304,dangling_wire_1305,dangling_wire_1306,dangling_wire_1307,dangling_wire_1308,dangling_wire_1309,dangling_wire_1310,dangling_wire_1311,dangling_wire_1312,dangling_wire_1313}),
            .WDATA({dangling_wire_1314,dangling_wire_1315,dangling_wire_1316,dangling_wire_1317,N__17687,dangling_wire_1318,dangling_wire_1319,dangling_wire_1320,dangling_wire_1321,dangling_wire_1322,dangling_wire_1323,dangling_wire_1324,N__17789,dangling_wire_1325,dangling_wire_1326,dangling_wire_1327}),
            .RCLKE(),
            .RCLK(N__22844),
            .RE(N__18053),
            .WCLKE(),
            .WCLK(N__24632),
            .WE(N__9382));
    defparam \line_buffer.mem28_physical .WRITE_MODE=3;
    defparam \line_buffer.mem28_physical .READ_MODE=3;
    defparam \line_buffer.mem28_physical .INIT_F=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem28_physical .INIT_E=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem28_physical .INIT_D=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem28_physical .INIT_C=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem28_physical .INIT_B=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem28_physical .INIT_A=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem28_physical .INIT_9=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem28_physical .INIT_8=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem28_physical .INIT_7=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem28_physical .INIT_6=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem28_physical .INIT_5=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem28_physical .INIT_4=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem28_physical .INIT_3=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    defparam \line_buffer.mem28_physical .INIT_2=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    defparam \line_buffer.mem28_physical .INIT_1=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    defparam \line_buffer.mem28_physical .INIT_0=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    SB_RAM40_4K \line_buffer.mem28_physical  (
            .RDATA({dangling_wire_1328,dangling_wire_1329,dangling_wire_1330,dangling_wire_1331,\line_buffer.n556 ,dangling_wire_1332,dangling_wire_1333,dangling_wire_1334,dangling_wire_1335,dangling_wire_1336,dangling_wire_1337,dangling_wire_1338,\line_buffer.n555 ,dangling_wire_1339,dangling_wire_1340,dangling_wire_1341}),
            .RADDR({N__16261,N__19057,N__19507,N__17185,N__17449,N__16912,N__9196,N__14071,N__18793,N__15751,N__16009}),
            .WADDR({N__12412,N__10513,N__10768,N__11017,N__11275,N__11539,N__11902,N__12160,N__12985,N__10009,N__10264}),
            .MASK({dangling_wire_1342,dangling_wire_1343,dangling_wire_1344,dangling_wire_1345,dangling_wire_1346,dangling_wire_1347,dangling_wire_1348,dangling_wire_1349,dangling_wire_1350,dangling_wire_1351,dangling_wire_1352,dangling_wire_1353,dangling_wire_1354,dangling_wire_1355,dangling_wire_1356,dangling_wire_1357}),
            .WDATA({dangling_wire_1358,dangling_wire_1359,dangling_wire_1360,dangling_wire_1361,N__14305,dangling_wire_1362,dangling_wire_1363,dangling_wire_1364,dangling_wire_1365,dangling_wire_1366,dangling_wire_1367,dangling_wire_1368,N__11722,dangling_wire_1369,dangling_wire_1370,dangling_wire_1371}),
            .RCLKE(),
            .RCLK(N__22833),
            .RE(N__18156),
            .WCLKE(),
            .WCLK(N__24610),
            .WE(N__9636));
    defparam \line_buffer.mem18_physical .WRITE_MODE=3;
    defparam \line_buffer.mem18_physical .READ_MODE=3;
    defparam \line_buffer.mem18_physical .INIT_F=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem18_physical .INIT_E=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem18_physical .INIT_D=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem18_physical .INIT_C=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem18_physical .INIT_B=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem18_physical .INIT_A=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem18_physical .INIT_9=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem18_physical .INIT_8=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem18_physical .INIT_7=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem18_physical .INIT_6=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem18_physical .INIT_5=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem18_physical .INIT_4=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem18_physical .INIT_3=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem18_physical .INIT_2=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem18_physical .INIT_1=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem18_physical .INIT_0=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    SB_RAM40_4K \line_buffer.mem18_physical  (
            .RDATA({dangling_wire_1372,dangling_wire_1373,dangling_wire_1374,dangling_wire_1375,\line_buffer.n461 ,dangling_wire_1376,dangling_wire_1377,dangling_wire_1378,dangling_wire_1379,dangling_wire_1380,dangling_wire_1381,dangling_wire_1382,\line_buffer.n460 ,dangling_wire_1383,dangling_wire_1384,dangling_wire_1385}),
            .RADDR({N__16210,N__18988,N__19444,N__17128,N__17398,N__16861,N__9145,N__14032,N__18736,N__15694,N__15946}),
            .WADDR({N__12373,N__10462,N__10705,N__10960,N__11218,N__11476,N__11857,N__12115,N__12916,N__9946,N__10207}),
            .MASK({dangling_wire_1386,dangling_wire_1387,dangling_wire_1388,dangling_wire_1389,dangling_wire_1390,dangling_wire_1391,dangling_wire_1392,dangling_wire_1393,dangling_wire_1394,dangling_wire_1395,dangling_wire_1396,dangling_wire_1397,dangling_wire_1398,dangling_wire_1399,dangling_wire_1400,dangling_wire_1401}),
            .WDATA({dangling_wire_1402,dangling_wire_1403,dangling_wire_1404,dangling_wire_1405,N__17920,dangling_wire_1406,dangling_wire_1407,dangling_wire_1408,dangling_wire_1409,dangling_wire_1410,dangling_wire_1411,dangling_wire_1412,N__19777,dangling_wire_1413,dangling_wire_1414,dangling_wire_1415}),
            .RCLKE(),
            .RCLK(N__23328),
            .RE(N__18109),
            .WCLKE(),
            .WCLK(N__24621),
            .WE(N__14175));
    PRE_IO_GBUF DEBUG_c_2_pad_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__25254),
            .GLOBALBUFFEROUTPUT(DEBUG_c_2_c));
    defparam DEBUG_c_2_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_c_2_pad_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_c_2_pad_iopad (
            .OE(N__25256),
            .DIN(N__25255),
            .DOUT(N__25254),
            .PACKAGEPIN(TVP_CLK));
    defparam DEBUG_c_2_pad_preio.PIN_TYPE=6'b000001;
    defparam DEBUG_c_2_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_c_2_pad_preio (
            .PADOEN(N__25256),
            .PADOUT(N__25255),
            .PADIN(N__25254),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_CLK_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_CLK_pad_iopad.PULLUP=1'b0;
    IO_PAD ADV_CLK_pad_iopad (
            .OE(N__25245),
            .DIN(N__25244),
            .DOUT(N__25243),
            .PACKAGEPIN(ADV_CLK));
    defparam ADV_CLK_pad_preio.PIN_TYPE=6'b011001;
    defparam ADV_CLK_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_CLK_pad_preio (
            .PADOEN(N__25245),
            .PADOUT(N__25244),
            .PADIN(N__25243),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__22910),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_3_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_3_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_3_iopad (
            .OE(N__25236),
            .DIN(N__25235),
            .DOUT(N__25234),
            .PACKAGEPIN(DEBUG[3]));
    defparam DEBUG_pad_3_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_3_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_3_preio (
            .PADOEN(N__25236),
            .PADOUT(N__25235),
            .PADIN(N__25234),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__15601),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_VIDEO_pad_2_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_VIDEO_pad_2_iopad.PULLUP=1'b1;
    IO_PAD TVP_VIDEO_pad_2_iopad (
            .OE(N__25227),
            .DIN(N__25226),
            .DOUT(N__25225),
            .PACKAGEPIN(TVP_VIDEO[2]));
    defparam TVP_VIDEO_pad_2_preio.PIN_TYPE=6'b000001;
    defparam TVP_VIDEO_pad_2_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_VIDEO_pad_2_preio (
            .PADOEN(N__25227),
            .PADOUT(N__25226),
            .PADIN(N__25225),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_VIDEO_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_5_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_5_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_5_iopad (
            .OE(N__25218),
            .DIN(N__25217),
            .DOUT(N__25216),
            .PACKAGEPIN(ADV_G[5]));
    defparam ADV_G_pad_5_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_5_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_5_preio (
            .PADOEN(N__25218),
            .PADOUT(N__25217),
            .PADIN(N__25216),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__21310),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_3_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_3_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_3_iopad (
            .OE(N__25209),
            .DIN(N__25208),
            .DOUT(N__25207),
            .PACKAGEPIN(ADV_R[3]));
    defparam ADV_R_pad_3_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_3_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_3_preio (
            .PADOEN(N__25209),
            .PADOUT(N__25208),
            .PADIN(N__25207),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__23592),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_c_3_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_c_3_pad_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_c_3_pad_iopad (
            .OE(N__25200),
            .DIN(N__25199),
            .DOUT(N__25198),
            .PACKAGEPIN(TVP_VIDEO[5]));
    defparam DEBUG_c_3_pad_preio.PIN_TYPE=6'b000001;
    defparam DEBUG_c_3_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_c_3_pad_preio (
            .PADOEN(N__25200),
            .PADOUT(N__25199),
            .PADIN(N__25198),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DEBUG_c_3_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_0_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_0_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_0_iopad (
            .OE(N__25191),
            .DIN(N__25190),
            .DOUT(N__25189),
            .PACKAGEPIN(ADV_R[0]));
    defparam ADV_R_pad_0_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_0_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_0_preio (
            .PADOEN(N__25191),
            .PADOUT(N__25190),
            .PADIN(N__25189),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__21431),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_2_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_2_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_2_iopad (
            .OE(N__25182),
            .DIN(N__25181),
            .DOUT(N__25180),
            .PACKAGEPIN(DEBUG[2]));
    defparam DEBUG_pad_2_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_2_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_2_preio (
            .PADOEN(N__25182),
            .PADOUT(N__25181),
            .PADIN(N__25180),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8395),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_VIDEO_pad_3_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_VIDEO_pad_3_iopad.PULLUP=1'b1;
    IO_PAD TVP_VIDEO_pad_3_iopad (
            .OE(N__25173),
            .DIN(N__25172),
            .DOUT(N__25171),
            .PACKAGEPIN(TVP_VIDEO[3]));
    defparam TVP_VIDEO_pad_3_preio.PIN_TYPE=6'b000001;
    defparam TVP_VIDEO_pad_3_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_VIDEO_pad_3_preio (
            .PADOEN(N__25173),
            .PADOUT(N__25172),
            .PADIN(N__25171),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_VIDEO_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_4_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_4_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_4_iopad (
            .OE(N__25164),
            .DIN(N__25163),
            .DOUT(N__25162),
            .PACKAGEPIN(ADV_G[4]));
    defparam ADV_G_pad_4_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_4_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_4_preio (
            .PADOEN(N__25164),
            .PADOUT(N__25163),
            .PADIN(N__25162),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__24140),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_5_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_5_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_5_iopad (
            .OE(N__25155),
            .DIN(N__25154),
            .DOUT(N__25153),
            .PACKAGEPIN(ADV_R[5]));
    defparam ADV_R_pad_5_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_5_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_5_preio (
            .PADOEN(N__25155),
            .PADOUT(N__25154),
            .PADIN(N__25153),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__21317),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_1_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_1_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_1_iopad (
            .OE(N__25146),
            .DIN(N__25145),
            .DOUT(N__25144),
            .PACKAGEPIN(DEBUG[1]));
    defparam DEBUG_pad_1_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_1_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_1_preio (
            .PADOEN(N__25146),
            .PADOUT(N__25145),
            .PADIN(N__25144),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8798),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_c_6_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_c_6_pad_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_c_6_pad_iopad (
            .OE(N__25137),
            .DIN(N__25136),
            .DOUT(N__25135),
            .PACKAGEPIN(TVP_VIDEO[8]));
    defparam DEBUG_c_6_pad_preio.PIN_TYPE=6'b000001;
    defparam DEBUG_c_6_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_c_6_pad_preio (
            .PADOEN(N__25137),
            .PADOUT(N__25136),
            .PADIN(N__25135),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DEBUG_c_6_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_1_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_1_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_1_iopad (
            .OE(N__25128),
            .DIN(N__25127),
            .DOUT(N__25126),
            .PACKAGEPIN(ADV_B[1]));
    defparam ADV_B_pad_1_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_1_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_1_preio (
            .PADOEN(N__25128),
            .PADOUT(N__25127),
            .PADIN(N__25126),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__21355),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_SYNC_N_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_SYNC_N_pad_iopad.PULLUP=1'b1;
    IO_PAD ADV_SYNC_N_pad_iopad (
            .OE(N__25119),
            .DIN(N__25118),
            .DOUT(N__25117),
            .PACKAGEPIN(ADV_SYNC_N));
    defparam ADV_SYNC_N_pad_preio.PIN_TYPE=6'b011001;
    defparam ADV_SYNC_N_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_SYNC_N_pad_preio (
            .PADOEN(N__25119),
            .PADOUT(N__25118),
            .PADIN(N__25117),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_6_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_6_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_6_iopad (
            .OE(N__25110),
            .DIN(N__25109),
            .DOUT(N__25108),
            .PACKAGEPIN(ADV_B[6]));
    defparam ADV_B_pad_6_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_6_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_6_preio (
            .PADOEN(N__25110),
            .PADOUT(N__25109),
            .PADIN(N__25108),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__21855),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_6_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_6_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_6_iopad (
            .OE(N__25101),
            .DIN(N__25100),
            .DOUT(N__25099),
            .PACKAGEPIN(DEBUG[6]));
    defparam DEBUG_pad_6_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_6_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_6_preio (
            .PADOEN(N__25101),
            .PADOUT(N__25100),
            .PADIN(N__25099),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__18470),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_0_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_0_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_0_iopad (
            .OE(N__25092),
            .DIN(N__25091),
            .DOUT(N__25090),
            .PACKAGEPIN(ADV_G[0]));
    defparam ADV_G_pad_0_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_0_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_0_preio (
            .PADOEN(N__25092),
            .PADOUT(N__25091),
            .PADIN(N__25090),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__21423),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_1_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_1_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_1_iopad (
            .OE(N__25083),
            .DIN(N__25082),
            .DOUT(N__25081),
            .PACKAGEPIN(ADV_R[1]));
    defparam ADV_R_pad_1_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_1_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_1_preio (
            .PADOEN(N__25083),
            .PADOUT(N__25082),
            .PADIN(N__25081),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__21373),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_5_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_5_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_5_iopad (
            .OE(N__25074),
            .DIN(N__25073),
            .DOUT(N__25072),
            .PACKAGEPIN(DEBUG[5]));
    defparam DEBUG_pad_5_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_5_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_5_preio (
            .PADOEN(N__25074),
            .PADOUT(N__25073),
            .PADIN(N__25072),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__16592),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_7_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_7_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_7_iopad (
            .OE(N__25065),
            .DIN(N__25064),
            .DOUT(N__25063),
            .PACKAGEPIN(ADV_G[7]));
    defparam ADV_G_pad_7_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_7_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_7_preio (
            .PADOEN(N__25065),
            .PADOUT(N__25064),
            .PADIN(N__25063),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__22207),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_6_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_6_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_6_iopad (
            .OE(N__25056),
            .DIN(N__25055),
            .DOUT(N__25054),
            .PACKAGEPIN(ADV_R[6]));
    defparam ADV_R_pad_6_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_6_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_6_preio (
            .PADOEN(N__25056),
            .PADOUT(N__25055),
            .PADIN(N__25054),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__21869),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_BLANK_N_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_BLANK_N_pad_iopad.PULLUP=1'b1;
    IO_PAD ADV_BLANK_N_pad_iopad (
            .OE(N__25047),
            .DIN(N__25046),
            .DOUT(N__25045),
            .PACKAGEPIN(ADV_BLANK_N));
    defparam ADV_BLANK_N_pad_preio.PIN_TYPE=6'b011001;
    defparam ADV_BLANK_N_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_BLANK_N_pad_preio (
            .PADOEN(N__25047),
            .PADOUT(N__25046),
            .PADIN(N__25045),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__18071),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_0_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_0_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_0_iopad (
            .OE(N__25038),
            .DIN(N__25037),
            .DOUT(N__25036),
            .PACKAGEPIN(DEBUG[0]));
    defparam DEBUG_pad_0_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_0_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_0_preio (
            .PADOEN(N__25038),
            .PADOUT(N__25037),
            .PADIN(N__25036),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9479),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_2_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_2_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_2_iopad (
            .OE(N__25029),
            .DIN(N__25028),
            .DOUT(N__25027),
            .PACKAGEPIN(ADV_B[2]));
    defparam ADV_B_pad_2_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_2_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_2_preio (
            .PADOEN(N__25029),
            .PADOUT(N__25028),
            .PADIN(N__25027),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__22243),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_c_7_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_c_7_pad_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_c_7_pad_iopad (
            .OE(N__25020),
            .DIN(N__25019),
            .DOUT(N__25018),
            .PACKAGEPIN(TVP_VIDEO[9]));
    defparam DEBUG_c_7_pad_preio.PIN_TYPE=6'b000001;
    defparam DEBUG_c_7_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_c_7_pad_preio (
            .PADOEN(N__25020),
            .PADOUT(N__25019),
            .PADIN(N__25018),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DEBUG_c_7_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_c_1_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_c_1_pad_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_c_1_pad_iopad (
            .OE(N__25011),
            .DIN(N__25010),
            .DOUT(N__25009),
            .PACKAGEPIN(TVP_HSYNC));
    defparam DEBUG_c_1_pad_preio.PIN_TYPE=6'b000001;
    defparam DEBUG_c_1_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_c_1_pad_preio (
            .PADOEN(N__25011),
            .PADOUT(N__25010),
            .PADIN(N__25009),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DEBUG_c_1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_c_5_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_c_5_pad_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_c_5_pad_iopad (
            .OE(N__25002),
            .DIN(N__25001),
            .DOUT(N__25000),
            .PACKAGEPIN(TVP_VIDEO[7]));
    defparam DEBUG_c_5_pad_preio.PIN_TYPE=6'b000001;
    defparam DEBUG_c_5_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_c_5_pad_preio (
            .PADOEN(N__25002),
            .PADOUT(N__25001),
            .PADIN(N__25000),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DEBUG_c_5_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_7_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_7_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_7_iopad (
            .OE(N__24993),
            .DIN(N__24992),
            .DOUT(N__24991),
            .PACKAGEPIN(ADV_B[7]));
    defparam ADV_B_pad_7_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_7_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_7_preio (
            .PADOEN(N__24993),
            .PADOUT(N__24992),
            .PADIN(N__24991),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__22197),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam LED_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam LED_pad_iopad.PULLUP=1'b1;
    IO_PAD LED_pad_iopad (
            .OE(N__24984),
            .DIN(N__24983),
            .DOUT(N__24982),
            .PACKAGEPIN(LED));
    defparam LED_pad_preio.PIN_TYPE=6'b011001;
    defparam LED_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO LED_pad_preio (
            .PADOEN(N__24984),
            .PADOUT(N__24983),
            .PADIN(N__24982),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8816),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_VIDEO_pad_4_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_VIDEO_pad_4_iopad.PULLUP=1'b1;
    IO_PAD TVP_VIDEO_pad_4_iopad (
            .OE(N__24975),
            .DIN(N__24974),
            .DOUT(N__24973),
            .PACKAGEPIN(TVP_VIDEO[4]));
    defparam TVP_VIDEO_pad_4_preio.PIN_TYPE=6'b000001;
    defparam TVP_VIDEO_pad_4_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_VIDEO_pad_4_preio (
            .PADOEN(N__24975),
            .PADOUT(N__24974),
            .PADIN(N__24973),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_VIDEO_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_3_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_3_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_3_iopad (
            .OE(N__24966),
            .DIN(N__24965),
            .DOUT(N__24964),
            .PACKAGEPIN(ADV_G[3]));
    defparam ADV_G_pad_3_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_3_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_3_preio (
            .PADOEN(N__24966),
            .PADOUT(N__24965),
            .PADIN(N__24964),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__23606),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_HSYNC_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_HSYNC_pad_iopad.PULLUP=1'b0;
    IO_PAD ADV_HSYNC_pad_iopad (
            .OE(N__24957),
            .DIN(N__24956),
            .DOUT(N__24955),
            .PACKAGEPIN(ADV_HSYNC));
    defparam ADV_HSYNC_pad_preio.PIN_TYPE=6'b011001;
    defparam ADV_HSYNC_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_HSYNC_pad_preio (
            .PADOEN(N__24957),
            .PADOUT(N__24956),
            .PADIN(N__24955),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__16379),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_2_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_2_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_2_iopad (
            .OE(N__24948),
            .DIN(N__24947),
            .DOUT(N__24946),
            .PACKAGEPIN(ADV_R[2]));
    defparam ADV_R_pad_2_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_2_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_2_preio (
            .PADOEN(N__24948),
            .PADOUT(N__24947),
            .PADIN(N__24946),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__22258),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_c_0_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_c_0_pad_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_c_0_pad_iopad (
            .OE(N__24939),
            .DIN(N__24938),
            .DOUT(N__24937),
            .PACKAGEPIN(TVP_VSYNC));
    defparam DEBUG_c_0_pad_preio.PIN_TYPE=6'b000001;
    defparam DEBUG_c_0_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_c_0_pad_preio (
            .PADOEN(N__24939),
            .PADOUT(N__24938),
            .PADIN(N__24937),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DEBUG_c_0_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_4_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_4_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_4_iopad (
            .OE(N__24930),
            .DIN(N__24929),
            .DOUT(N__24928),
            .PACKAGEPIN(ADV_B[4]));
    defparam ADV_B_pad_4_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_4_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_4_preio (
            .PADOEN(N__24930),
            .PADOUT(N__24929),
            .PADIN(N__24928),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__24136),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_4_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_4_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_4_iopad (
            .OE(N__24921),
            .DIN(N__24920),
            .DOUT(N__24919),
            .PACKAGEPIN(DEBUG[4]));
    defparam DEBUG_pad_4_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_4_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_4_preio (
            .PADOEN(N__24921),
            .PADOUT(N__24920),
            .PADIN(N__24919),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__15575),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_6_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_6_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_6_iopad (
            .OE(N__24912),
            .DIN(N__24911),
            .DOUT(N__24910),
            .PACKAGEPIN(ADV_G[6]));
    defparam ADV_G_pad_6_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_6_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_6_preio (
            .PADOEN(N__24912),
            .PADOUT(N__24911),
            .PADIN(N__24910),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__21862),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_7_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_7_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_7_iopad (
            .OE(N__24903),
            .DIN(N__24902),
            .DOUT(N__24901),
            .PACKAGEPIN(ADV_R[7]));
    defparam ADV_R_pad_7_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_7_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_7_preio (
            .PADOEN(N__24903),
            .PADOUT(N__24902),
            .PADIN(N__24901),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__22208),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_3_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_3_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_3_iopad (
            .OE(N__24894),
            .DIN(N__24893),
            .DOUT(N__24892),
            .PACKAGEPIN(ADV_B[3]));
    defparam ADV_B_pad_3_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_3_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_3_preio (
            .PADOEN(N__24894),
            .PADOUT(N__24893),
            .PADIN(N__24892),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__23602),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_4_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_4_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_4_iopad (
            .OE(N__24885),
            .DIN(N__24884),
            .DOUT(N__24883),
            .PACKAGEPIN(ADV_R[4]));
    defparam ADV_R_pad_4_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_4_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_4_preio (
            .PADOEN(N__24885),
            .PADOUT(N__24884),
            .PADIN(N__24883),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__24126),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_0_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_0_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_0_iopad (
            .OE(N__24876),
            .DIN(N__24875),
            .DOUT(N__24874),
            .PACKAGEPIN(ADV_B[0]));
    defparam ADV_B_pad_0_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_0_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_0_preio (
            .PADOEN(N__24876),
            .PADOUT(N__24875),
            .PADIN(N__24874),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__21430),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_2_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_2_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_2_iopad (
            .OE(N__24867),
            .DIN(N__24866),
            .DOUT(N__24865),
            .PACKAGEPIN(ADV_G[2]));
    defparam ADV_G_pad_2_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_2_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_2_preio (
            .PADOEN(N__24867),
            .PADOUT(N__24866),
            .PADIN(N__24865),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__22268),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_VSYNC_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_VSYNC_pad_iopad.PULLUP=1'b0;
    IO_PAD ADV_VSYNC_pad_iopad (
            .OE(N__24858),
            .DIN(N__24857),
            .DOUT(N__24856),
            .PACKAGEPIN(ADV_VSYNC));
    defparam ADV_VSYNC_pad_preio.PIN_TYPE=6'b011001;
    defparam ADV_VSYNC_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_VSYNC_pad_preio (
            .PADOEN(N__24858),
            .PADOUT(N__24857),
            .PADIN(N__24856),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__20420),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_c_4_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_c_4_pad_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_c_4_pad_iopad (
            .OE(N__24849),
            .DIN(N__24848),
            .DOUT(N__24847),
            .PACKAGEPIN(TVP_VIDEO[6]));
    defparam DEBUG_c_4_pad_preio.PIN_TYPE=6'b000001;
    defparam DEBUG_c_4_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_c_4_pad_preio (
            .PADOEN(N__24849),
            .PADOUT(N__24848),
            .PADIN(N__24847),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DEBUG_c_4_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_5_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_5_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_5_iopad (
            .OE(N__24840),
            .DIN(N__24839),
            .DOUT(N__24838),
            .PACKAGEPIN(ADV_B[5]));
    defparam ADV_B_pad_5_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_5_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_5_preio (
            .PADOEN(N__24840),
            .PADOUT(N__24839),
            .PADIN(N__24838),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__21303),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_7_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_7_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_7_iopad (
            .OE(N__24831),
            .DIN(N__24830),
            .DOUT(N__24829),
            .PACKAGEPIN(DEBUG[7]));
    defparam DEBUG_pad_7_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_7_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_7_preio (
            .PADOEN(N__24831),
            .PADOUT(N__24830),
            .PADIN(N__24829),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__24683),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_1_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_1_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_1_iopad (
            .OE(N__24822),
            .DIN(N__24821),
            .DOUT(N__24820),
            .PACKAGEPIN(ADV_G[1]));
    defparam ADV_G_pad_1_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_1_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_1_preio (
            .PADOEN(N__24822),
            .PADOUT(N__24821),
            .PADIN(N__24820),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__21377),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    SRMux I__6017 (
            .O(N__24803),
            .I(N__24800));
    LocalMux I__6016 (
            .O(N__24800),
            .I(N__24793));
    SRMux I__6015 (
            .O(N__24799),
            .I(N__24789));
    SRMux I__6014 (
            .O(N__24798),
            .I(N__24786));
    SRMux I__6013 (
            .O(N__24797),
            .I(N__24781));
    SRMux I__6012 (
            .O(N__24796),
            .I(N__24778));
    Span4Mux_h I__6011 (
            .O(N__24793),
            .I(N__24775));
    SRMux I__6010 (
            .O(N__24792),
            .I(N__24772));
    LocalMux I__6009 (
            .O(N__24789),
            .I(N__24769));
    LocalMux I__6008 (
            .O(N__24786),
            .I(N__24766));
    SRMux I__6007 (
            .O(N__24785),
            .I(N__24763));
    SRMux I__6006 (
            .O(N__24784),
            .I(N__24760));
    LocalMux I__6005 (
            .O(N__24781),
            .I(N__24751));
    LocalMux I__6004 (
            .O(N__24778),
            .I(N__24751));
    Span4Mux_h I__6003 (
            .O(N__24775),
            .I(N__24751));
    LocalMux I__6002 (
            .O(N__24772),
            .I(N__24751));
    Span4Mux_v I__6001 (
            .O(N__24769),
            .I(N__24748));
    Span4Mux_v I__6000 (
            .O(N__24766),
            .I(N__24741));
    LocalMux I__5999 (
            .O(N__24763),
            .I(N__24741));
    LocalMux I__5998 (
            .O(N__24760),
            .I(N__24741));
    Span4Mux_v I__5997 (
            .O(N__24751),
            .I(N__24738));
    Sp12to4 I__5996 (
            .O(N__24748),
            .I(N__24733));
    Sp12to4 I__5995 (
            .O(N__24741),
            .I(N__24733));
    Odrv4 I__5994 (
            .O(N__24738),
            .I(\transmit_module.n2367 ));
    Odrv12 I__5993 (
            .O(N__24733),
            .I(\transmit_module.n2367 ));
    InMux I__5992 (
            .O(N__24728),
            .I(N__24725));
    LocalMux I__5991 (
            .O(N__24725),
            .I(N__24722));
    Odrv4 I__5990 (
            .O(N__24722),
            .I(\tvp_video_buffer.BUFFER_1_9 ));
    InMux I__5989 (
            .O(N__24719),
            .I(N__24716));
    LocalMux I__5988 (
            .O(N__24716),
            .I(N__24713));
    Span12Mux_h I__5987 (
            .O(N__24713),
            .I(N__24710));
    Span12Mux_v I__5986 (
            .O(N__24710),
            .I(N__24707));
    Odrv12 I__5985 (
            .O(N__24707),
            .I(\line_buffer.n526 ));
    InMux I__5984 (
            .O(N__24704),
            .I(N__24701));
    LocalMux I__5983 (
            .O(N__24701),
            .I(N__24698));
    Span4Mux_h I__5982 (
            .O(N__24698),
            .I(N__24695));
    Span4Mux_v I__5981 (
            .O(N__24695),
            .I(N__24692));
    Odrv4 I__5980 (
            .O(N__24692),
            .I(\line_buffer.n518 ));
    InMux I__5979 (
            .O(N__24689),
            .I(N__24686));
    LocalMux I__5978 (
            .O(N__24686),
            .I(\line_buffer.n3479 ));
    IoInMux I__5977 (
            .O(N__24683),
            .I(N__24680));
    LocalMux I__5976 (
            .O(N__24680),
            .I(N__24677));
    IoSpan4Mux I__5975 (
            .O(N__24677),
            .I(N__24674));
    Span4Mux_s0_h I__5974 (
            .O(N__24674),
            .I(N__24671));
    Sp12to4 I__5973 (
            .O(N__24671),
            .I(N__24668));
    Span12Mux_s11_h I__5972 (
            .O(N__24668),
            .I(N__24665));
    Span12Mux_v I__5971 (
            .O(N__24665),
            .I(N__24661));
    InMux I__5970 (
            .O(N__24664),
            .I(N__24658));
    Span12Mux_h I__5969 (
            .O(N__24661),
            .I(N__24655));
    LocalMux I__5968 (
            .O(N__24658),
            .I(N__24652));
    Odrv12 I__5967 (
            .O(N__24655),
            .I(DEBUG_c_7_c));
    Odrv4 I__5966 (
            .O(N__24652),
            .I(DEBUG_c_7_c));
    InMux I__5965 (
            .O(N__24647),
            .I(N__24644));
    LocalMux I__5964 (
            .O(N__24644),
            .I(\tvp_video_buffer.BUFFER_0_9 ));
    InMux I__5963 (
            .O(N__24641),
            .I(N__24638));
    LocalMux I__5962 (
            .O(N__24638),
            .I(N__24633));
    ClkMux I__5961 (
            .O(N__24637),
            .I(N__24419));
    ClkMux I__5960 (
            .O(N__24636),
            .I(N__24419));
    Glb2LocalMux I__5959 (
            .O(N__24633),
            .I(N__24419));
    ClkMux I__5958 (
            .O(N__24632),
            .I(N__24419));
    ClkMux I__5957 (
            .O(N__24631),
            .I(N__24419));
    ClkMux I__5956 (
            .O(N__24630),
            .I(N__24419));
    ClkMux I__5955 (
            .O(N__24629),
            .I(N__24419));
    ClkMux I__5954 (
            .O(N__24628),
            .I(N__24419));
    ClkMux I__5953 (
            .O(N__24627),
            .I(N__24419));
    ClkMux I__5952 (
            .O(N__24626),
            .I(N__24419));
    ClkMux I__5951 (
            .O(N__24625),
            .I(N__24419));
    ClkMux I__5950 (
            .O(N__24624),
            .I(N__24419));
    ClkMux I__5949 (
            .O(N__24623),
            .I(N__24419));
    ClkMux I__5948 (
            .O(N__24622),
            .I(N__24419));
    ClkMux I__5947 (
            .O(N__24621),
            .I(N__24419));
    ClkMux I__5946 (
            .O(N__24620),
            .I(N__24419));
    ClkMux I__5945 (
            .O(N__24619),
            .I(N__24419));
    ClkMux I__5944 (
            .O(N__24618),
            .I(N__24419));
    ClkMux I__5943 (
            .O(N__24617),
            .I(N__24419));
    ClkMux I__5942 (
            .O(N__24616),
            .I(N__24419));
    ClkMux I__5941 (
            .O(N__24615),
            .I(N__24419));
    ClkMux I__5940 (
            .O(N__24614),
            .I(N__24419));
    ClkMux I__5939 (
            .O(N__24613),
            .I(N__24419));
    ClkMux I__5938 (
            .O(N__24612),
            .I(N__24419));
    ClkMux I__5937 (
            .O(N__24611),
            .I(N__24419));
    ClkMux I__5936 (
            .O(N__24610),
            .I(N__24419));
    ClkMux I__5935 (
            .O(N__24609),
            .I(N__24419));
    ClkMux I__5934 (
            .O(N__24608),
            .I(N__24419));
    ClkMux I__5933 (
            .O(N__24607),
            .I(N__24419));
    ClkMux I__5932 (
            .O(N__24606),
            .I(N__24419));
    ClkMux I__5931 (
            .O(N__24605),
            .I(N__24419));
    ClkMux I__5930 (
            .O(N__24604),
            .I(N__24419));
    ClkMux I__5929 (
            .O(N__24603),
            .I(N__24419));
    ClkMux I__5928 (
            .O(N__24602),
            .I(N__24419));
    ClkMux I__5927 (
            .O(N__24601),
            .I(N__24419));
    ClkMux I__5926 (
            .O(N__24600),
            .I(N__24419));
    ClkMux I__5925 (
            .O(N__24599),
            .I(N__24419));
    ClkMux I__5924 (
            .O(N__24598),
            .I(N__24419));
    ClkMux I__5923 (
            .O(N__24597),
            .I(N__24419));
    ClkMux I__5922 (
            .O(N__24596),
            .I(N__24419));
    ClkMux I__5921 (
            .O(N__24595),
            .I(N__24419));
    ClkMux I__5920 (
            .O(N__24594),
            .I(N__24419));
    ClkMux I__5919 (
            .O(N__24593),
            .I(N__24419));
    ClkMux I__5918 (
            .O(N__24592),
            .I(N__24419));
    ClkMux I__5917 (
            .O(N__24591),
            .I(N__24419));
    ClkMux I__5916 (
            .O(N__24590),
            .I(N__24419));
    ClkMux I__5915 (
            .O(N__24589),
            .I(N__24419));
    ClkMux I__5914 (
            .O(N__24588),
            .I(N__24419));
    ClkMux I__5913 (
            .O(N__24587),
            .I(N__24419));
    ClkMux I__5912 (
            .O(N__24586),
            .I(N__24419));
    ClkMux I__5911 (
            .O(N__24585),
            .I(N__24419));
    ClkMux I__5910 (
            .O(N__24584),
            .I(N__24419));
    ClkMux I__5909 (
            .O(N__24583),
            .I(N__24419));
    ClkMux I__5908 (
            .O(N__24582),
            .I(N__24419));
    ClkMux I__5907 (
            .O(N__24581),
            .I(N__24419));
    ClkMux I__5906 (
            .O(N__24580),
            .I(N__24419));
    ClkMux I__5905 (
            .O(N__24579),
            .I(N__24419));
    ClkMux I__5904 (
            .O(N__24578),
            .I(N__24419));
    ClkMux I__5903 (
            .O(N__24577),
            .I(N__24419));
    ClkMux I__5902 (
            .O(N__24576),
            .I(N__24419));
    ClkMux I__5901 (
            .O(N__24575),
            .I(N__24419));
    ClkMux I__5900 (
            .O(N__24574),
            .I(N__24419));
    ClkMux I__5899 (
            .O(N__24573),
            .I(N__24419));
    ClkMux I__5898 (
            .O(N__24572),
            .I(N__24419));
    ClkMux I__5897 (
            .O(N__24571),
            .I(N__24419));
    ClkMux I__5896 (
            .O(N__24570),
            .I(N__24419));
    ClkMux I__5895 (
            .O(N__24569),
            .I(N__24419));
    ClkMux I__5894 (
            .O(N__24568),
            .I(N__24419));
    ClkMux I__5893 (
            .O(N__24567),
            .I(N__24419));
    ClkMux I__5892 (
            .O(N__24566),
            .I(N__24419));
    ClkMux I__5891 (
            .O(N__24565),
            .I(N__24419));
    ClkMux I__5890 (
            .O(N__24564),
            .I(N__24419));
    GlobalMux I__5889 (
            .O(N__24419),
            .I(N__24416));
    gio2CtrlBuf I__5888 (
            .O(N__24416),
            .I(DEBUG_c_2_c));
    InMux I__5887 (
            .O(N__24413),
            .I(N__24410));
    LocalMux I__5886 (
            .O(N__24410),
            .I(N__24407));
    Span4Mux_h I__5885 (
            .O(N__24407),
            .I(N__24404));
    Odrv4 I__5884 (
            .O(N__24404),
            .I(\line_buffer.n459 ));
    InMux I__5883 (
            .O(N__24401),
            .I(N__24398));
    LocalMux I__5882 (
            .O(N__24398),
            .I(N__24395));
    Sp12to4 I__5881 (
            .O(N__24395),
            .I(N__24392));
    Span12Mux_v I__5880 (
            .O(N__24392),
            .I(N__24389));
    Odrv12 I__5879 (
            .O(N__24389),
            .I(\line_buffer.n451 ));
    InMux I__5878 (
            .O(N__24386),
            .I(N__24381));
    InMux I__5877 (
            .O(N__24385),
            .I(N__24374));
    InMux I__5876 (
            .O(N__24384),
            .I(N__24370));
    LocalMux I__5875 (
            .O(N__24381),
            .I(N__24364));
    InMux I__5874 (
            .O(N__24380),
            .I(N__24359));
    InMux I__5873 (
            .O(N__24379),
            .I(N__24359));
    InMux I__5872 (
            .O(N__24378),
            .I(N__24354));
    InMux I__5871 (
            .O(N__24377),
            .I(N__24351));
    LocalMux I__5870 (
            .O(N__24374),
            .I(N__24348));
    InMux I__5869 (
            .O(N__24373),
            .I(N__24345));
    LocalMux I__5868 (
            .O(N__24370),
            .I(N__24332));
    InMux I__5867 (
            .O(N__24369),
            .I(N__24329));
    InMux I__5866 (
            .O(N__24368),
            .I(N__24326));
    InMux I__5865 (
            .O(N__24367),
            .I(N__24323));
    Span4Mux_v I__5864 (
            .O(N__24364),
            .I(N__24320));
    LocalMux I__5863 (
            .O(N__24359),
            .I(N__24317));
    InMux I__5862 (
            .O(N__24358),
            .I(N__24314));
    InMux I__5861 (
            .O(N__24357),
            .I(N__24311));
    LocalMux I__5860 (
            .O(N__24354),
            .I(N__24307));
    LocalMux I__5859 (
            .O(N__24351),
            .I(N__24304));
    Span4Mux_v I__5858 (
            .O(N__24348),
            .I(N__24299));
    LocalMux I__5857 (
            .O(N__24345),
            .I(N__24299));
    InMux I__5856 (
            .O(N__24344),
            .I(N__24296));
    InMux I__5855 (
            .O(N__24343),
            .I(N__24291));
    InMux I__5854 (
            .O(N__24342),
            .I(N__24291));
    InMux I__5853 (
            .O(N__24341),
            .I(N__24285));
    InMux I__5852 (
            .O(N__24340),
            .I(N__24285));
    InMux I__5851 (
            .O(N__24339),
            .I(N__24282));
    InMux I__5850 (
            .O(N__24338),
            .I(N__24279));
    InMux I__5849 (
            .O(N__24337),
            .I(N__24276));
    InMux I__5848 (
            .O(N__24336),
            .I(N__24273));
    InMux I__5847 (
            .O(N__24335),
            .I(N__24270));
    Span4Mux_v I__5846 (
            .O(N__24332),
            .I(N__24265));
    LocalMux I__5845 (
            .O(N__24329),
            .I(N__24265));
    LocalMux I__5844 (
            .O(N__24326),
            .I(N__24262));
    LocalMux I__5843 (
            .O(N__24323),
            .I(N__24254));
    Span4Mux_h I__5842 (
            .O(N__24320),
            .I(N__24254));
    Span4Mux_v I__5841 (
            .O(N__24317),
            .I(N__24254));
    LocalMux I__5840 (
            .O(N__24314),
            .I(N__24251));
    LocalMux I__5839 (
            .O(N__24311),
            .I(N__24248));
    InMux I__5838 (
            .O(N__24310),
            .I(N__24245));
    Span4Mux_h I__5837 (
            .O(N__24307),
            .I(N__24242));
    Span4Mux_v I__5836 (
            .O(N__24304),
            .I(N__24233));
    Span4Mux_v I__5835 (
            .O(N__24299),
            .I(N__24233));
    LocalMux I__5834 (
            .O(N__24296),
            .I(N__24233));
    LocalMux I__5833 (
            .O(N__24291),
            .I(N__24233));
    InMux I__5832 (
            .O(N__24290),
            .I(N__24230));
    LocalMux I__5831 (
            .O(N__24285),
            .I(N__24227));
    LocalMux I__5830 (
            .O(N__24282),
            .I(N__24224));
    LocalMux I__5829 (
            .O(N__24279),
            .I(N__24217));
    LocalMux I__5828 (
            .O(N__24276),
            .I(N__24217));
    LocalMux I__5827 (
            .O(N__24273),
            .I(N__24217));
    LocalMux I__5826 (
            .O(N__24270),
            .I(N__24210));
    Span4Mux_v I__5825 (
            .O(N__24265),
            .I(N__24210));
    Span4Mux_h I__5824 (
            .O(N__24262),
            .I(N__24210));
    InMux I__5823 (
            .O(N__24261),
            .I(N__24207));
    Span4Mux_h I__5822 (
            .O(N__24254),
            .I(N__24202));
    Span4Mux_v I__5821 (
            .O(N__24251),
            .I(N__24202));
    Span4Mux_h I__5820 (
            .O(N__24248),
            .I(N__24197));
    LocalMux I__5819 (
            .O(N__24245),
            .I(N__24197));
    Span4Mux_v I__5818 (
            .O(N__24242),
            .I(N__24194));
    Sp12to4 I__5817 (
            .O(N__24233),
            .I(N__24189));
    LocalMux I__5816 (
            .O(N__24230),
            .I(N__24189));
    Span4Mux_h I__5815 (
            .O(N__24227),
            .I(N__24184));
    Span4Mux_h I__5814 (
            .O(N__24224),
            .I(N__24184));
    Span12Mux_h I__5813 (
            .O(N__24217),
            .I(N__24181));
    Span4Mux_h I__5812 (
            .O(N__24210),
            .I(N__24178));
    LocalMux I__5811 (
            .O(N__24207),
            .I(TX_ADDR_11));
    Odrv4 I__5810 (
            .O(N__24202),
            .I(TX_ADDR_11));
    Odrv4 I__5809 (
            .O(N__24197),
            .I(TX_ADDR_11));
    Odrv4 I__5808 (
            .O(N__24194),
            .I(TX_ADDR_11));
    Odrv12 I__5807 (
            .O(N__24189),
            .I(TX_ADDR_11));
    Odrv4 I__5806 (
            .O(N__24184),
            .I(TX_ADDR_11));
    Odrv12 I__5805 (
            .O(N__24181),
            .I(TX_ADDR_11));
    Odrv4 I__5804 (
            .O(N__24178),
            .I(TX_ADDR_11));
    InMux I__5803 (
            .O(N__24161),
            .I(N__24158));
    LocalMux I__5802 (
            .O(N__24158),
            .I(N__24155));
    Odrv12 I__5801 (
            .O(N__24155),
            .I(\line_buffer.n3518 ));
    InMux I__5800 (
            .O(N__24152),
            .I(N__24149));
    LocalMux I__5799 (
            .O(N__24149),
            .I(N__24146));
    Span4Mux_v I__5798 (
            .O(N__24146),
            .I(N__24143));
    Odrv4 I__5797 (
            .O(N__24143),
            .I(TX_DATA_4));
    IoInMux I__5796 (
            .O(N__24140),
            .I(N__24137));
    LocalMux I__5795 (
            .O(N__24137),
            .I(N__24133));
    IoInMux I__5794 (
            .O(N__24136),
            .I(N__24130));
    IoSpan4Mux I__5793 (
            .O(N__24133),
            .I(N__24127));
    LocalMux I__5792 (
            .O(N__24130),
            .I(N__24123));
    Span4Mux_s2_v I__5791 (
            .O(N__24127),
            .I(N__24120));
    IoInMux I__5790 (
            .O(N__24126),
            .I(N__24117));
    IoSpan4Mux I__5789 (
            .O(N__24123),
            .I(N__24114));
    Sp12to4 I__5788 (
            .O(N__24120),
            .I(N__24111));
    LocalMux I__5787 (
            .O(N__24117),
            .I(N__24108));
    Span4Mux_s0_v I__5786 (
            .O(N__24114),
            .I(N__24105));
    Span12Mux_s7_v I__5785 (
            .O(N__24111),
            .I(N__24100));
    Span12Mux_s7_h I__5784 (
            .O(N__24108),
            .I(N__24100));
    Span4Mux_v I__5783 (
            .O(N__24105),
            .I(N__24097));
    Span12Mux_h I__5782 (
            .O(N__24100),
            .I(N__24094));
    Span4Mux_v I__5781 (
            .O(N__24097),
            .I(N__24091));
    Odrv12 I__5780 (
            .O(N__24094),
            .I(n1810));
    Odrv4 I__5779 (
            .O(N__24091),
            .I(n1810));
    InMux I__5778 (
            .O(N__24086),
            .I(N__24083));
    LocalMux I__5777 (
            .O(N__24083),
            .I(N__24080));
    Span12Mux_h I__5776 (
            .O(N__24080),
            .I(N__24077));
    Span12Mux_v I__5775 (
            .O(N__24077),
            .I(N__24074));
    Odrv12 I__5774 (
            .O(N__24074),
            .I(\line_buffer.n554 ));
    InMux I__5773 (
            .O(N__24071),
            .I(N__24068));
    LocalMux I__5772 (
            .O(N__24068),
            .I(N__24065));
    Span12Mux_h I__5771 (
            .O(N__24065),
            .I(N__24062));
    Span12Mux_h I__5770 (
            .O(N__24062),
            .I(N__24059));
    Odrv12 I__5769 (
            .O(N__24059),
            .I(\line_buffer.n562 ));
    InMux I__5768 (
            .O(N__24056),
            .I(N__24053));
    LocalMux I__5767 (
            .O(N__24053),
            .I(\line_buffer.n3585 ));
    InMux I__5766 (
            .O(N__24050),
            .I(N__24047));
    LocalMux I__5765 (
            .O(N__24047),
            .I(N__24044));
    Span4Mux_v I__5764 (
            .O(N__24044),
            .I(N__24041));
    Span4Mux_v I__5763 (
            .O(N__24041),
            .I(N__24038));
    Sp12to4 I__5762 (
            .O(N__24038),
            .I(N__24035));
    Odrv12 I__5761 (
            .O(N__24035),
            .I(\line_buffer.n558 ));
    InMux I__5760 (
            .O(N__24032),
            .I(N__24029));
    LocalMux I__5759 (
            .O(N__24029),
            .I(N__24026));
    Span4Mux_v I__5758 (
            .O(N__24026),
            .I(N__24023));
    Span4Mux_h I__5757 (
            .O(N__24023),
            .I(N__24020));
    Odrv4 I__5756 (
            .O(N__24020),
            .I(\line_buffer.n550 ));
    CascadeMux I__5755 (
            .O(N__24017),
            .I(N__24012));
    InMux I__5754 (
            .O(N__24016),
            .I(N__24005));
    InMux I__5753 (
            .O(N__24015),
            .I(N__24002));
    InMux I__5752 (
            .O(N__24012),
            .I(N__23999));
    InMux I__5751 (
            .O(N__24011),
            .I(N__23993));
    InMux I__5750 (
            .O(N__24010),
            .I(N__23990));
    CascadeMux I__5749 (
            .O(N__24009),
            .I(N__23987));
    CascadeMux I__5748 (
            .O(N__24008),
            .I(N__23983));
    LocalMux I__5747 (
            .O(N__24005),
            .I(N__23980));
    LocalMux I__5746 (
            .O(N__24002),
            .I(N__23975));
    LocalMux I__5745 (
            .O(N__23999),
            .I(N__23975));
    InMux I__5744 (
            .O(N__23998),
            .I(N__23971));
    InMux I__5743 (
            .O(N__23997),
            .I(N__23968));
    InMux I__5742 (
            .O(N__23996),
            .I(N__23965));
    LocalMux I__5741 (
            .O(N__23993),
            .I(N__23960));
    LocalMux I__5740 (
            .O(N__23990),
            .I(N__23960));
    InMux I__5739 (
            .O(N__23987),
            .I(N__23957));
    InMux I__5738 (
            .O(N__23986),
            .I(N__23954));
    InMux I__5737 (
            .O(N__23983),
            .I(N__23951));
    Span4Mux_v I__5736 (
            .O(N__23980),
            .I(N__23946));
    Span4Mux_h I__5735 (
            .O(N__23975),
            .I(N__23943));
    InMux I__5734 (
            .O(N__23974),
            .I(N__23940));
    LocalMux I__5733 (
            .O(N__23971),
            .I(N__23937));
    LocalMux I__5732 (
            .O(N__23968),
            .I(N__23928));
    LocalMux I__5731 (
            .O(N__23965),
            .I(N__23928));
    Span4Mux_h I__5730 (
            .O(N__23960),
            .I(N__23928));
    LocalMux I__5729 (
            .O(N__23957),
            .I(N__23928));
    LocalMux I__5728 (
            .O(N__23954),
            .I(N__23923));
    LocalMux I__5727 (
            .O(N__23951),
            .I(N__23923));
    InMux I__5726 (
            .O(N__23950),
            .I(N__23920));
    InMux I__5725 (
            .O(N__23949),
            .I(N__23917));
    Span4Mux_h I__5724 (
            .O(N__23946),
            .I(N__23914));
    Span4Mux_h I__5723 (
            .O(N__23943),
            .I(N__23911));
    LocalMux I__5722 (
            .O(N__23940),
            .I(N__23902));
    Span4Mux_v I__5721 (
            .O(N__23937),
            .I(N__23902));
    Span4Mux_v I__5720 (
            .O(N__23928),
            .I(N__23902));
    Span4Mux_h I__5719 (
            .O(N__23923),
            .I(N__23902));
    LocalMux I__5718 (
            .O(N__23920),
            .I(N__23899));
    LocalMux I__5717 (
            .O(N__23917),
            .I(TX_ADDR_13));
    Odrv4 I__5716 (
            .O(N__23914),
            .I(TX_ADDR_13));
    Odrv4 I__5715 (
            .O(N__23911),
            .I(TX_ADDR_13));
    Odrv4 I__5714 (
            .O(N__23902),
            .I(TX_ADDR_13));
    Odrv4 I__5713 (
            .O(N__23899),
            .I(TX_ADDR_13));
    InMux I__5712 (
            .O(N__23888),
            .I(N__23885));
    LocalMux I__5711 (
            .O(N__23885),
            .I(N__23882));
    Odrv4 I__5710 (
            .O(N__23882),
            .I(\line_buffer.n3482 ));
    CascadeMux I__5709 (
            .O(N__23879),
            .I(\line_buffer.n3567_cascade_ ));
    InMux I__5708 (
            .O(N__23876),
            .I(N__23873));
    LocalMux I__5707 (
            .O(N__23873),
            .I(\line_buffer.n3483 ));
    InMux I__5706 (
            .O(N__23870),
            .I(N__23867));
    LocalMux I__5705 (
            .O(N__23867),
            .I(N__23864));
    Span4Mux_v I__5704 (
            .O(N__23864),
            .I(N__23861));
    Span4Mux_v I__5703 (
            .O(N__23861),
            .I(N__23858));
    Span4Mux_v I__5702 (
            .O(N__23858),
            .I(N__23855));
    Sp12to4 I__5701 (
            .O(N__23855),
            .I(N__23852));
    Odrv12 I__5700 (
            .O(N__23852),
            .I(\line_buffer.n559 ));
    CascadeMux I__5699 (
            .O(N__23849),
            .I(N__23837));
    CascadeMux I__5698 (
            .O(N__23848),
            .I(N__23834));
    CascadeMux I__5697 (
            .O(N__23847),
            .I(N__23828));
    CascadeMux I__5696 (
            .O(N__23846),
            .I(N__23823));
    InMux I__5695 (
            .O(N__23845),
            .I(N__23820));
    CascadeMux I__5694 (
            .O(N__23844),
            .I(N__23813));
    CascadeMux I__5693 (
            .O(N__23843),
            .I(N__23810));
    CascadeMux I__5692 (
            .O(N__23842),
            .I(N__23807));
    CascadeMux I__5691 (
            .O(N__23841),
            .I(N__23803));
    InMux I__5690 (
            .O(N__23840),
            .I(N__23798));
    InMux I__5689 (
            .O(N__23837),
            .I(N__23798));
    InMux I__5688 (
            .O(N__23834),
            .I(N__23795));
    InMux I__5687 (
            .O(N__23833),
            .I(N__23792));
    InMux I__5686 (
            .O(N__23832),
            .I(N__23789));
    InMux I__5685 (
            .O(N__23831),
            .I(N__23784));
    InMux I__5684 (
            .O(N__23828),
            .I(N__23784));
    InMux I__5683 (
            .O(N__23827),
            .I(N__23780));
    InMux I__5682 (
            .O(N__23826),
            .I(N__23777));
    InMux I__5681 (
            .O(N__23823),
            .I(N__23774));
    LocalMux I__5680 (
            .O(N__23820),
            .I(N__23771));
    InMux I__5679 (
            .O(N__23819),
            .I(N__23768));
    InMux I__5678 (
            .O(N__23818),
            .I(N__23759));
    InMux I__5677 (
            .O(N__23817),
            .I(N__23759));
    InMux I__5676 (
            .O(N__23816),
            .I(N__23759));
    InMux I__5675 (
            .O(N__23813),
            .I(N__23759));
    InMux I__5674 (
            .O(N__23810),
            .I(N__23756));
    InMux I__5673 (
            .O(N__23807),
            .I(N__23753));
    InMux I__5672 (
            .O(N__23806),
            .I(N__23750));
    InMux I__5671 (
            .O(N__23803),
            .I(N__23747));
    LocalMux I__5670 (
            .O(N__23798),
            .I(N__23742));
    LocalMux I__5669 (
            .O(N__23795),
            .I(N__23742));
    LocalMux I__5668 (
            .O(N__23792),
            .I(N__23737));
    LocalMux I__5667 (
            .O(N__23789),
            .I(N__23737));
    LocalMux I__5666 (
            .O(N__23784),
            .I(N__23734));
    InMux I__5665 (
            .O(N__23783),
            .I(N__23730));
    LocalMux I__5664 (
            .O(N__23780),
            .I(N__23723));
    LocalMux I__5663 (
            .O(N__23777),
            .I(N__23723));
    LocalMux I__5662 (
            .O(N__23774),
            .I(N__23723));
    Span4Mux_v I__5661 (
            .O(N__23771),
            .I(N__23712));
    LocalMux I__5660 (
            .O(N__23768),
            .I(N__23712));
    LocalMux I__5659 (
            .O(N__23759),
            .I(N__23712));
    LocalMux I__5658 (
            .O(N__23756),
            .I(N__23712));
    LocalMux I__5657 (
            .O(N__23753),
            .I(N__23712));
    LocalMux I__5656 (
            .O(N__23750),
            .I(N__23707));
    LocalMux I__5655 (
            .O(N__23747),
            .I(N__23707));
    Span4Mux_h I__5654 (
            .O(N__23742),
            .I(N__23704));
    Span4Mux_v I__5653 (
            .O(N__23737),
            .I(N__23699));
    Span4Mux_h I__5652 (
            .O(N__23734),
            .I(N__23699));
    InMux I__5651 (
            .O(N__23733),
            .I(N__23696));
    LocalMux I__5650 (
            .O(N__23730),
            .I(N__23693));
    Span4Mux_v I__5649 (
            .O(N__23723),
            .I(N__23686));
    Span4Mux_h I__5648 (
            .O(N__23712),
            .I(N__23686));
    Span4Mux_v I__5647 (
            .O(N__23707),
            .I(N__23686));
    Span4Mux_h I__5646 (
            .O(N__23704),
            .I(N__23683));
    Span4Mux_h I__5645 (
            .O(N__23699),
            .I(N__23680));
    LocalMux I__5644 (
            .O(N__23696),
            .I(TX_ADDR_12));
    Odrv4 I__5643 (
            .O(N__23693),
            .I(TX_ADDR_12));
    Odrv4 I__5642 (
            .O(N__23686),
            .I(TX_ADDR_12));
    Odrv4 I__5641 (
            .O(N__23683),
            .I(TX_ADDR_12));
    Odrv4 I__5640 (
            .O(N__23680),
            .I(TX_ADDR_12));
    InMux I__5639 (
            .O(N__23669),
            .I(N__23666));
    LocalMux I__5638 (
            .O(N__23666),
            .I(N__23663));
    Span4Mux_h I__5637 (
            .O(N__23663),
            .I(N__23660));
    Odrv4 I__5636 (
            .O(N__23660),
            .I(\line_buffer.n551 ));
    InMux I__5635 (
            .O(N__23657),
            .I(N__23654));
    LocalMux I__5634 (
            .O(N__23654),
            .I(\line_buffer.n3543 ));
    InMux I__5633 (
            .O(N__23651),
            .I(N__23648));
    LocalMux I__5632 (
            .O(N__23648),
            .I(N__23645));
    Span12Mux_h I__5631 (
            .O(N__23645),
            .I(N__23642));
    Span12Mux_v I__5630 (
            .O(N__23642),
            .I(N__23639));
    Odrv12 I__5629 (
            .O(N__23639),
            .I(\line_buffer.n582 ));
    InMux I__5628 (
            .O(N__23636),
            .I(N__23633));
    LocalMux I__5627 (
            .O(N__23633),
            .I(N__23630));
    Span12Mux_h I__5626 (
            .O(N__23630),
            .I(N__23627));
    Odrv12 I__5625 (
            .O(N__23627),
            .I(\line_buffer.n590 ));
    InMux I__5624 (
            .O(N__23624),
            .I(N__23621));
    LocalMux I__5623 (
            .O(N__23621),
            .I(\line_buffer.n3480 ));
    InMux I__5622 (
            .O(N__23618),
            .I(N__23615));
    LocalMux I__5621 (
            .O(N__23615),
            .I(N__23612));
    Span4Mux_v I__5620 (
            .O(N__23612),
            .I(N__23609));
    Odrv4 I__5619 (
            .O(N__23609),
            .I(TX_DATA_3));
    IoInMux I__5618 (
            .O(N__23606),
            .I(N__23603));
    LocalMux I__5617 (
            .O(N__23603),
            .I(N__23599));
    IoInMux I__5616 (
            .O(N__23602),
            .I(N__23596));
    IoSpan4Mux I__5615 (
            .O(N__23599),
            .I(N__23593));
    LocalMux I__5614 (
            .O(N__23596),
            .I(N__23589));
    Span4Mux_s3_v I__5613 (
            .O(N__23593),
            .I(N__23586));
    IoInMux I__5612 (
            .O(N__23592),
            .I(N__23583));
    Span4Mux_s3_v I__5611 (
            .O(N__23589),
            .I(N__23580));
    Sp12to4 I__5610 (
            .O(N__23586),
            .I(N__23577));
    LocalMux I__5609 (
            .O(N__23583),
            .I(N__23574));
    Span4Mux_h I__5608 (
            .O(N__23580),
            .I(N__23571));
    Span12Mux_s11_v I__5607 (
            .O(N__23577),
            .I(N__23568));
    Span12Mux_s8_h I__5606 (
            .O(N__23574),
            .I(N__23565));
    Span4Mux_v I__5605 (
            .O(N__23571),
            .I(N__23562));
    Span12Mux_h I__5604 (
            .O(N__23568),
            .I(N__23559));
    Span12Mux_h I__5603 (
            .O(N__23565),
            .I(N__23556));
    Span4Mux_v I__5602 (
            .O(N__23562),
            .I(N__23553));
    Odrv12 I__5601 (
            .O(N__23559),
            .I(n1811));
    Odrv12 I__5600 (
            .O(N__23556),
            .I(n1811));
    Odrv4 I__5599 (
            .O(N__23553),
            .I(n1811));
    ClkMux I__5598 (
            .O(N__23546),
            .I(N__23543));
    LocalMux I__5597 (
            .O(N__23543),
            .I(N__23539));
    ClkMux I__5596 (
            .O(N__23542),
            .I(N__23536));
    Span4Mux_h I__5595 (
            .O(N__23539),
            .I(N__23530));
    LocalMux I__5594 (
            .O(N__23536),
            .I(N__23530));
    ClkMux I__5593 (
            .O(N__23535),
            .I(N__23527));
    Span4Mux_v I__5592 (
            .O(N__23530),
            .I(N__23521));
    LocalMux I__5591 (
            .O(N__23527),
            .I(N__23521));
    ClkMux I__5590 (
            .O(N__23526),
            .I(N__23518));
    Span4Mux_h I__5589 (
            .O(N__23521),
            .I(N__23511));
    LocalMux I__5588 (
            .O(N__23518),
            .I(N__23511));
    ClkMux I__5587 (
            .O(N__23517),
            .I(N__23508));
    ClkMux I__5586 (
            .O(N__23516),
            .I(N__23502));
    Span4Mux_v I__5585 (
            .O(N__23511),
            .I(N__23493));
    LocalMux I__5584 (
            .O(N__23508),
            .I(N__23493));
    ClkMux I__5583 (
            .O(N__23507),
            .I(N__23490));
    ClkMux I__5582 (
            .O(N__23506),
            .I(N__23487));
    ClkMux I__5581 (
            .O(N__23505),
            .I(N__23479));
    LocalMux I__5580 (
            .O(N__23502),
            .I(N__23476));
    ClkMux I__5579 (
            .O(N__23501),
            .I(N__23473));
    ClkMux I__5578 (
            .O(N__23500),
            .I(N__23469));
    ClkMux I__5577 (
            .O(N__23499),
            .I(N__23465));
    ClkMux I__5576 (
            .O(N__23498),
            .I(N__23460));
    Span4Mux_h I__5575 (
            .O(N__23493),
            .I(N__23450));
    LocalMux I__5574 (
            .O(N__23490),
            .I(N__23450));
    LocalMux I__5573 (
            .O(N__23487),
            .I(N__23447));
    ClkMux I__5572 (
            .O(N__23486),
            .I(N__23444));
    ClkMux I__5571 (
            .O(N__23485),
            .I(N__23441));
    ClkMux I__5570 (
            .O(N__23484),
            .I(N__23437));
    ClkMux I__5569 (
            .O(N__23483),
            .I(N__23430));
    ClkMux I__5568 (
            .O(N__23482),
            .I(N__23423));
    LocalMux I__5567 (
            .O(N__23479),
            .I(N__23419));
    Span4Mux_h I__5566 (
            .O(N__23476),
            .I(N__23414));
    LocalMux I__5565 (
            .O(N__23473),
            .I(N__23414));
    ClkMux I__5564 (
            .O(N__23472),
            .I(N__23411));
    LocalMux I__5563 (
            .O(N__23469),
            .I(N__23408));
    ClkMux I__5562 (
            .O(N__23468),
            .I(N__23405));
    LocalMux I__5561 (
            .O(N__23465),
            .I(N__23401));
    ClkMux I__5560 (
            .O(N__23464),
            .I(N__23398));
    ClkMux I__5559 (
            .O(N__23463),
            .I(N__23394));
    LocalMux I__5558 (
            .O(N__23460),
            .I(N__23386));
    ClkMux I__5557 (
            .O(N__23459),
            .I(N__23383));
    ClkMux I__5556 (
            .O(N__23458),
            .I(N__23380));
    ClkMux I__5555 (
            .O(N__23457),
            .I(N__23373));
    ClkMux I__5554 (
            .O(N__23456),
            .I(N__23368));
    ClkMux I__5553 (
            .O(N__23455),
            .I(N__23365));
    Span4Mux_h I__5552 (
            .O(N__23450),
            .I(N__23361));
    Span4Mux_h I__5551 (
            .O(N__23447),
            .I(N__23354));
    LocalMux I__5550 (
            .O(N__23444),
            .I(N__23354));
    LocalMux I__5549 (
            .O(N__23441),
            .I(N__23354));
    ClkMux I__5548 (
            .O(N__23440),
            .I(N__23351));
    LocalMux I__5547 (
            .O(N__23437),
            .I(N__23348));
    ClkMux I__5546 (
            .O(N__23436),
            .I(N__23345));
    ClkMux I__5545 (
            .O(N__23435),
            .I(N__23342));
    ClkMux I__5544 (
            .O(N__23434),
            .I(N__23339));
    ClkMux I__5543 (
            .O(N__23433),
            .I(N__23336));
    LocalMux I__5542 (
            .O(N__23430),
            .I(N__23332));
    ClkMux I__5541 (
            .O(N__23429),
            .I(N__23329));
    ClkMux I__5540 (
            .O(N__23428),
            .I(N__23325));
    ClkMux I__5539 (
            .O(N__23427),
            .I(N__23322));
    ClkMux I__5538 (
            .O(N__23426),
            .I(N__23313));
    LocalMux I__5537 (
            .O(N__23423),
            .I(N__23309));
    ClkMux I__5536 (
            .O(N__23422),
            .I(N__23306));
    Span4Mux_h I__5535 (
            .O(N__23419),
            .I(N__23295));
    Span4Mux_h I__5534 (
            .O(N__23414),
            .I(N__23295));
    LocalMux I__5533 (
            .O(N__23411),
            .I(N__23295));
    Span4Mux_h I__5532 (
            .O(N__23408),
            .I(N__23290));
    LocalMux I__5531 (
            .O(N__23405),
            .I(N__23290));
    ClkMux I__5530 (
            .O(N__23404),
            .I(N__23287));
    Span4Mux_h I__5529 (
            .O(N__23401),
            .I(N__23282));
    LocalMux I__5528 (
            .O(N__23398),
            .I(N__23282));
    ClkMux I__5527 (
            .O(N__23397),
            .I(N__23279));
    LocalMux I__5526 (
            .O(N__23394),
            .I(N__23276));
    ClkMux I__5525 (
            .O(N__23393),
            .I(N__23273));
    ClkMux I__5524 (
            .O(N__23392),
            .I(N__23270));
    ClkMux I__5523 (
            .O(N__23391),
            .I(N__23267));
    ClkMux I__5522 (
            .O(N__23390),
            .I(N__23264));
    ClkMux I__5521 (
            .O(N__23389),
            .I(N__23259));
    Span4Mux_h I__5520 (
            .O(N__23386),
            .I(N__23254));
    LocalMux I__5519 (
            .O(N__23383),
            .I(N__23254));
    LocalMux I__5518 (
            .O(N__23380),
            .I(N__23251));
    ClkMux I__5517 (
            .O(N__23379),
            .I(N__23248));
    ClkMux I__5516 (
            .O(N__23378),
            .I(N__23245));
    ClkMux I__5515 (
            .O(N__23377),
            .I(N__23242));
    ClkMux I__5514 (
            .O(N__23376),
            .I(N__23239));
    LocalMux I__5513 (
            .O(N__23373),
            .I(N__23236));
    ClkMux I__5512 (
            .O(N__23372),
            .I(N__23233));
    ClkMux I__5511 (
            .O(N__23371),
            .I(N__23230));
    LocalMux I__5510 (
            .O(N__23368),
            .I(N__23222));
    LocalMux I__5509 (
            .O(N__23365),
            .I(N__23222));
    ClkMux I__5508 (
            .O(N__23364),
            .I(N__23219));
    Span4Mux_v I__5507 (
            .O(N__23361),
            .I(N__23213));
    Span4Mux_h I__5506 (
            .O(N__23354),
            .I(N__23213));
    LocalMux I__5505 (
            .O(N__23351),
            .I(N__23206));
    Span4Mux_v I__5504 (
            .O(N__23348),
            .I(N__23206));
    LocalMux I__5503 (
            .O(N__23345),
            .I(N__23206));
    LocalMux I__5502 (
            .O(N__23342),
            .I(N__23201));
    LocalMux I__5501 (
            .O(N__23339),
            .I(N__23201));
    LocalMux I__5500 (
            .O(N__23336),
            .I(N__23198));
    ClkMux I__5499 (
            .O(N__23335),
            .I(N__23195));
    Span4Mux_h I__5498 (
            .O(N__23332),
            .I(N__23191));
    LocalMux I__5497 (
            .O(N__23329),
            .I(N__23188));
    ClkMux I__5496 (
            .O(N__23328),
            .I(N__23185));
    LocalMux I__5495 (
            .O(N__23325),
            .I(N__23179));
    LocalMux I__5494 (
            .O(N__23322),
            .I(N__23176));
    ClkMux I__5493 (
            .O(N__23321),
            .I(N__23173));
    ClkMux I__5492 (
            .O(N__23320),
            .I(N__23170));
    ClkMux I__5491 (
            .O(N__23319),
            .I(N__23166));
    ClkMux I__5490 (
            .O(N__23318),
            .I(N__23162));
    ClkMux I__5489 (
            .O(N__23317),
            .I(N__23158));
    ClkMux I__5488 (
            .O(N__23316),
            .I(N__23155));
    LocalMux I__5487 (
            .O(N__23313),
            .I(N__23151));
    ClkMux I__5486 (
            .O(N__23312),
            .I(N__23148));
    Span4Mux_h I__5485 (
            .O(N__23309),
            .I(N__23142));
    LocalMux I__5484 (
            .O(N__23306),
            .I(N__23142));
    ClkMux I__5483 (
            .O(N__23305),
            .I(N__23139));
    ClkMux I__5482 (
            .O(N__23304),
            .I(N__23136));
    ClkMux I__5481 (
            .O(N__23303),
            .I(N__23133));
    ClkMux I__5480 (
            .O(N__23302),
            .I(N__23126));
    Span4Mux_v I__5479 (
            .O(N__23295),
            .I(N__23112));
    Span4Mux_h I__5478 (
            .O(N__23290),
            .I(N__23112));
    LocalMux I__5477 (
            .O(N__23287),
            .I(N__23112));
    Span4Mux_h I__5476 (
            .O(N__23282),
            .I(N__23112));
    LocalMux I__5475 (
            .O(N__23279),
            .I(N__23112));
    Span4Mux_h I__5474 (
            .O(N__23276),
            .I(N__23105));
    LocalMux I__5473 (
            .O(N__23273),
            .I(N__23105));
    LocalMux I__5472 (
            .O(N__23270),
            .I(N__23105));
    LocalMux I__5471 (
            .O(N__23267),
            .I(N__23102));
    LocalMux I__5470 (
            .O(N__23264),
            .I(N__23099));
    ClkMux I__5469 (
            .O(N__23263),
            .I(N__23096));
    ClkMux I__5468 (
            .O(N__23262),
            .I(N__23093));
    LocalMux I__5467 (
            .O(N__23259),
            .I(N__23088));
    Span4Mux_v I__5466 (
            .O(N__23254),
            .I(N__23081));
    Span4Mux_h I__5465 (
            .O(N__23251),
            .I(N__23081));
    LocalMux I__5464 (
            .O(N__23248),
            .I(N__23081));
    LocalMux I__5463 (
            .O(N__23245),
            .I(N__23078));
    LocalMux I__5462 (
            .O(N__23242),
            .I(N__23075));
    LocalMux I__5461 (
            .O(N__23239),
            .I(N__23072));
    Span4Mux_v I__5460 (
            .O(N__23236),
            .I(N__23065));
    LocalMux I__5459 (
            .O(N__23233),
            .I(N__23065));
    LocalMux I__5458 (
            .O(N__23230),
            .I(N__23065));
    ClkMux I__5457 (
            .O(N__23229),
            .I(N__23062));
    ClkMux I__5456 (
            .O(N__23228),
            .I(N__23058));
    ClkMux I__5455 (
            .O(N__23227),
            .I(N__23054));
    Span4Mux_h I__5454 (
            .O(N__23222),
            .I(N__23049));
    LocalMux I__5453 (
            .O(N__23219),
            .I(N__23049));
    ClkMux I__5452 (
            .O(N__23218),
            .I(N__23046));
    Span4Mux_v I__5451 (
            .O(N__23213),
            .I(N__23035));
    Span4Mux_h I__5450 (
            .O(N__23206),
            .I(N__23035));
    Span4Mux_h I__5449 (
            .O(N__23201),
            .I(N__23035));
    Span4Mux_h I__5448 (
            .O(N__23198),
            .I(N__23035));
    LocalMux I__5447 (
            .O(N__23195),
            .I(N__23035));
    ClkMux I__5446 (
            .O(N__23194),
            .I(N__23032));
    Span4Mux_v I__5445 (
            .O(N__23191),
            .I(N__23026));
    Span4Mux_h I__5444 (
            .O(N__23188),
            .I(N__23026));
    LocalMux I__5443 (
            .O(N__23185),
            .I(N__23023));
    ClkMux I__5442 (
            .O(N__23184),
            .I(N__23020));
    ClkMux I__5441 (
            .O(N__23183),
            .I(N__23016));
    ClkMux I__5440 (
            .O(N__23182),
            .I(N__23012));
    Span4Mux_s2_v I__5439 (
            .O(N__23179),
            .I(N__23004));
    Span4Mux_h I__5438 (
            .O(N__23176),
            .I(N__23004));
    LocalMux I__5437 (
            .O(N__23173),
            .I(N__23004));
    LocalMux I__5436 (
            .O(N__23170),
            .I(N__23001));
    ClkMux I__5435 (
            .O(N__23169),
            .I(N__22998));
    LocalMux I__5434 (
            .O(N__23166),
            .I(N__22994));
    ClkMux I__5433 (
            .O(N__23165),
            .I(N__22991));
    LocalMux I__5432 (
            .O(N__23162),
            .I(N__22988));
    ClkMux I__5431 (
            .O(N__23161),
            .I(N__22985));
    LocalMux I__5430 (
            .O(N__23158),
            .I(N__22980));
    LocalMux I__5429 (
            .O(N__23155),
            .I(N__22980));
    ClkMux I__5428 (
            .O(N__23154),
            .I(N__22977));
    Span4Mux_h I__5427 (
            .O(N__23151),
            .I(N__22973));
    LocalMux I__5426 (
            .O(N__23148),
            .I(N__22970));
    ClkMux I__5425 (
            .O(N__23147),
            .I(N__22966));
    Span4Mux_h I__5424 (
            .O(N__23142),
            .I(N__22961));
    LocalMux I__5423 (
            .O(N__23139),
            .I(N__22961));
    LocalMux I__5422 (
            .O(N__23136),
            .I(N__22956));
    LocalMux I__5421 (
            .O(N__23133),
            .I(N__22956));
    ClkMux I__5420 (
            .O(N__23132),
            .I(N__22953));
    ClkMux I__5419 (
            .O(N__23131),
            .I(N__22950));
    ClkMux I__5418 (
            .O(N__23130),
            .I(N__22947));
    ClkMux I__5417 (
            .O(N__23129),
            .I(N__22944));
    LocalMux I__5416 (
            .O(N__23126),
            .I(N__22941));
    ClkMux I__5415 (
            .O(N__23125),
            .I(N__22938));
    ClkMux I__5414 (
            .O(N__23124),
            .I(N__22933));
    ClkMux I__5413 (
            .O(N__23123),
            .I(N__22929));
    Span4Mux_h I__5412 (
            .O(N__23112),
            .I(N__22922));
    Span4Mux_v I__5411 (
            .O(N__23105),
            .I(N__22922));
    Span4Mux_h I__5410 (
            .O(N__23102),
            .I(N__22922));
    Span4Mux_v I__5409 (
            .O(N__23099),
            .I(N__22915));
    LocalMux I__5408 (
            .O(N__23096),
            .I(N__22915));
    LocalMux I__5407 (
            .O(N__23093),
            .I(N__22915));
    ClkMux I__5406 (
            .O(N__23092),
            .I(N__22912));
    ClkMux I__5405 (
            .O(N__23091),
            .I(N__22907));
    Span4Mux_h I__5404 (
            .O(N__23088),
            .I(N__22900));
    Span4Mux_h I__5403 (
            .O(N__23081),
            .I(N__22900));
    Span4Mux_h I__5402 (
            .O(N__23078),
            .I(N__22900));
    Span4Mux_v I__5401 (
            .O(N__23075),
            .I(N__22891));
    Span4Mux_h I__5400 (
            .O(N__23072),
            .I(N__22891));
    Span4Mux_h I__5399 (
            .O(N__23065),
            .I(N__22891));
    LocalMux I__5398 (
            .O(N__23062),
            .I(N__22891));
    ClkMux I__5397 (
            .O(N__23061),
            .I(N__22888));
    LocalMux I__5396 (
            .O(N__23058),
            .I(N__22885));
    ClkMux I__5395 (
            .O(N__23057),
            .I(N__22882));
    LocalMux I__5394 (
            .O(N__23054),
            .I(N__22879));
    Span4Mux_h I__5393 (
            .O(N__23049),
            .I(N__22870));
    LocalMux I__5392 (
            .O(N__23046),
            .I(N__22870));
    Span4Mux_h I__5391 (
            .O(N__23035),
            .I(N__22870));
    LocalMux I__5390 (
            .O(N__23032),
            .I(N__22870));
    ClkMux I__5389 (
            .O(N__23031),
            .I(N__22867));
    Span4Mux_v I__5388 (
            .O(N__23026),
            .I(N__22860));
    Span4Mux_h I__5387 (
            .O(N__23023),
            .I(N__22860));
    LocalMux I__5386 (
            .O(N__23020),
            .I(N__22860));
    ClkMux I__5385 (
            .O(N__23019),
            .I(N__22857));
    LocalMux I__5384 (
            .O(N__23016),
            .I(N__22854));
    ClkMux I__5383 (
            .O(N__23015),
            .I(N__22851));
    LocalMux I__5382 (
            .O(N__23012),
            .I(N__22848));
    ClkMux I__5381 (
            .O(N__23011),
            .I(N__22845));
    Span4Mux_v I__5380 (
            .O(N__23004),
            .I(N__22837));
    Span4Mux_h I__5379 (
            .O(N__23001),
            .I(N__22837));
    LocalMux I__5378 (
            .O(N__22998),
            .I(N__22837));
    ClkMux I__5377 (
            .O(N__22997),
            .I(N__22834));
    Span4Mux_v I__5376 (
            .O(N__22994),
            .I(N__22824));
    LocalMux I__5375 (
            .O(N__22991),
            .I(N__22824));
    Span4Mux_v I__5374 (
            .O(N__22988),
            .I(N__22824));
    LocalMux I__5373 (
            .O(N__22985),
            .I(N__22824));
    Span4Mux_v I__5372 (
            .O(N__22980),
            .I(N__22819));
    LocalMux I__5371 (
            .O(N__22977),
            .I(N__22819));
    ClkMux I__5370 (
            .O(N__22976),
            .I(N__22816));
    Span4Mux_v I__5369 (
            .O(N__22973),
            .I(N__22811));
    Span4Mux_h I__5368 (
            .O(N__22970),
            .I(N__22811));
    ClkMux I__5367 (
            .O(N__22969),
            .I(N__22808));
    LocalMux I__5366 (
            .O(N__22966),
            .I(N__22805));
    Span4Mux_v I__5365 (
            .O(N__22961),
            .I(N__22796));
    Span4Mux_h I__5364 (
            .O(N__22956),
            .I(N__22796));
    LocalMux I__5363 (
            .O(N__22953),
            .I(N__22796));
    LocalMux I__5362 (
            .O(N__22950),
            .I(N__22796));
    LocalMux I__5361 (
            .O(N__22947),
            .I(N__22793));
    LocalMux I__5360 (
            .O(N__22944),
            .I(N__22786));
    Span4Mux_v I__5359 (
            .O(N__22941),
            .I(N__22786));
    LocalMux I__5358 (
            .O(N__22938),
            .I(N__22786));
    ClkMux I__5357 (
            .O(N__22937),
            .I(N__22783));
    ClkMux I__5356 (
            .O(N__22936),
            .I(N__22780));
    LocalMux I__5355 (
            .O(N__22933),
            .I(N__22776));
    ClkMux I__5354 (
            .O(N__22932),
            .I(N__22773));
    LocalMux I__5353 (
            .O(N__22929),
            .I(N__22769));
    Span4Mux_v I__5352 (
            .O(N__22922),
            .I(N__22764));
    Span4Mux_h I__5351 (
            .O(N__22915),
            .I(N__22764));
    LocalMux I__5350 (
            .O(N__22912),
            .I(N__22761));
    ClkMux I__5349 (
            .O(N__22911),
            .I(N__22758));
    IoInMux I__5348 (
            .O(N__22910),
            .I(N__22755));
    LocalMux I__5347 (
            .O(N__22907),
            .I(N__22752));
    Span4Mux_v I__5346 (
            .O(N__22900),
            .I(N__22748));
    Span4Mux_h I__5345 (
            .O(N__22891),
            .I(N__22745));
    LocalMux I__5344 (
            .O(N__22888),
            .I(N__22742));
    Span4Mux_h I__5343 (
            .O(N__22885),
            .I(N__22739));
    LocalMux I__5342 (
            .O(N__22882),
            .I(N__22736));
    Span4Mux_v I__5341 (
            .O(N__22879),
            .I(N__22729));
    Span4Mux_v I__5340 (
            .O(N__22870),
            .I(N__22729));
    LocalMux I__5339 (
            .O(N__22867),
            .I(N__22729));
    Span4Mux_h I__5338 (
            .O(N__22860),
            .I(N__22724));
    LocalMux I__5337 (
            .O(N__22857),
            .I(N__22724));
    Span4Mux_v I__5336 (
            .O(N__22854),
            .I(N__22719));
    LocalMux I__5335 (
            .O(N__22851),
            .I(N__22719));
    Span4Mux_h I__5334 (
            .O(N__22848),
            .I(N__22714));
    LocalMux I__5333 (
            .O(N__22845),
            .I(N__22714));
    ClkMux I__5332 (
            .O(N__22844),
            .I(N__22711));
    Span4Mux_v I__5331 (
            .O(N__22837),
            .I(N__22707));
    LocalMux I__5330 (
            .O(N__22834),
            .I(N__22704));
    ClkMux I__5329 (
            .O(N__22833),
            .I(N__22701));
    Span4Mux_h I__5328 (
            .O(N__22824),
            .I(N__22693));
    Span4Mux_h I__5327 (
            .O(N__22819),
            .I(N__22693));
    LocalMux I__5326 (
            .O(N__22816),
            .I(N__22693));
    Span4Mux_h I__5325 (
            .O(N__22811),
            .I(N__22688));
    LocalMux I__5324 (
            .O(N__22808),
            .I(N__22688));
    Span4Mux_h I__5323 (
            .O(N__22805),
            .I(N__22675));
    Span4Mux_h I__5322 (
            .O(N__22796),
            .I(N__22675));
    Span4Mux_v I__5321 (
            .O(N__22793),
            .I(N__22675));
    Span4Mux_h I__5320 (
            .O(N__22786),
            .I(N__22675));
    LocalMux I__5319 (
            .O(N__22783),
            .I(N__22675));
    LocalMux I__5318 (
            .O(N__22780),
            .I(N__22675));
    ClkMux I__5317 (
            .O(N__22779),
            .I(N__22672));
    Span4Mux_h I__5316 (
            .O(N__22776),
            .I(N__22669));
    LocalMux I__5315 (
            .O(N__22773),
            .I(N__22666));
    ClkMux I__5314 (
            .O(N__22772),
            .I(N__22663));
    Span4Mux_v I__5313 (
            .O(N__22769),
            .I(N__22654));
    Span4Mux_v I__5312 (
            .O(N__22764),
            .I(N__22654));
    Span4Mux_h I__5311 (
            .O(N__22761),
            .I(N__22654));
    LocalMux I__5310 (
            .O(N__22758),
            .I(N__22654));
    LocalMux I__5309 (
            .O(N__22755),
            .I(N__22651));
    Span4Mux_h I__5308 (
            .O(N__22752),
            .I(N__22648));
    ClkMux I__5307 (
            .O(N__22751),
            .I(N__22645));
    Span4Mux_v I__5306 (
            .O(N__22748),
            .I(N__22637));
    Span4Mux_v I__5305 (
            .O(N__22745),
            .I(N__22637));
    Span4Mux_h I__5304 (
            .O(N__22742),
            .I(N__22637));
    Span4Mux_v I__5303 (
            .O(N__22739),
            .I(N__22632));
    Span4Mux_h I__5302 (
            .O(N__22736),
            .I(N__22632));
    Span4Mux_v I__5301 (
            .O(N__22729),
            .I(N__22625));
    Span4Mux_h I__5300 (
            .O(N__22724),
            .I(N__22625));
    Span4Mux_h I__5299 (
            .O(N__22719),
            .I(N__22625));
    Span4Mux_v I__5298 (
            .O(N__22714),
            .I(N__22620));
    LocalMux I__5297 (
            .O(N__22711),
            .I(N__22620));
    ClkMux I__5296 (
            .O(N__22710),
            .I(N__22617));
    Sp12to4 I__5295 (
            .O(N__22707),
            .I(N__22612));
    Sp12to4 I__5294 (
            .O(N__22704),
            .I(N__22612));
    LocalMux I__5293 (
            .O(N__22701),
            .I(N__22609));
    ClkMux I__5292 (
            .O(N__22700),
            .I(N__22606));
    Span4Mux_h I__5291 (
            .O(N__22693),
            .I(N__22597));
    Span4Mux_h I__5290 (
            .O(N__22688),
            .I(N__22597));
    Span4Mux_v I__5289 (
            .O(N__22675),
            .I(N__22597));
    LocalMux I__5288 (
            .O(N__22672),
            .I(N__22597));
    Span4Mux_h I__5287 (
            .O(N__22669),
            .I(N__22590));
    Span4Mux_v I__5286 (
            .O(N__22666),
            .I(N__22590));
    LocalMux I__5285 (
            .O(N__22663),
            .I(N__22590));
    Span4Mux_h I__5284 (
            .O(N__22654),
            .I(N__22587));
    Span4Mux_s1_v I__5283 (
            .O(N__22651),
            .I(N__22584));
    Span4Mux_v I__5282 (
            .O(N__22648),
            .I(N__22579));
    LocalMux I__5281 (
            .O(N__22645),
            .I(N__22579));
    ClkMux I__5280 (
            .O(N__22644),
            .I(N__22576));
    Span4Mux_v I__5279 (
            .O(N__22637),
            .I(N__22573));
    Span4Mux_h I__5278 (
            .O(N__22632),
            .I(N__22570));
    Span4Mux_v I__5277 (
            .O(N__22625),
            .I(N__22567));
    Span4Mux_h I__5276 (
            .O(N__22620),
            .I(N__22564));
    LocalMux I__5275 (
            .O(N__22617),
            .I(N__22561));
    Span12Mux_h I__5274 (
            .O(N__22612),
            .I(N__22554));
    Span12Mux_h I__5273 (
            .O(N__22609),
            .I(N__22554));
    LocalMux I__5272 (
            .O(N__22606),
            .I(N__22554));
    Span4Mux_v I__5271 (
            .O(N__22597),
            .I(N__22549));
    Span4Mux_h I__5270 (
            .O(N__22590),
            .I(N__22549));
    Span4Mux_v I__5269 (
            .O(N__22587),
            .I(N__22546));
    Sp12to4 I__5268 (
            .O(N__22584),
            .I(N__22541));
    Sp12to4 I__5267 (
            .O(N__22579),
            .I(N__22541));
    LocalMux I__5266 (
            .O(N__22576),
            .I(N__22538));
    Span4Mux_v I__5265 (
            .O(N__22573),
            .I(N__22535));
    Span4Mux_h I__5264 (
            .O(N__22570),
            .I(N__22528));
    Span4Mux_v I__5263 (
            .O(N__22567),
            .I(N__22528));
    Span4Mux_h I__5262 (
            .O(N__22564),
            .I(N__22528));
    Span12Mux_h I__5261 (
            .O(N__22561),
            .I(N__22521));
    Span12Mux_v I__5260 (
            .O(N__22554),
            .I(N__22521));
    Sp12to4 I__5259 (
            .O(N__22549),
            .I(N__22521));
    Span4Mux_v I__5258 (
            .O(N__22546),
            .I(N__22518));
    Span12Mux_h I__5257 (
            .O(N__22541),
            .I(N__22513));
    Span12Mux_h I__5256 (
            .O(N__22538),
            .I(N__22513));
    Odrv4 I__5255 (
            .O(N__22535),
            .I(ADV_CLK_c));
    Odrv4 I__5254 (
            .O(N__22528),
            .I(ADV_CLK_c));
    Odrv12 I__5253 (
            .O(N__22521),
            .I(ADV_CLK_c));
    Odrv4 I__5252 (
            .O(N__22518),
            .I(ADV_CLK_c));
    Odrv12 I__5251 (
            .O(N__22513),
            .I(ADV_CLK_c));
    InMux I__5250 (
            .O(N__22502),
            .I(N__22499));
    LocalMux I__5249 (
            .O(N__22499),
            .I(N__22496));
    Span4Mux_v I__5248 (
            .O(N__22496),
            .I(N__22493));
    Span4Mux_h I__5247 (
            .O(N__22493),
            .I(N__22490));
    Odrv4 I__5246 (
            .O(N__22490),
            .I(\line_buffer.n517 ));
    InMux I__5245 (
            .O(N__22487),
            .I(N__22484));
    LocalMux I__5244 (
            .O(N__22484),
            .I(N__22481));
    Span12Mux_v I__5243 (
            .O(N__22481),
            .I(N__22478));
    Span12Mux_v I__5242 (
            .O(N__22478),
            .I(N__22475));
    Odrv12 I__5241 (
            .O(N__22475),
            .I(\line_buffer.n525 ));
    CascadeMux I__5240 (
            .O(N__22472),
            .I(\line_buffer.n3603_cascade_ ));
    InMux I__5239 (
            .O(N__22469),
            .I(N__22466));
    LocalMux I__5238 (
            .O(N__22466),
            .I(\line_buffer.n3606 ));
    InMux I__5237 (
            .O(N__22463),
            .I(N__22460));
    LocalMux I__5236 (
            .O(N__22460),
            .I(N__22457));
    Span4Mux_h I__5235 (
            .O(N__22457),
            .I(N__22454));
    Span4Mux_h I__5234 (
            .O(N__22454),
            .I(N__22451));
    Odrv4 I__5233 (
            .O(N__22451),
            .I(\line_buffer.n462 ));
    CascadeMux I__5232 (
            .O(N__22448),
            .I(N__22445));
    InMux I__5231 (
            .O(N__22445),
            .I(N__22442));
    LocalMux I__5230 (
            .O(N__22442),
            .I(N__22439));
    Span12Mux_h I__5229 (
            .O(N__22439),
            .I(N__22436));
    Span12Mux_v I__5228 (
            .O(N__22436),
            .I(N__22433));
    Odrv12 I__5227 (
            .O(N__22433),
            .I(\line_buffer.n454 ));
    CascadeMux I__5226 (
            .O(N__22430),
            .I(\line_buffer.n3546_cascade_ ));
    InMux I__5225 (
            .O(N__22427),
            .I(N__22424));
    LocalMux I__5224 (
            .O(N__22424),
            .I(\line_buffer.n3576 ));
    InMux I__5223 (
            .O(N__22421),
            .I(N__22418));
    LocalMux I__5222 (
            .O(N__22418),
            .I(N__22415));
    Span12Mux_v I__5221 (
            .O(N__22415),
            .I(N__22412));
    Odrv12 I__5220 (
            .O(N__22412),
            .I(\line_buffer.n555 ));
    InMux I__5219 (
            .O(N__22409),
            .I(N__22406));
    LocalMux I__5218 (
            .O(N__22406),
            .I(N__22403));
    Odrv12 I__5217 (
            .O(N__22403),
            .I(\line_buffer.n547 ));
    InMux I__5216 (
            .O(N__22400),
            .I(N__22397));
    LocalMux I__5215 (
            .O(N__22397),
            .I(N__22394));
    Span4Mux_h I__5214 (
            .O(N__22394),
            .I(N__22391));
    Span4Mux_h I__5213 (
            .O(N__22391),
            .I(N__22388));
    Odrv4 I__5212 (
            .O(N__22388),
            .I(\line_buffer.n461 ));
    InMux I__5211 (
            .O(N__22385),
            .I(N__22382));
    LocalMux I__5210 (
            .O(N__22382),
            .I(N__22379));
    Span12Mux_h I__5209 (
            .O(N__22379),
            .I(N__22376));
    Span12Mux_v I__5208 (
            .O(N__22376),
            .I(N__22373));
    Odrv12 I__5207 (
            .O(N__22373),
            .I(\line_buffer.n453 ));
    InMux I__5206 (
            .O(N__22370),
            .I(N__22367));
    LocalMux I__5205 (
            .O(N__22367),
            .I(N__22364));
    Span12Mux_h I__5204 (
            .O(N__22364),
            .I(N__22361));
    Odrv12 I__5203 (
            .O(N__22361),
            .I(\line_buffer.n588 ));
    InMux I__5202 (
            .O(N__22358),
            .I(N__22355));
    LocalMux I__5201 (
            .O(N__22355),
            .I(N__22352));
    Span12Mux_h I__5200 (
            .O(N__22352),
            .I(N__22349));
    Span12Mux_v I__5199 (
            .O(N__22349),
            .I(N__22346));
    Odrv12 I__5198 (
            .O(N__22346),
            .I(\line_buffer.n580 ));
    InMux I__5197 (
            .O(N__22343),
            .I(N__22340));
    LocalMux I__5196 (
            .O(N__22340),
            .I(N__22337));
    Odrv4 I__5195 (
            .O(N__22337),
            .I(\line_buffer.n3522 ));
    InMux I__5194 (
            .O(N__22334),
            .I(N__22331));
    LocalMux I__5193 (
            .O(N__22331),
            .I(N__22328));
    Span4Mux_h I__5192 (
            .O(N__22328),
            .I(N__22325));
    Span4Mux_h I__5191 (
            .O(N__22325),
            .I(N__22322));
    Odrv4 I__5190 (
            .O(N__22322),
            .I(\line_buffer.n458 ));
    CascadeMux I__5189 (
            .O(N__22319),
            .I(N__22316));
    InMux I__5188 (
            .O(N__22316),
            .I(N__22313));
    LocalMux I__5187 (
            .O(N__22313),
            .I(N__22310));
    Span4Mux_v I__5186 (
            .O(N__22310),
            .I(N__22307));
    Span4Mux_h I__5185 (
            .O(N__22307),
            .I(N__22304));
    Span4Mux_v I__5184 (
            .O(N__22304),
            .I(N__22301));
    Span4Mux_v I__5183 (
            .O(N__22301),
            .I(N__22298));
    Odrv4 I__5182 (
            .O(N__22298),
            .I(\line_buffer.n450 ));
    InMux I__5181 (
            .O(N__22295),
            .I(N__22292));
    LocalMux I__5180 (
            .O(N__22292),
            .I(N__22289));
    Odrv4 I__5179 (
            .O(N__22289),
            .I(\line_buffer.n3579 ));
    InMux I__5178 (
            .O(N__22286),
            .I(N__22283));
    LocalMux I__5177 (
            .O(N__22283),
            .I(\line_buffer.n3582 ));
    InMux I__5176 (
            .O(N__22280),
            .I(N__22277));
    LocalMux I__5175 (
            .O(N__22277),
            .I(N__22274));
    Span4Mux_v I__5174 (
            .O(N__22274),
            .I(N__22271));
    Odrv4 I__5173 (
            .O(N__22271),
            .I(TX_DATA_2));
    IoInMux I__5172 (
            .O(N__22268),
            .I(N__22265));
    LocalMux I__5171 (
            .O(N__22265),
            .I(N__22262));
    IoSpan4Mux I__5170 (
            .O(N__22262),
            .I(N__22259));
    IoSpan4Mux I__5169 (
            .O(N__22259),
            .I(N__22255));
    IoInMux I__5168 (
            .O(N__22258),
            .I(N__22252));
    IoSpan4Mux I__5167 (
            .O(N__22255),
            .I(N__22247));
    LocalMux I__5166 (
            .O(N__22252),
            .I(N__22247));
    IoSpan4Mux I__5165 (
            .O(N__22247),
            .I(N__22244));
    Span4Mux_s0_h I__5164 (
            .O(N__22244),
            .I(N__22240));
    IoInMux I__5163 (
            .O(N__22243),
            .I(N__22237));
    Sp12to4 I__5162 (
            .O(N__22240),
            .I(N__22234));
    LocalMux I__5161 (
            .O(N__22237),
            .I(N__22231));
    Span12Mux_s11_h I__5160 (
            .O(N__22234),
            .I(N__22228));
    Span12Mux_s11_v I__5159 (
            .O(N__22231),
            .I(N__22225));
    Odrv12 I__5158 (
            .O(N__22228),
            .I(n1812));
    Odrv12 I__5157 (
            .O(N__22225),
            .I(n1812));
    InMux I__5156 (
            .O(N__22220),
            .I(N__22217));
    LocalMux I__5155 (
            .O(N__22217),
            .I(N__22214));
    Span4Mux_v I__5154 (
            .O(N__22214),
            .I(N__22211));
    Odrv4 I__5153 (
            .O(N__22211),
            .I(TX_DATA_7));
    IoInMux I__5152 (
            .O(N__22208),
            .I(N__22204));
    IoInMux I__5151 (
            .O(N__22207),
            .I(N__22201));
    LocalMux I__5150 (
            .O(N__22204),
            .I(N__22198));
    LocalMux I__5149 (
            .O(N__22201),
            .I(N__22194));
    IoSpan4Mux I__5148 (
            .O(N__22198),
            .I(N__22191));
    IoInMux I__5147 (
            .O(N__22197),
            .I(N__22188));
    Span4Mux_s3_v I__5146 (
            .O(N__22194),
            .I(N__22185));
    Sp12to4 I__5145 (
            .O(N__22191),
            .I(N__22182));
    LocalMux I__5144 (
            .O(N__22188),
            .I(N__22179));
    Span4Mux_h I__5143 (
            .O(N__22185),
            .I(N__22176));
    Span12Mux_s6_h I__5142 (
            .O(N__22182),
            .I(N__22173));
    Span12Mux_s4_v I__5141 (
            .O(N__22179),
            .I(N__22170));
    Span4Mux_h I__5140 (
            .O(N__22176),
            .I(N__22167));
    Span12Mux_h I__5139 (
            .O(N__22173),
            .I(N__22162));
    Span12Mux_h I__5138 (
            .O(N__22170),
            .I(N__22162));
    Span4Mux_v I__5137 (
            .O(N__22167),
            .I(N__22159));
    Odrv12 I__5136 (
            .O(N__22162),
            .I(ADV_B_c));
    Odrv4 I__5135 (
            .O(N__22159),
            .I(ADV_B_c));
    InMux I__5134 (
            .O(N__22154),
            .I(N__22151));
    LocalMux I__5133 (
            .O(N__22151),
            .I(N__22145));
    InMux I__5132 (
            .O(N__22150),
            .I(N__22142));
    InMux I__5131 (
            .O(N__22149),
            .I(N__22139));
    InMux I__5130 (
            .O(N__22148),
            .I(N__22136));
    Span4Mux_v I__5129 (
            .O(N__22145),
            .I(N__22129));
    LocalMux I__5128 (
            .O(N__22142),
            .I(N__22122));
    LocalMux I__5127 (
            .O(N__22139),
            .I(N__22122));
    LocalMux I__5126 (
            .O(N__22136),
            .I(N__22122));
    InMux I__5125 (
            .O(N__22135),
            .I(N__22119));
    InMux I__5124 (
            .O(N__22134),
            .I(N__22116));
    InMux I__5123 (
            .O(N__22133),
            .I(N__22113));
    InMux I__5122 (
            .O(N__22132),
            .I(N__22110));
    Sp12to4 I__5121 (
            .O(N__22129),
            .I(N__22107));
    Span12Mux_s11_v I__5120 (
            .O(N__22122),
            .I(N__22100));
    LocalMux I__5119 (
            .O(N__22119),
            .I(N__22100));
    LocalMux I__5118 (
            .O(N__22116),
            .I(N__22100));
    LocalMux I__5117 (
            .O(N__22113),
            .I(N__22095));
    LocalMux I__5116 (
            .O(N__22110),
            .I(N__22095));
    Span12Mux_h I__5115 (
            .O(N__22107),
            .I(N__22092));
    Span12Mux_v I__5114 (
            .O(N__22100),
            .I(N__22089));
    Span4Mux_s2_v I__5113 (
            .O(N__22095),
            .I(N__22086));
    Span12Mux_v I__5112 (
            .O(N__22092),
            .I(N__22081));
    Span12Mux_h I__5111 (
            .O(N__22089),
            .I(N__22081));
    Span4Mux_h I__5110 (
            .O(N__22086),
            .I(N__22078));
    Odrv12 I__5109 (
            .O(N__22081),
            .I(RX_DATA_7));
    Odrv4 I__5108 (
            .O(N__22078),
            .I(RX_DATA_7));
    InMux I__5107 (
            .O(N__22073),
            .I(N__22070));
    LocalMux I__5106 (
            .O(N__22070),
            .I(N__22067));
    Span4Mux_v I__5105 (
            .O(N__22067),
            .I(N__22064));
    Span4Mux_v I__5104 (
            .O(N__22064),
            .I(N__22061));
    Span4Mux_h I__5103 (
            .O(N__22061),
            .I(N__22058));
    Odrv4 I__5102 (
            .O(N__22058),
            .I(\line_buffer.n465 ));
    CascadeMux I__5101 (
            .O(N__22055),
            .I(N__22052));
    InMux I__5100 (
            .O(N__22052),
            .I(N__22049));
    LocalMux I__5099 (
            .O(N__22049),
            .I(N__22046));
    Sp12to4 I__5098 (
            .O(N__22046),
            .I(N__22043));
    Span12Mux_v I__5097 (
            .O(N__22043),
            .I(N__22040));
    Odrv12 I__5096 (
            .O(N__22040),
            .I(\line_buffer.n457 ));
    InMux I__5095 (
            .O(N__22037),
            .I(N__22034));
    LocalMux I__5094 (
            .O(N__22034),
            .I(\line_buffer.n3588 ));
    InMux I__5093 (
            .O(N__22031),
            .I(N__22028));
    LocalMux I__5092 (
            .O(N__22028),
            .I(N__22025));
    Span12Mux_v I__5091 (
            .O(N__22025),
            .I(N__22022));
    Odrv12 I__5090 (
            .O(N__22022),
            .I(\line_buffer.n557 ));
    InMux I__5089 (
            .O(N__22019),
            .I(N__22016));
    LocalMux I__5088 (
            .O(N__22016),
            .I(N__22013));
    Span4Mux_h I__5087 (
            .O(N__22013),
            .I(N__22010));
    Span4Mux_h I__5086 (
            .O(N__22010),
            .I(N__22007));
    Odrv4 I__5085 (
            .O(N__22007),
            .I(\line_buffer.n549 ));
    InMux I__5084 (
            .O(N__22004),
            .I(N__22001));
    LocalMux I__5083 (
            .O(N__22001),
            .I(N__21998));
    Span4Mux_v I__5082 (
            .O(N__21998),
            .I(N__21995));
    Span4Mux_h I__5081 (
            .O(N__21995),
            .I(N__21992));
    Odrv4 I__5080 (
            .O(N__21992),
            .I(\line_buffer.n460 ));
    CascadeMux I__5079 (
            .O(N__21989),
            .I(N__21986));
    InMux I__5078 (
            .O(N__21986),
            .I(N__21983));
    LocalMux I__5077 (
            .O(N__21983),
            .I(N__21980));
    Span4Mux_v I__5076 (
            .O(N__21980),
            .I(N__21977));
    Span4Mux_v I__5075 (
            .O(N__21977),
            .I(N__21974));
    Sp12to4 I__5074 (
            .O(N__21974),
            .I(N__21971));
    Span12Mux_h I__5073 (
            .O(N__21971),
            .I(N__21968));
    Odrv12 I__5072 (
            .O(N__21968),
            .I(\line_buffer.n452 ));
    InMux I__5071 (
            .O(N__21965),
            .I(N__21962));
    LocalMux I__5070 (
            .O(N__21962),
            .I(N__21959));
    Odrv4 I__5069 (
            .O(N__21959),
            .I(\line_buffer.n3549 ));
    CascadeMux I__5068 (
            .O(N__21956),
            .I(\line_buffer.n3552_cascade_ ));
    InMux I__5067 (
            .O(N__21953),
            .I(N__21950));
    LocalMux I__5066 (
            .O(N__21950),
            .I(N__21947));
    Span12Mux_v I__5065 (
            .O(N__21947),
            .I(N__21944));
    Span12Mux_h I__5064 (
            .O(N__21944),
            .I(N__21941));
    Odrv12 I__5063 (
            .O(N__21941),
            .I(\line_buffer.n527 ));
    CascadeMux I__5062 (
            .O(N__21938),
            .I(N__21935));
    InMux I__5061 (
            .O(N__21935),
            .I(N__21932));
    LocalMux I__5060 (
            .O(N__21932),
            .I(N__21929));
    Span4Mux_v I__5059 (
            .O(N__21929),
            .I(N__21926));
    Span4Mux_h I__5058 (
            .O(N__21926),
            .I(N__21923));
    Span4Mux_v I__5057 (
            .O(N__21923),
            .I(N__21920));
    Odrv4 I__5056 (
            .O(N__21920),
            .I(\line_buffer.n519 ));
    InMux I__5055 (
            .O(N__21917),
            .I(N__21914));
    LocalMux I__5054 (
            .O(N__21914),
            .I(\line_buffer.n3573 ));
    InMux I__5053 (
            .O(N__21911),
            .I(N__21908));
    LocalMux I__5052 (
            .O(N__21908),
            .I(N__21905));
    Span4Mux_v I__5051 (
            .O(N__21905),
            .I(N__21902));
    Sp12to4 I__5050 (
            .O(N__21902),
            .I(N__21899));
    Odrv12 I__5049 (
            .O(N__21899),
            .I(\line_buffer.n589 ));
    InMux I__5048 (
            .O(N__21896),
            .I(N__21893));
    LocalMux I__5047 (
            .O(N__21893),
            .I(N__21890));
    Span4Mux_v I__5046 (
            .O(N__21890),
            .I(N__21887));
    Span4Mux_h I__5045 (
            .O(N__21887),
            .I(N__21884));
    Sp12to4 I__5044 (
            .O(N__21884),
            .I(N__21881));
    Odrv12 I__5043 (
            .O(N__21881),
            .I(\line_buffer.n581 ));
    InMux I__5042 (
            .O(N__21878),
            .I(N__21875));
    LocalMux I__5041 (
            .O(N__21875),
            .I(N__21872));
    Odrv4 I__5040 (
            .O(N__21872),
            .I(TX_DATA_6));
    IoInMux I__5039 (
            .O(N__21869),
            .I(N__21866));
    LocalMux I__5038 (
            .O(N__21866),
            .I(N__21863));
    Span4Mux_s1_h I__5037 (
            .O(N__21863),
            .I(N__21859));
    IoInMux I__5036 (
            .O(N__21862),
            .I(N__21856));
    Span4Mux_h I__5035 (
            .O(N__21859),
            .I(N__21852));
    LocalMux I__5034 (
            .O(N__21856),
            .I(N__21849));
    IoInMux I__5033 (
            .O(N__21855),
            .I(N__21846));
    Span4Mux_h I__5032 (
            .O(N__21852),
            .I(N__21843));
    IoSpan4Mux I__5031 (
            .O(N__21849),
            .I(N__21840));
    LocalMux I__5030 (
            .O(N__21846),
            .I(N__21837));
    Span4Mux_h I__5029 (
            .O(N__21843),
            .I(N__21832));
    Span4Mux_s2_v I__5028 (
            .O(N__21840),
            .I(N__21832));
    Span12Mux_s11_v I__5027 (
            .O(N__21837),
            .I(N__21829));
    Span4Mux_h I__5026 (
            .O(N__21832),
            .I(N__21826));
    Span12Mux_h I__5025 (
            .O(N__21829),
            .I(N__21823));
    Span4Mux_v I__5024 (
            .O(N__21826),
            .I(N__21820));
    Odrv12 I__5023 (
            .O(N__21823),
            .I(n1808));
    Odrv4 I__5022 (
            .O(N__21820),
            .I(n1808));
    InMux I__5021 (
            .O(N__21815),
            .I(N__21812));
    LocalMux I__5020 (
            .O(N__21812),
            .I(N__21809));
    Sp12to4 I__5019 (
            .O(N__21809),
            .I(N__21806));
    Span12Mux_v I__5018 (
            .O(N__21806),
            .I(N__21803));
    Odrv12 I__5017 (
            .O(N__21803),
            .I(\line_buffer.n528 ));
    InMux I__5016 (
            .O(N__21800),
            .I(N__21797));
    LocalMux I__5015 (
            .O(N__21797),
            .I(N__21794));
    Span4Mux_h I__5014 (
            .O(N__21794),
            .I(N__21791));
    Span4Mux_h I__5013 (
            .O(N__21791),
            .I(N__21788));
    Odrv4 I__5012 (
            .O(N__21788),
            .I(\line_buffer.n520 ));
    InMux I__5011 (
            .O(N__21785),
            .I(N__21782));
    LocalMux I__5010 (
            .O(N__21782),
            .I(N__21779));
    Odrv12 I__5009 (
            .O(N__21779),
            .I(\line_buffer.n3594 ));
    InMux I__5008 (
            .O(N__21776),
            .I(N__21773));
    LocalMux I__5007 (
            .O(N__21773),
            .I(N__21770));
    Span4Mux_v I__5006 (
            .O(N__21770),
            .I(N__21767));
    Sp12to4 I__5005 (
            .O(N__21767),
            .I(N__21764));
    Odrv12 I__5004 (
            .O(N__21764),
            .I(\line_buffer.n592 ));
    InMux I__5003 (
            .O(N__21761),
            .I(N__21758));
    LocalMux I__5002 (
            .O(N__21758),
            .I(N__21755));
    Span4Mux_v I__5001 (
            .O(N__21755),
            .I(N__21752));
    Span4Mux_v I__5000 (
            .O(N__21752),
            .I(N__21749));
    Span4Mux_v I__4999 (
            .O(N__21749),
            .I(N__21746));
    Span4Mux_h I__4998 (
            .O(N__21746),
            .I(N__21743));
    Odrv4 I__4997 (
            .O(N__21743),
            .I(\line_buffer.n584 ));
    InMux I__4996 (
            .O(N__21740),
            .I(N__21737));
    LocalMux I__4995 (
            .O(N__21737),
            .I(\line_buffer.n3489 ));
    InMux I__4994 (
            .O(N__21734),
            .I(N__21731));
    LocalMux I__4993 (
            .O(N__21731),
            .I(N__21728));
    Odrv12 I__4992 (
            .O(N__21728),
            .I(\line_buffer.n3488 ));
    InMux I__4991 (
            .O(N__21725),
            .I(N__21722));
    LocalMux I__4990 (
            .O(N__21722),
            .I(\line_buffer.n3561 ));
    InMux I__4989 (
            .O(N__21719),
            .I(N__21716));
    LocalMux I__4988 (
            .O(N__21716),
            .I(N__21713));
    Span4Mux_v I__4987 (
            .O(N__21713),
            .I(N__21710));
    Sp12to4 I__4986 (
            .O(N__21710),
            .I(N__21707));
    Odrv12 I__4985 (
            .O(N__21707),
            .I(\line_buffer.n591 ));
    InMux I__4984 (
            .O(N__21704),
            .I(N__21701));
    LocalMux I__4983 (
            .O(N__21701),
            .I(N__21698));
    Span4Mux_v I__4982 (
            .O(N__21698),
            .I(N__21695));
    Span4Mux_v I__4981 (
            .O(N__21695),
            .I(N__21692));
    Span4Mux_v I__4980 (
            .O(N__21692),
            .I(N__21689));
    Span4Mux_h I__4979 (
            .O(N__21689),
            .I(N__21686));
    Odrv4 I__4978 (
            .O(N__21686),
            .I(\line_buffer.n583 ));
    InMux I__4977 (
            .O(N__21683),
            .I(N__21680));
    LocalMux I__4976 (
            .O(N__21680),
            .I(N__21677));
    Span4Mux_h I__4975 (
            .O(N__21677),
            .I(N__21674));
    Span4Mux_h I__4974 (
            .O(N__21674),
            .I(N__21671));
    Span4Mux_h I__4973 (
            .O(N__21671),
            .I(N__21668));
    Sp12to4 I__4972 (
            .O(N__21668),
            .I(N__21665));
    Span12Mux_v I__4971 (
            .O(N__21665),
            .I(N__21662));
    Odrv12 I__4970 (
            .O(N__21662),
            .I(\line_buffer.n523 ));
    CascadeMux I__4969 (
            .O(N__21659),
            .I(N__21656));
    InMux I__4968 (
            .O(N__21656),
            .I(N__21653));
    LocalMux I__4967 (
            .O(N__21653),
            .I(N__21650));
    Span4Mux_h I__4966 (
            .O(N__21650),
            .I(N__21647));
    Span4Mux_v I__4965 (
            .O(N__21647),
            .I(N__21644));
    Span4Mux_v I__4964 (
            .O(N__21644),
            .I(N__21641));
    Odrv4 I__4963 (
            .O(N__21641),
            .I(\line_buffer.n515 ));
    InMux I__4962 (
            .O(N__21638),
            .I(N__21635));
    LocalMux I__4961 (
            .O(N__21635),
            .I(\line_buffer.n3597 ));
    CascadeMux I__4960 (
            .O(N__21632),
            .I(\line_buffer.n3600_cascade_ ));
    InMux I__4959 (
            .O(N__21629),
            .I(N__21626));
    LocalMux I__4958 (
            .O(N__21626),
            .I(TX_DATA_0));
    InMux I__4957 (
            .O(N__21623),
            .I(N__21619));
    InMux I__4956 (
            .O(N__21622),
            .I(N__21615));
    LocalMux I__4955 (
            .O(N__21619),
            .I(N__21608));
    InMux I__4954 (
            .O(N__21618),
            .I(N__21599));
    LocalMux I__4953 (
            .O(N__21615),
            .I(N__21596));
    InMux I__4952 (
            .O(N__21614),
            .I(N__21593));
    InMux I__4951 (
            .O(N__21613),
            .I(N__21586));
    InMux I__4950 (
            .O(N__21612),
            .I(N__21586));
    InMux I__4949 (
            .O(N__21611),
            .I(N__21586));
    Span4Mux_v I__4948 (
            .O(N__21608),
            .I(N__21582));
    InMux I__4947 (
            .O(N__21607),
            .I(N__21579));
    InMux I__4946 (
            .O(N__21606),
            .I(N__21572));
    InMux I__4945 (
            .O(N__21605),
            .I(N__21572));
    InMux I__4944 (
            .O(N__21604),
            .I(N__21572));
    InMux I__4943 (
            .O(N__21603),
            .I(N__21569));
    InMux I__4942 (
            .O(N__21602),
            .I(N__21566));
    LocalMux I__4941 (
            .O(N__21599),
            .I(N__21563));
    Span4Mux_h I__4940 (
            .O(N__21596),
            .I(N__21558));
    LocalMux I__4939 (
            .O(N__21593),
            .I(N__21558));
    LocalMux I__4938 (
            .O(N__21586),
            .I(N__21555));
    InMux I__4937 (
            .O(N__21585),
            .I(N__21552));
    Span4Mux_h I__4936 (
            .O(N__21582),
            .I(N__21543));
    LocalMux I__4935 (
            .O(N__21579),
            .I(N__21543));
    LocalMux I__4934 (
            .O(N__21572),
            .I(N__21543));
    LocalMux I__4933 (
            .O(N__21569),
            .I(N__21543));
    LocalMux I__4932 (
            .O(N__21566),
            .I(\transmit_module.VGA_VISIBLE ));
    Odrv12 I__4931 (
            .O(N__21563),
            .I(\transmit_module.VGA_VISIBLE ));
    Odrv4 I__4930 (
            .O(N__21558),
            .I(\transmit_module.VGA_VISIBLE ));
    Odrv4 I__4929 (
            .O(N__21555),
            .I(\transmit_module.VGA_VISIBLE ));
    LocalMux I__4928 (
            .O(N__21552),
            .I(\transmit_module.VGA_VISIBLE ));
    Odrv4 I__4927 (
            .O(N__21543),
            .I(\transmit_module.VGA_VISIBLE ));
    InMux I__4926 (
            .O(N__21530),
            .I(N__21527));
    LocalMux I__4925 (
            .O(N__21527),
            .I(N__21524));
    Odrv12 I__4924 (
            .O(N__21524),
            .I(\line_buffer.n3525 ));
    CascadeMux I__4923 (
            .O(N__21521),
            .I(\line_buffer.n3524_cascade_ ));
    InMux I__4922 (
            .O(N__21518),
            .I(N__21515));
    LocalMux I__4921 (
            .O(N__21515),
            .I(N__21512));
    Odrv12 I__4920 (
            .O(N__21512),
            .I(\line_buffer.n3521 ));
    CascadeMux I__4919 (
            .O(N__21509),
            .I(\line_buffer.n3555_cascade_ ));
    InMux I__4918 (
            .O(N__21506),
            .I(N__21503));
    LocalMux I__4917 (
            .O(N__21503),
            .I(\line_buffer.n3519 ));
    InMux I__4916 (
            .O(N__21500),
            .I(N__21497));
    LocalMux I__4915 (
            .O(N__21497),
            .I(N__21494));
    Span4Mux_h I__4914 (
            .O(N__21494),
            .I(N__21491));
    Span4Mux_h I__4913 (
            .O(N__21491),
            .I(N__21488));
    Span4Mux_h I__4912 (
            .O(N__21488),
            .I(N__21485));
    Odrv4 I__4911 (
            .O(N__21485),
            .I(\line_buffer.n561 ));
    InMux I__4910 (
            .O(N__21482),
            .I(N__21479));
    LocalMux I__4909 (
            .O(N__21479),
            .I(N__21476));
    Span4Mux_h I__4908 (
            .O(N__21476),
            .I(N__21473));
    Span4Mux_h I__4907 (
            .O(N__21473),
            .I(N__21470));
    Sp12to4 I__4906 (
            .O(N__21470),
            .I(N__21467));
    Span12Mux_v I__4905 (
            .O(N__21467),
            .I(N__21464));
    Odrv12 I__4904 (
            .O(N__21464),
            .I(\line_buffer.n553 ));
    InMux I__4903 (
            .O(N__21461),
            .I(N__21458));
    LocalMux I__4902 (
            .O(N__21458),
            .I(\line_buffer.n3498 ));
    InMux I__4901 (
            .O(N__21455),
            .I(N__21452));
    LocalMux I__4900 (
            .O(N__21452),
            .I(N__21449));
    Odrv12 I__4899 (
            .O(N__21449),
            .I(\line_buffer.n587 ));
    InMux I__4898 (
            .O(N__21446),
            .I(N__21443));
    LocalMux I__4897 (
            .O(N__21443),
            .I(N__21440));
    Span12Mux_h I__4896 (
            .O(N__21440),
            .I(N__21437));
    Span12Mux_v I__4895 (
            .O(N__21437),
            .I(N__21434));
    Odrv12 I__4894 (
            .O(N__21434),
            .I(\line_buffer.n579 ));
    IoInMux I__4893 (
            .O(N__21431),
            .I(N__21427));
    IoInMux I__4892 (
            .O(N__21430),
            .I(N__21424));
    LocalMux I__4891 (
            .O(N__21427),
            .I(N__21420));
    LocalMux I__4890 (
            .O(N__21424),
            .I(N__21417));
    IoInMux I__4889 (
            .O(N__21423),
            .I(N__21414));
    Span4Mux_s1_h I__4888 (
            .O(N__21420),
            .I(N__21411));
    IoSpan4Mux I__4887 (
            .O(N__21417),
            .I(N__21408));
    LocalMux I__4886 (
            .O(N__21414),
            .I(N__21403));
    Sp12to4 I__4885 (
            .O(N__21411),
            .I(N__21403));
    Span4Mux_s3_v I__4884 (
            .O(N__21408),
            .I(N__21400));
    Span12Mux_s11_v I__4883 (
            .O(N__21403),
            .I(N__21397));
    Sp12to4 I__4882 (
            .O(N__21400),
            .I(N__21394));
    Span12Mux_h I__4881 (
            .O(N__21397),
            .I(N__21389));
    Span12Mux_s11_v I__4880 (
            .O(N__21394),
            .I(N__21389));
    Odrv12 I__4879 (
            .O(N__21389),
            .I(n1814));
    InMux I__4878 (
            .O(N__21386),
            .I(N__21383));
    LocalMux I__4877 (
            .O(N__21383),
            .I(N__21380));
    Odrv4 I__4876 (
            .O(N__21380),
            .I(TX_DATA_1));
    IoInMux I__4875 (
            .O(N__21377),
            .I(N__21374));
    LocalMux I__4874 (
            .O(N__21374),
            .I(N__21370));
    IoInMux I__4873 (
            .O(N__21373),
            .I(N__21367));
    Span4Mux_s1_v I__4872 (
            .O(N__21370),
            .I(N__21364));
    LocalMux I__4871 (
            .O(N__21367),
            .I(N__21361));
    Span4Mux_v I__4870 (
            .O(N__21364),
            .I(N__21356));
    Span4Mux_s2_h I__4869 (
            .O(N__21361),
            .I(N__21356));
    Span4Mux_h I__4868 (
            .O(N__21356),
            .I(N__21352));
    IoInMux I__4867 (
            .O(N__21355),
            .I(N__21349));
    Span4Mux_h I__4866 (
            .O(N__21352),
            .I(N__21346));
    LocalMux I__4865 (
            .O(N__21349),
            .I(N__21343));
    Sp12to4 I__4864 (
            .O(N__21346),
            .I(N__21340));
    Span4Mux_s3_v I__4863 (
            .O(N__21343),
            .I(N__21337));
    Span12Mux_s10_v I__4862 (
            .O(N__21340),
            .I(N__21334));
    Span4Mux_v I__4861 (
            .O(N__21337),
            .I(N__21331));
    Odrv12 I__4860 (
            .O(N__21334),
            .I(n1813));
    Odrv4 I__4859 (
            .O(N__21331),
            .I(n1813));
    InMux I__4858 (
            .O(N__21326),
            .I(N__21323));
    LocalMux I__4857 (
            .O(N__21323),
            .I(N__21320));
    Odrv12 I__4856 (
            .O(N__21320),
            .I(TX_DATA_5));
    IoInMux I__4855 (
            .O(N__21317),
            .I(N__21314));
    LocalMux I__4854 (
            .O(N__21314),
            .I(N__21311));
    Span4Mux_s0_h I__4853 (
            .O(N__21311),
            .I(N__21307));
    IoInMux I__4852 (
            .O(N__21310),
            .I(N__21304));
    Span4Mux_h I__4851 (
            .O(N__21307),
            .I(N__21300));
    LocalMux I__4850 (
            .O(N__21304),
            .I(N__21297));
    IoInMux I__4849 (
            .O(N__21303),
            .I(N__21294));
    Span4Mux_v I__4848 (
            .O(N__21300),
            .I(N__21289));
    Span4Mux_s3_v I__4847 (
            .O(N__21297),
            .I(N__21289));
    LocalMux I__4846 (
            .O(N__21294),
            .I(N__21286));
    Sp12to4 I__4845 (
            .O(N__21289),
            .I(N__21283));
    Span12Mux_s9_v I__4844 (
            .O(N__21286),
            .I(N__21280));
    Span12Mux_h I__4843 (
            .O(N__21283),
            .I(N__21277));
    Odrv12 I__4842 (
            .O(N__21280),
            .I(n1809));
    Odrv12 I__4841 (
            .O(N__21277),
            .I(n1809));
    InMux I__4840 (
            .O(N__21272),
            .I(N__21269));
    LocalMux I__4839 (
            .O(N__21269),
            .I(N__21266));
    Span4Mux_h I__4838 (
            .O(N__21266),
            .I(N__21263));
    Span4Mux_h I__4837 (
            .O(N__21263),
            .I(N__21260));
    Odrv4 I__4836 (
            .O(N__21260),
            .I(\line_buffer.n464 ));
    InMux I__4835 (
            .O(N__21257),
            .I(N__21254));
    LocalMux I__4834 (
            .O(N__21254),
            .I(N__21251));
    Span4Mux_v I__4833 (
            .O(N__21251),
            .I(N__21248));
    Span4Mux_h I__4832 (
            .O(N__21248),
            .I(N__21245));
    Span4Mux_h I__4831 (
            .O(N__21245),
            .I(N__21242));
    Odrv4 I__4830 (
            .O(N__21242),
            .I(\line_buffer.n456 ));
    InMux I__4829 (
            .O(N__21239),
            .I(N__21236));
    LocalMux I__4828 (
            .O(N__21236),
            .I(\line_buffer.n3497 ));
    InMux I__4827 (
            .O(N__21233),
            .I(N__21230));
    LocalMux I__4826 (
            .O(N__21230),
            .I(N__21227));
    Span4Mux_v I__4825 (
            .O(N__21227),
            .I(N__21224));
    Span4Mux_v I__4824 (
            .O(N__21224),
            .I(N__21221));
    Sp12to4 I__4823 (
            .O(N__21221),
            .I(N__21218));
    Odrv12 I__4822 (
            .O(N__21218),
            .I(\line_buffer.n524 ));
    InMux I__4821 (
            .O(N__21215),
            .I(N__21212));
    LocalMux I__4820 (
            .O(N__21212),
            .I(N__21209));
    Odrv12 I__4819 (
            .O(N__21209),
            .I(\line_buffer.n516 ));
    InMux I__4818 (
            .O(N__21206),
            .I(N__21203));
    LocalMux I__4817 (
            .O(N__21203),
            .I(N__21200));
    Span4Mux_v I__4816 (
            .O(N__21200),
            .I(N__21197));
    Span4Mux_v I__4815 (
            .O(N__21197),
            .I(N__21194));
    Sp12to4 I__4814 (
            .O(N__21194),
            .I(N__21191));
    Odrv12 I__4813 (
            .O(N__21191),
            .I(\line_buffer.n560 ));
    InMux I__4812 (
            .O(N__21188),
            .I(N__21185));
    LocalMux I__4811 (
            .O(N__21185),
            .I(N__21182));
    Odrv12 I__4810 (
            .O(N__21182),
            .I(\line_buffer.n552 ));
    InMux I__4809 (
            .O(N__21179),
            .I(N__21176));
    LocalMux I__4808 (
            .O(N__21176),
            .I(N__21173));
    Span4Mux_v I__4807 (
            .O(N__21173),
            .I(N__21170));
    Odrv4 I__4806 (
            .O(N__21170),
            .I(\transmit_module.X_DELTA_PATTERN_1 ));
    InMux I__4805 (
            .O(N__21167),
            .I(N__21164));
    LocalMux I__4804 (
            .O(N__21164),
            .I(\transmit_module.X_DELTA_PATTERN_2 ));
    InMux I__4803 (
            .O(N__21161),
            .I(N__21158));
    LocalMux I__4802 (
            .O(N__21158),
            .I(\transmit_module.X_DELTA_PATTERN_3 ));
    InMux I__4801 (
            .O(N__21155),
            .I(N__21152));
    LocalMux I__4800 (
            .O(N__21152),
            .I(\transmit_module.X_DELTA_PATTERN_5 ));
    InMux I__4799 (
            .O(N__21149),
            .I(N__21146));
    LocalMux I__4798 (
            .O(N__21146),
            .I(\transmit_module.X_DELTA_PATTERN_4 ));
    InMux I__4797 (
            .O(N__21143),
            .I(N__21140));
    LocalMux I__4796 (
            .O(N__21140),
            .I(\transmit_module.X_DELTA_PATTERN_7 ));
    InMux I__4795 (
            .O(N__21137),
            .I(N__21134));
    LocalMux I__4794 (
            .O(N__21134),
            .I(\transmit_module.X_DELTA_PATTERN_6 ));
    CEMux I__4793 (
            .O(N__21131),
            .I(N__21126));
    CEMux I__4792 (
            .O(N__21130),
            .I(N__21123));
    CEMux I__4791 (
            .O(N__21129),
            .I(N__21120));
    LocalMux I__4790 (
            .O(N__21126),
            .I(N__21112));
    LocalMux I__4789 (
            .O(N__21123),
            .I(N__21112));
    LocalMux I__4788 (
            .O(N__21120),
            .I(N__21108));
    CEMux I__4787 (
            .O(N__21119),
            .I(N__21105));
    CEMux I__4786 (
            .O(N__21118),
            .I(N__21102));
    CEMux I__4785 (
            .O(N__21117),
            .I(N__21099));
    Span4Mux_v I__4784 (
            .O(N__21112),
            .I(N__21096));
    CEMux I__4783 (
            .O(N__21111),
            .I(N__21093));
    Span4Mux_h I__4782 (
            .O(N__21108),
            .I(N__21086));
    LocalMux I__4781 (
            .O(N__21105),
            .I(N__21086));
    LocalMux I__4780 (
            .O(N__21102),
            .I(N__21086));
    LocalMux I__4779 (
            .O(N__21099),
            .I(N__21083));
    Span4Mux_h I__4778 (
            .O(N__21096),
            .I(N__21080));
    LocalMux I__4777 (
            .O(N__21093),
            .I(N__21077));
    Span4Mux_v I__4776 (
            .O(N__21086),
            .I(N__21074));
    Odrv4 I__4775 (
            .O(N__21083),
            .I(\transmit_module.n2115 ));
    Odrv4 I__4774 (
            .O(N__21080),
            .I(\transmit_module.n2115 ));
    Odrv4 I__4773 (
            .O(N__21077),
            .I(\transmit_module.n2115 ));
    Odrv4 I__4772 (
            .O(N__21074),
            .I(\transmit_module.n2115 ));
    SRMux I__4771 (
            .O(N__21065),
            .I(N__21058));
    SRMux I__4770 (
            .O(N__21064),
            .I(N__21051));
    SRMux I__4769 (
            .O(N__21063),
            .I(N__21048));
    CEMux I__4768 (
            .O(N__21062),
            .I(N__21043));
    CEMux I__4767 (
            .O(N__21061),
            .I(N__21040));
    LocalMux I__4766 (
            .O(N__21058),
            .I(N__21037));
    SRMux I__4765 (
            .O(N__21057),
            .I(N__21034));
    CEMux I__4764 (
            .O(N__21056),
            .I(N__21029));
    SRMux I__4763 (
            .O(N__21055),
            .I(N__21026));
    SRMux I__4762 (
            .O(N__21054),
            .I(N__21023));
    LocalMux I__4761 (
            .O(N__21051),
            .I(N__21019));
    LocalMux I__4760 (
            .O(N__21048),
            .I(N__21016));
    CEMux I__4759 (
            .O(N__21047),
            .I(N__21013));
    CEMux I__4758 (
            .O(N__21046),
            .I(N__21010));
    LocalMux I__4757 (
            .O(N__21043),
            .I(N__21006));
    LocalMux I__4756 (
            .O(N__21040),
            .I(N__21003));
    Span4Mux_h I__4755 (
            .O(N__21037),
            .I(N__21000));
    LocalMux I__4754 (
            .O(N__21034),
            .I(N__20997));
    CEMux I__4753 (
            .O(N__21033),
            .I(N__20994));
    CEMux I__4752 (
            .O(N__21032),
            .I(N__20991));
    LocalMux I__4751 (
            .O(N__21029),
            .I(N__20987));
    LocalMux I__4750 (
            .O(N__21026),
            .I(N__20984));
    LocalMux I__4749 (
            .O(N__21023),
            .I(N__20981));
    CEMux I__4748 (
            .O(N__21022),
            .I(N__20978));
    Span4Mux_h I__4747 (
            .O(N__21019),
            .I(N__20973));
    Span4Mux_h I__4746 (
            .O(N__21016),
            .I(N__20973));
    LocalMux I__4745 (
            .O(N__21013),
            .I(N__20968));
    LocalMux I__4744 (
            .O(N__21010),
            .I(N__20968));
    CEMux I__4743 (
            .O(N__21009),
            .I(N__20965));
    Span4Mux_h I__4742 (
            .O(N__21006),
            .I(N__20956));
    Span4Mux_v I__4741 (
            .O(N__21003),
            .I(N__20956));
    Span4Mux_v I__4740 (
            .O(N__21000),
            .I(N__20956));
    Span4Mux_h I__4739 (
            .O(N__20997),
            .I(N__20956));
    LocalMux I__4738 (
            .O(N__20994),
            .I(N__20953));
    LocalMux I__4737 (
            .O(N__20991),
            .I(N__20950));
    CEMux I__4736 (
            .O(N__20990),
            .I(N__20947));
    Span4Mux_v I__4735 (
            .O(N__20987),
            .I(N__20940));
    Span4Mux_h I__4734 (
            .O(N__20984),
            .I(N__20940));
    Span4Mux_h I__4733 (
            .O(N__20981),
            .I(N__20940));
    LocalMux I__4732 (
            .O(N__20978),
            .I(N__20937));
    Span4Mux_h I__4731 (
            .O(N__20973),
            .I(N__20934));
    Span4Mux_h I__4730 (
            .O(N__20968),
            .I(N__20927));
    LocalMux I__4729 (
            .O(N__20965),
            .I(N__20927));
    Span4Mux_h I__4728 (
            .O(N__20956),
            .I(N__20927));
    Span4Mux_v I__4727 (
            .O(N__20953),
            .I(N__20918));
    Span4Mux_h I__4726 (
            .O(N__20950),
            .I(N__20918));
    LocalMux I__4725 (
            .O(N__20947),
            .I(N__20918));
    Span4Mux_h I__4724 (
            .O(N__20940),
            .I(N__20918));
    Odrv12 I__4723 (
            .O(N__20937),
            .I(\transmit_module.n3635 ));
    Odrv4 I__4722 (
            .O(N__20934),
            .I(\transmit_module.n3635 ));
    Odrv4 I__4721 (
            .O(N__20927),
            .I(\transmit_module.n3635 ));
    Odrv4 I__4720 (
            .O(N__20918),
            .I(\transmit_module.n3635 ));
    InMux I__4719 (
            .O(N__20909),
            .I(N__20906));
    LocalMux I__4718 (
            .O(N__20906),
            .I(N__20903));
    Span4Mux_h I__4717 (
            .O(N__20903),
            .I(N__20900));
    Span4Mux_h I__4716 (
            .O(N__20900),
            .I(N__20897));
    Odrv4 I__4715 (
            .O(N__20897),
            .I(\line_buffer.n463 ));
    InMux I__4714 (
            .O(N__20894),
            .I(N__20891));
    LocalMux I__4713 (
            .O(N__20891),
            .I(N__20888));
    Span12Mux_h I__4712 (
            .O(N__20888),
            .I(N__20885));
    Span12Mux_v I__4711 (
            .O(N__20885),
            .I(N__20882));
    Odrv12 I__4710 (
            .O(N__20882),
            .I(\line_buffer.n455 ));
    CascadeMux I__4709 (
            .O(N__20879),
            .I(N__20872));
    InMux I__4708 (
            .O(N__20878),
            .I(N__20865));
    InMux I__4707 (
            .O(N__20877),
            .I(N__20862));
    InMux I__4706 (
            .O(N__20876),
            .I(N__20859));
    CascadeMux I__4705 (
            .O(N__20875),
            .I(N__20856));
    InMux I__4704 (
            .O(N__20872),
            .I(N__20850));
    InMux I__4703 (
            .O(N__20871),
            .I(N__20850));
    InMux I__4702 (
            .O(N__20870),
            .I(N__20845));
    InMux I__4701 (
            .O(N__20869),
            .I(N__20845));
    InMux I__4700 (
            .O(N__20868),
            .I(N__20842));
    LocalMux I__4699 (
            .O(N__20865),
            .I(N__20836));
    LocalMux I__4698 (
            .O(N__20862),
            .I(N__20833));
    LocalMux I__4697 (
            .O(N__20859),
            .I(N__20830));
    InMux I__4696 (
            .O(N__20856),
            .I(N__20825));
    InMux I__4695 (
            .O(N__20855),
            .I(N__20825));
    LocalMux I__4694 (
            .O(N__20850),
            .I(N__20812));
    LocalMux I__4693 (
            .O(N__20845),
            .I(N__20812));
    LocalMux I__4692 (
            .O(N__20842),
            .I(N__20809));
    InMux I__4691 (
            .O(N__20841),
            .I(N__20806));
    InMux I__4690 (
            .O(N__20840),
            .I(N__20801));
    InMux I__4689 (
            .O(N__20839),
            .I(N__20801));
    Span4Mux_s3_v I__4688 (
            .O(N__20836),
            .I(N__20798));
    Span4Mux_h I__4687 (
            .O(N__20833),
            .I(N__20793));
    Span4Mux_h I__4686 (
            .O(N__20830),
            .I(N__20793));
    LocalMux I__4685 (
            .O(N__20825),
            .I(N__20790));
    InMux I__4684 (
            .O(N__20824),
            .I(N__20787));
    InMux I__4683 (
            .O(N__20823),
            .I(N__20782));
    InMux I__4682 (
            .O(N__20822),
            .I(N__20782));
    InMux I__4681 (
            .O(N__20821),
            .I(N__20773));
    InMux I__4680 (
            .O(N__20820),
            .I(N__20773));
    InMux I__4679 (
            .O(N__20819),
            .I(N__20773));
    InMux I__4678 (
            .O(N__20818),
            .I(N__20773));
    CascadeMux I__4677 (
            .O(N__20817),
            .I(N__20766));
    Span4Mux_h I__4676 (
            .O(N__20812),
            .I(N__20756));
    Span4Mux_v I__4675 (
            .O(N__20809),
            .I(N__20756));
    LocalMux I__4674 (
            .O(N__20806),
            .I(N__20756));
    LocalMux I__4673 (
            .O(N__20801),
            .I(N__20753));
    Sp12to4 I__4672 (
            .O(N__20798),
            .I(N__20748));
    Sp12to4 I__4671 (
            .O(N__20793),
            .I(N__20748));
    Span4Mux_h I__4670 (
            .O(N__20790),
            .I(N__20743));
    LocalMux I__4669 (
            .O(N__20787),
            .I(N__20743));
    LocalMux I__4668 (
            .O(N__20782),
            .I(N__20738));
    LocalMux I__4667 (
            .O(N__20773),
            .I(N__20738));
    InMux I__4666 (
            .O(N__20772),
            .I(N__20731));
    InMux I__4665 (
            .O(N__20771),
            .I(N__20731));
    InMux I__4664 (
            .O(N__20770),
            .I(N__20731));
    InMux I__4663 (
            .O(N__20769),
            .I(N__20728));
    InMux I__4662 (
            .O(N__20766),
            .I(N__20725));
    InMux I__4661 (
            .O(N__20765),
            .I(N__20720));
    InMux I__4660 (
            .O(N__20764),
            .I(N__20720));
    InMux I__4659 (
            .O(N__20763),
            .I(N__20717));
    Span4Mux_v I__4658 (
            .O(N__20756),
            .I(N__20712));
    Span4Mux_v I__4657 (
            .O(N__20753),
            .I(N__20712));
    Span12Mux_v I__4656 (
            .O(N__20748),
            .I(N__20709));
    Span4Mux_v I__4655 (
            .O(N__20743),
            .I(N__20704));
    Span4Mux_v I__4654 (
            .O(N__20738),
            .I(N__20704));
    LocalMux I__4653 (
            .O(N__20731),
            .I(\transmit_module.n3627 ));
    LocalMux I__4652 (
            .O(N__20728),
            .I(\transmit_module.n3627 ));
    LocalMux I__4651 (
            .O(N__20725),
            .I(\transmit_module.n3627 ));
    LocalMux I__4650 (
            .O(N__20720),
            .I(\transmit_module.n3627 ));
    LocalMux I__4649 (
            .O(N__20717),
            .I(\transmit_module.n3627 ));
    Odrv4 I__4648 (
            .O(N__20712),
            .I(\transmit_module.n3627 ));
    Odrv12 I__4647 (
            .O(N__20709),
            .I(\transmit_module.n3627 ));
    Odrv4 I__4646 (
            .O(N__20704),
            .I(\transmit_module.n3627 ));
    InMux I__4645 (
            .O(N__20687),
            .I(N__20684));
    LocalMux I__4644 (
            .O(N__20684),
            .I(N__20681));
    Span4Mux_v I__4643 (
            .O(N__20681),
            .I(N__20678));
    Span4Mux_h I__4642 (
            .O(N__20678),
            .I(N__20675));
    Span4Mux_h I__4641 (
            .O(N__20675),
            .I(N__20672));
    Odrv4 I__4640 (
            .O(N__20672),
            .I(\line_buffer.n556 ));
    InMux I__4639 (
            .O(N__20669),
            .I(N__20666));
    LocalMux I__4638 (
            .O(N__20666),
            .I(N__20663));
    Span12Mux_v I__4637 (
            .O(N__20663),
            .I(N__20660));
    Odrv12 I__4636 (
            .O(N__20660),
            .I(\line_buffer.n548 ));
    InMux I__4635 (
            .O(N__20657),
            .I(N__20649));
    InMux I__4634 (
            .O(N__20656),
            .I(N__20646));
    InMux I__4633 (
            .O(N__20655),
            .I(N__20643));
    InMux I__4632 (
            .O(N__20654),
            .I(N__20636));
    InMux I__4631 (
            .O(N__20653),
            .I(N__20636));
    InMux I__4630 (
            .O(N__20652),
            .I(N__20636));
    LocalMux I__4629 (
            .O(N__20649),
            .I(N__20631));
    LocalMux I__4628 (
            .O(N__20646),
            .I(N__20628));
    LocalMux I__4627 (
            .O(N__20643),
            .I(N__20625));
    LocalMux I__4626 (
            .O(N__20636),
            .I(N__20622));
    InMux I__4625 (
            .O(N__20635),
            .I(N__20617));
    InMux I__4624 (
            .O(N__20634),
            .I(N__20614));
    Span12Mux_h I__4623 (
            .O(N__20631),
            .I(N__20607));
    Span4Mux_h I__4622 (
            .O(N__20628),
            .I(N__20604));
    Span12Mux_h I__4621 (
            .O(N__20625),
            .I(N__20601));
    Span4Mux_v I__4620 (
            .O(N__20622),
            .I(N__20598));
    InMux I__4619 (
            .O(N__20621),
            .I(N__20595));
    InMux I__4618 (
            .O(N__20620),
            .I(N__20592));
    LocalMux I__4617 (
            .O(N__20617),
            .I(N__20587));
    LocalMux I__4616 (
            .O(N__20614),
            .I(N__20587));
    InMux I__4615 (
            .O(N__20613),
            .I(N__20584));
    InMux I__4614 (
            .O(N__20612),
            .I(N__20577));
    InMux I__4613 (
            .O(N__20611),
            .I(N__20577));
    InMux I__4612 (
            .O(N__20610),
            .I(N__20577));
    Odrv12 I__4611 (
            .O(N__20607),
            .I(\transmit_module.Y_DELTA_PATTERN_0 ));
    Odrv4 I__4610 (
            .O(N__20604),
            .I(\transmit_module.Y_DELTA_PATTERN_0 ));
    Odrv12 I__4609 (
            .O(N__20601),
            .I(\transmit_module.Y_DELTA_PATTERN_0 ));
    Odrv4 I__4608 (
            .O(N__20598),
            .I(\transmit_module.Y_DELTA_PATTERN_0 ));
    LocalMux I__4607 (
            .O(N__20595),
            .I(\transmit_module.Y_DELTA_PATTERN_0 ));
    LocalMux I__4606 (
            .O(N__20592),
            .I(\transmit_module.Y_DELTA_PATTERN_0 ));
    Odrv4 I__4605 (
            .O(N__20587),
            .I(\transmit_module.Y_DELTA_PATTERN_0 ));
    LocalMux I__4604 (
            .O(N__20584),
            .I(\transmit_module.Y_DELTA_PATTERN_0 ));
    LocalMux I__4603 (
            .O(N__20577),
            .I(\transmit_module.Y_DELTA_PATTERN_0 ));
    CascadeMux I__4602 (
            .O(N__20558),
            .I(N__20554));
    InMux I__4601 (
            .O(N__20557),
            .I(N__20551));
    InMux I__4600 (
            .O(N__20554),
            .I(N__20548));
    LocalMux I__4599 (
            .O(N__20551),
            .I(N__20545));
    LocalMux I__4598 (
            .O(N__20548),
            .I(N__20542));
    Span12Mux_h I__4597 (
            .O(N__20545),
            .I(N__20539));
    Span4Mux_h I__4596 (
            .O(N__20542),
            .I(N__20536));
    Span12Mux_v I__4595 (
            .O(N__20539),
            .I(N__20533));
    Odrv4 I__4594 (
            .O(N__20536),
            .I(\transmit_module.n112 ));
    Odrv12 I__4593 (
            .O(N__20533),
            .I(\transmit_module.n112 ));
    InMux I__4592 (
            .O(N__20528),
            .I(N__20525));
    LocalMux I__4591 (
            .O(N__20525),
            .I(N__20520));
    InMux I__4590 (
            .O(N__20524),
            .I(N__20517));
    CascadeMux I__4589 (
            .O(N__20523),
            .I(N__20513));
    Span4Mux_v I__4588 (
            .O(N__20520),
            .I(N__20508));
    LocalMux I__4587 (
            .O(N__20517),
            .I(N__20508));
    InMux I__4586 (
            .O(N__20516),
            .I(N__20505));
    InMux I__4585 (
            .O(N__20513),
            .I(N__20502));
    Span4Mux_v I__4584 (
            .O(N__20508),
            .I(N__20499));
    LocalMux I__4583 (
            .O(N__20505),
            .I(N__20496));
    LocalMux I__4582 (
            .O(N__20502),
            .I(N__20493));
    Odrv4 I__4581 (
            .O(N__20499),
            .I(\transmit_module.TX_ADDR_4 ));
    Odrv12 I__4580 (
            .O(N__20496),
            .I(\transmit_module.TX_ADDR_4 ));
    Odrv4 I__4579 (
            .O(N__20493),
            .I(\transmit_module.TX_ADDR_4 ));
    InMux I__4578 (
            .O(N__20486),
            .I(N__20483));
    LocalMux I__4577 (
            .O(N__20483),
            .I(\transmit_module.ADDR_Y_COMPONENT_4 ));
    CEMux I__4576 (
            .O(N__20480),
            .I(N__20476));
    CEMux I__4575 (
            .O(N__20479),
            .I(N__20473));
    LocalMux I__4574 (
            .O(N__20476),
            .I(N__20469));
    LocalMux I__4573 (
            .O(N__20473),
            .I(N__20466));
    CEMux I__4572 (
            .O(N__20472),
            .I(N__20463));
    Span4Mux_h I__4571 (
            .O(N__20469),
            .I(N__20456));
    Span4Mux_h I__4570 (
            .O(N__20466),
            .I(N__20456));
    LocalMux I__4569 (
            .O(N__20463),
            .I(N__20456));
    Span4Mux_v I__4568 (
            .O(N__20456),
            .I(N__20451));
    CEMux I__4567 (
            .O(N__20455),
            .I(N__20448));
    CEMux I__4566 (
            .O(N__20454),
            .I(N__20445));
    Span4Mux_h I__4565 (
            .O(N__20451),
            .I(N__20439));
    LocalMux I__4564 (
            .O(N__20448),
            .I(N__20439));
    LocalMux I__4563 (
            .O(N__20445),
            .I(N__20436));
    CEMux I__4562 (
            .O(N__20444),
            .I(N__20433));
    Span4Mux_v I__4561 (
            .O(N__20439),
            .I(N__20430));
    Span12Mux_v I__4560 (
            .O(N__20436),
            .I(N__20425));
    LocalMux I__4559 (
            .O(N__20433),
            .I(N__20425));
    Odrv4 I__4558 (
            .O(N__20430),
            .I(\transmit_module.n2069 ));
    Odrv12 I__4557 (
            .O(N__20425),
            .I(\transmit_module.n2069 ));
    IoInMux I__4556 (
            .O(N__20420),
            .I(N__20417));
    LocalMux I__4555 (
            .O(N__20417),
            .I(N__20410));
    SRMux I__4554 (
            .O(N__20416),
            .I(N__20404));
    SRMux I__4553 (
            .O(N__20415),
            .I(N__20401));
    SRMux I__4552 (
            .O(N__20414),
            .I(N__20398));
    SRMux I__4551 (
            .O(N__20413),
            .I(N__20394));
    Span4Mux_s1_h I__4550 (
            .O(N__20410),
            .I(N__20389));
    SRMux I__4549 (
            .O(N__20409),
            .I(N__20386));
    CascadeMux I__4548 (
            .O(N__20408),
            .I(N__20381));
    CascadeMux I__4547 (
            .O(N__20407),
            .I(N__20378));
    LocalMux I__4546 (
            .O(N__20404),
            .I(N__20375));
    LocalMux I__4545 (
            .O(N__20401),
            .I(N__20372));
    LocalMux I__4544 (
            .O(N__20398),
            .I(N__20369));
    SRMux I__4543 (
            .O(N__20397),
            .I(N__20366));
    LocalMux I__4542 (
            .O(N__20394),
            .I(N__20363));
    SRMux I__4541 (
            .O(N__20393),
            .I(N__20360));
    SRMux I__4540 (
            .O(N__20392),
            .I(N__20357));
    Span4Mux_h I__4539 (
            .O(N__20389),
            .I(N__20349));
    LocalMux I__4538 (
            .O(N__20386),
            .I(N__20346));
    SRMux I__4537 (
            .O(N__20385),
            .I(N__20343));
    SRMux I__4536 (
            .O(N__20384),
            .I(N__20340));
    InMux I__4535 (
            .O(N__20381),
            .I(N__20332));
    InMux I__4534 (
            .O(N__20378),
            .I(N__20329));
    Span4Mux_h I__4533 (
            .O(N__20375),
            .I(N__20321));
    Span4Mux_v I__4532 (
            .O(N__20372),
            .I(N__20321));
    Span4Mux_h I__4531 (
            .O(N__20369),
            .I(N__20316));
    LocalMux I__4530 (
            .O(N__20366),
            .I(N__20316));
    Span4Mux_v I__4529 (
            .O(N__20363),
            .I(N__20309));
    LocalMux I__4528 (
            .O(N__20360),
            .I(N__20309));
    LocalMux I__4527 (
            .O(N__20357),
            .I(N__20309));
    SRMux I__4526 (
            .O(N__20356),
            .I(N__20306));
    CascadeMux I__4525 (
            .O(N__20355),
            .I(N__20302));
    SRMux I__4524 (
            .O(N__20354),
            .I(N__20299));
    CascadeMux I__4523 (
            .O(N__20353),
            .I(N__20289));
    SRMux I__4522 (
            .O(N__20352),
            .I(N__20281));
    Span4Mux_v I__4521 (
            .O(N__20349),
            .I(N__20272));
    Span4Mux_v I__4520 (
            .O(N__20346),
            .I(N__20272));
    LocalMux I__4519 (
            .O(N__20343),
            .I(N__20272));
    LocalMux I__4518 (
            .O(N__20340),
            .I(N__20272));
    SRMux I__4517 (
            .O(N__20339),
            .I(N__20269));
    SRMux I__4516 (
            .O(N__20338),
            .I(N__20264));
    SRMux I__4515 (
            .O(N__20337),
            .I(N__20261));
    SRMux I__4514 (
            .O(N__20336),
            .I(N__20255));
    SRMux I__4513 (
            .O(N__20335),
            .I(N__20252));
    LocalMux I__4512 (
            .O(N__20332),
            .I(N__20247));
    LocalMux I__4511 (
            .O(N__20329),
            .I(N__20244));
    CascadeMux I__4510 (
            .O(N__20328),
            .I(N__20241));
    SRMux I__4509 (
            .O(N__20327),
            .I(N__20233));
    CascadeMux I__4508 (
            .O(N__20326),
            .I(N__20230));
    Span4Mux_v I__4507 (
            .O(N__20321),
            .I(N__20220));
    Span4Mux_h I__4506 (
            .O(N__20316),
            .I(N__20220));
    Span4Mux_h I__4505 (
            .O(N__20309),
            .I(N__20220));
    LocalMux I__4504 (
            .O(N__20306),
            .I(N__20220));
    InMux I__4503 (
            .O(N__20305),
            .I(N__20217));
    InMux I__4502 (
            .O(N__20302),
            .I(N__20214));
    LocalMux I__4501 (
            .O(N__20299),
            .I(N__20211));
    SRMux I__4500 (
            .O(N__20298),
            .I(N__20208));
    SRMux I__4499 (
            .O(N__20297),
            .I(N__20205));
    SRMux I__4498 (
            .O(N__20296),
            .I(N__20202));
    SRMux I__4497 (
            .O(N__20295),
            .I(N__20199));
    SRMux I__4496 (
            .O(N__20294),
            .I(N__20196));
    SRMux I__4495 (
            .O(N__20293),
            .I(N__20193));
    SRMux I__4494 (
            .O(N__20292),
            .I(N__20190));
    InMux I__4493 (
            .O(N__20289),
            .I(N__20183));
    CascadeMux I__4492 (
            .O(N__20288),
            .I(N__20180));
    CascadeMux I__4491 (
            .O(N__20287),
            .I(N__20176));
    CascadeMux I__4490 (
            .O(N__20286),
            .I(N__20173));
    SRMux I__4489 (
            .O(N__20285),
            .I(N__20165));
    SRMux I__4488 (
            .O(N__20284),
            .I(N__20160));
    LocalMux I__4487 (
            .O(N__20281),
            .I(N__20157));
    Span4Mux_h I__4486 (
            .O(N__20272),
            .I(N__20152));
    LocalMux I__4485 (
            .O(N__20269),
            .I(N__20152));
    SRMux I__4484 (
            .O(N__20268),
            .I(N__20149));
    SRMux I__4483 (
            .O(N__20267),
            .I(N__20146));
    LocalMux I__4482 (
            .O(N__20264),
            .I(N__20141));
    LocalMux I__4481 (
            .O(N__20261),
            .I(N__20141));
    SRMux I__4480 (
            .O(N__20260),
            .I(N__20138));
    InMux I__4479 (
            .O(N__20259),
            .I(N__20135));
    CascadeMux I__4478 (
            .O(N__20258),
            .I(N__20132));
    LocalMux I__4477 (
            .O(N__20255),
            .I(N__20127));
    LocalMux I__4476 (
            .O(N__20252),
            .I(N__20127));
    SRMux I__4475 (
            .O(N__20251),
            .I(N__20124));
    SRMux I__4474 (
            .O(N__20250),
            .I(N__20118));
    Span4Mux_h I__4473 (
            .O(N__20247),
            .I(N__20113));
    Span4Mux_h I__4472 (
            .O(N__20244),
            .I(N__20113));
    InMux I__4471 (
            .O(N__20241),
            .I(N__20110));
    SRMux I__4470 (
            .O(N__20240),
            .I(N__20107));
    SRMux I__4469 (
            .O(N__20239),
            .I(N__20104));
    SRMux I__4468 (
            .O(N__20238),
            .I(N__20101));
    InMux I__4467 (
            .O(N__20237),
            .I(N__20096));
    InMux I__4466 (
            .O(N__20236),
            .I(N__20096));
    LocalMux I__4465 (
            .O(N__20233),
            .I(N__20093));
    InMux I__4464 (
            .O(N__20230),
            .I(N__20090));
    InMux I__4463 (
            .O(N__20229),
            .I(N__20087));
    Span4Mux_h I__4462 (
            .O(N__20220),
            .I(N__20080));
    LocalMux I__4461 (
            .O(N__20217),
            .I(N__20080));
    LocalMux I__4460 (
            .O(N__20214),
            .I(N__20080));
    Span4Mux_v I__4459 (
            .O(N__20211),
            .I(N__20075));
    LocalMux I__4458 (
            .O(N__20208),
            .I(N__20075));
    LocalMux I__4457 (
            .O(N__20205),
            .I(N__20070));
    LocalMux I__4456 (
            .O(N__20202),
            .I(N__20070));
    LocalMux I__4455 (
            .O(N__20199),
            .I(N__20061));
    LocalMux I__4454 (
            .O(N__20196),
            .I(N__20061));
    LocalMux I__4453 (
            .O(N__20193),
            .I(N__20061));
    LocalMux I__4452 (
            .O(N__20190),
            .I(N__20061));
    InMux I__4451 (
            .O(N__20189),
            .I(N__20058));
    CascadeMux I__4450 (
            .O(N__20188),
            .I(N__20055));
    CascadeMux I__4449 (
            .O(N__20187),
            .I(N__20052));
    SRMux I__4448 (
            .O(N__20186),
            .I(N__20049));
    LocalMux I__4447 (
            .O(N__20183),
            .I(N__20046));
    InMux I__4446 (
            .O(N__20180),
            .I(N__20043));
    InMux I__4445 (
            .O(N__20179),
            .I(N__20038));
    InMux I__4444 (
            .O(N__20176),
            .I(N__20038));
    InMux I__4443 (
            .O(N__20173),
            .I(N__20029));
    InMux I__4442 (
            .O(N__20172),
            .I(N__20029));
    InMux I__4441 (
            .O(N__20171),
            .I(N__20029));
    InMux I__4440 (
            .O(N__20170),
            .I(N__20029));
    SRMux I__4439 (
            .O(N__20169),
            .I(N__20026));
    SRMux I__4438 (
            .O(N__20168),
            .I(N__20023));
    LocalMux I__4437 (
            .O(N__20165),
            .I(N__20020));
    SRMux I__4436 (
            .O(N__20164),
            .I(N__20017));
    CascadeMux I__4435 (
            .O(N__20163),
            .I(N__20012));
    LocalMux I__4434 (
            .O(N__20160),
            .I(N__20007));
    Span4Mux_h I__4433 (
            .O(N__20157),
            .I(N__20007));
    Span4Mux_h I__4432 (
            .O(N__20152),
            .I(N__20002));
    LocalMux I__4431 (
            .O(N__20149),
            .I(N__20002));
    LocalMux I__4430 (
            .O(N__20146),
            .I(N__19995));
    Span4Mux_v I__4429 (
            .O(N__20141),
            .I(N__19995));
    LocalMux I__4428 (
            .O(N__20138),
            .I(N__19995));
    LocalMux I__4427 (
            .O(N__20135),
            .I(N__19992));
    InMux I__4426 (
            .O(N__20132),
            .I(N__19989));
    Span4Mux_v I__4425 (
            .O(N__20127),
            .I(N__19984));
    LocalMux I__4424 (
            .O(N__20124),
            .I(N__19984));
    InMux I__4423 (
            .O(N__20123),
            .I(N__19981));
    CascadeMux I__4422 (
            .O(N__20122),
            .I(N__19978));
    CascadeMux I__4421 (
            .O(N__20121),
            .I(N__19975));
    LocalMux I__4420 (
            .O(N__20118),
            .I(N__19972));
    Span4Mux_v I__4419 (
            .O(N__20113),
            .I(N__19969));
    LocalMux I__4418 (
            .O(N__20110),
            .I(N__19966));
    LocalMux I__4417 (
            .O(N__20107),
            .I(N__19963));
    LocalMux I__4416 (
            .O(N__20104),
            .I(N__19956));
    LocalMux I__4415 (
            .O(N__20101),
            .I(N__19956));
    LocalMux I__4414 (
            .O(N__20096),
            .I(N__19956));
    Span4Mux_v I__4413 (
            .O(N__20093),
            .I(N__19951));
    LocalMux I__4412 (
            .O(N__20090),
            .I(N__19951));
    LocalMux I__4411 (
            .O(N__20087),
            .I(N__19946));
    Span4Mux_v I__4410 (
            .O(N__20080),
            .I(N__19946));
    Span4Mux_h I__4409 (
            .O(N__20075),
            .I(N__19939));
    Span4Mux_v I__4408 (
            .O(N__20070),
            .I(N__19939));
    Span4Mux_v I__4407 (
            .O(N__20061),
            .I(N__19939));
    LocalMux I__4406 (
            .O(N__20058),
            .I(N__19936));
    InMux I__4405 (
            .O(N__20055),
            .I(N__19931));
    InMux I__4404 (
            .O(N__20052),
            .I(N__19931));
    LocalMux I__4403 (
            .O(N__20049),
            .I(N__19920));
    Span4Mux_h I__4402 (
            .O(N__20046),
            .I(N__19920));
    LocalMux I__4401 (
            .O(N__20043),
            .I(N__19920));
    LocalMux I__4400 (
            .O(N__20038),
            .I(N__19920));
    LocalMux I__4399 (
            .O(N__20029),
            .I(N__19920));
    LocalMux I__4398 (
            .O(N__20026),
            .I(N__19915));
    LocalMux I__4397 (
            .O(N__20023),
            .I(N__19915));
    Span4Mux_h I__4396 (
            .O(N__20020),
            .I(N__19910));
    LocalMux I__4395 (
            .O(N__20017),
            .I(N__19910));
    InMux I__4394 (
            .O(N__20016),
            .I(N__19907));
    InMux I__4393 (
            .O(N__20015),
            .I(N__19902));
    InMux I__4392 (
            .O(N__20012),
            .I(N__19902));
    Span4Mux_h I__4391 (
            .O(N__20007),
            .I(N__19895));
    Span4Mux_h I__4390 (
            .O(N__20002),
            .I(N__19895));
    Span4Mux_h I__4389 (
            .O(N__19995),
            .I(N__19895));
    Span4Mux_h I__4388 (
            .O(N__19992),
            .I(N__19890));
    LocalMux I__4387 (
            .O(N__19989),
            .I(N__19890));
    Span4Mux_h I__4386 (
            .O(N__19984),
            .I(N__19885));
    LocalMux I__4385 (
            .O(N__19981),
            .I(N__19885));
    InMux I__4384 (
            .O(N__19978),
            .I(N__19882));
    InMux I__4383 (
            .O(N__19975),
            .I(N__19879));
    Span12Mux_h I__4382 (
            .O(N__19972),
            .I(N__19872));
    Sp12to4 I__4381 (
            .O(N__19969),
            .I(N__19872));
    Span12Mux_s4_v I__4380 (
            .O(N__19966),
            .I(N__19872));
    Span4Mux_v I__4379 (
            .O(N__19963),
            .I(N__19863));
    Span4Mux_v I__4378 (
            .O(N__19956),
            .I(N__19863));
    Span4Mux_h I__4377 (
            .O(N__19951),
            .I(N__19863));
    Span4Mux_h I__4376 (
            .O(N__19946),
            .I(N__19863));
    Span4Mux_h I__4375 (
            .O(N__19939),
            .I(N__19854));
    Span4Mux_v I__4374 (
            .O(N__19936),
            .I(N__19854));
    LocalMux I__4373 (
            .O(N__19931),
            .I(N__19854));
    Span4Mux_v I__4372 (
            .O(N__19920),
            .I(N__19854));
    Span4Mux_h I__4371 (
            .O(N__19915),
            .I(N__19845));
    Span4Mux_h I__4370 (
            .O(N__19910),
            .I(N__19845));
    LocalMux I__4369 (
            .O(N__19907),
            .I(N__19845));
    LocalMux I__4368 (
            .O(N__19902),
            .I(N__19845));
    Odrv4 I__4367 (
            .O(N__19895),
            .I(ADV_VSYNC_c));
    Odrv4 I__4366 (
            .O(N__19890),
            .I(ADV_VSYNC_c));
    Odrv4 I__4365 (
            .O(N__19885),
            .I(ADV_VSYNC_c));
    LocalMux I__4364 (
            .O(N__19882),
            .I(ADV_VSYNC_c));
    LocalMux I__4363 (
            .O(N__19879),
            .I(ADV_VSYNC_c));
    Odrv12 I__4362 (
            .O(N__19872),
            .I(ADV_VSYNC_c));
    Odrv4 I__4361 (
            .O(N__19863),
            .I(ADV_VSYNC_c));
    Odrv4 I__4360 (
            .O(N__19854),
            .I(ADV_VSYNC_c));
    Odrv4 I__4359 (
            .O(N__19845),
            .I(ADV_VSYNC_c));
    InMux I__4358 (
            .O(N__19826),
            .I(N__19823));
    LocalMux I__4357 (
            .O(N__19823),
            .I(N__19820));
    Span4Mux_v I__4356 (
            .O(N__19820),
            .I(N__19817));
    Sp12to4 I__4355 (
            .O(N__19817),
            .I(N__19814));
    Odrv12 I__4354 (
            .O(N__19814),
            .I(\line_buffer.n529 ));
    InMux I__4353 (
            .O(N__19811),
            .I(N__19808));
    LocalMux I__4352 (
            .O(N__19808),
            .I(N__19805));
    Span12Mux_v I__4351 (
            .O(N__19805),
            .I(N__19802));
    Span12Mux_v I__4350 (
            .O(N__19802),
            .I(N__19799));
    Odrv12 I__4349 (
            .O(N__19799),
            .I(\line_buffer.n521 ));
    CascadeMux I__4348 (
            .O(N__19796),
            .I(\line_buffer.n3500_cascade_ ));
    InMux I__4347 (
            .O(N__19793),
            .I(N__19790));
    LocalMux I__4346 (
            .O(N__19790),
            .I(N__19787));
    Span4Mux_h I__4345 (
            .O(N__19787),
            .I(N__19784));
    Odrv4 I__4344 (
            .O(N__19784),
            .I(\line_buffer.n3501 ));
    CascadeMux I__4343 (
            .O(N__19781),
            .I(\line_buffer.n3537_cascade_ ));
    InMux I__4342 (
            .O(N__19778),
            .I(N__19774));
    InMux I__4341 (
            .O(N__19777),
            .I(N__19771));
    LocalMux I__4340 (
            .O(N__19774),
            .I(N__19767));
    LocalMux I__4339 (
            .O(N__19771),
            .I(N__19762));
    InMux I__4338 (
            .O(N__19770),
            .I(N__19759));
    Span4Mux_s1_v I__4337 (
            .O(N__19767),
            .I(N__19756));
    InMux I__4336 (
            .O(N__19766),
            .I(N__19752));
    InMux I__4335 (
            .O(N__19765),
            .I(N__19749));
    Span4Mux_v I__4334 (
            .O(N__19762),
            .I(N__19743));
    LocalMux I__4333 (
            .O(N__19759),
            .I(N__19743));
    Span4Mux_h I__4332 (
            .O(N__19756),
            .I(N__19739));
    InMux I__4331 (
            .O(N__19755),
            .I(N__19736));
    LocalMux I__4330 (
            .O(N__19752),
            .I(N__19733));
    LocalMux I__4329 (
            .O(N__19749),
            .I(N__19730));
    InMux I__4328 (
            .O(N__19748),
            .I(N__19727));
    Span4Mux_v I__4327 (
            .O(N__19743),
            .I(N__19724));
    InMux I__4326 (
            .O(N__19742),
            .I(N__19721));
    Span4Mux_h I__4325 (
            .O(N__19739),
            .I(N__19718));
    LocalMux I__4324 (
            .O(N__19736),
            .I(N__19715));
    Span4Mux_v I__4323 (
            .O(N__19733),
            .I(N__19712));
    Span4Mux_v I__4322 (
            .O(N__19730),
            .I(N__19707));
    LocalMux I__4321 (
            .O(N__19727),
            .I(N__19707));
    Span4Mux_v I__4320 (
            .O(N__19724),
            .I(N__19702));
    LocalMux I__4319 (
            .O(N__19721),
            .I(N__19702));
    Sp12to4 I__4318 (
            .O(N__19718),
            .I(N__19697));
    Span12Mux_h I__4317 (
            .O(N__19715),
            .I(N__19697));
    Span4Mux_v I__4316 (
            .O(N__19712),
            .I(N__19692));
    Span4Mux_v I__4315 (
            .O(N__19707),
            .I(N__19692));
    Span4Mux_h I__4314 (
            .O(N__19702),
            .I(N__19689));
    Span12Mux_v I__4313 (
            .O(N__19697),
            .I(N__19686));
    Sp12to4 I__4312 (
            .O(N__19692),
            .I(N__19683));
    Span4Mux_h I__4311 (
            .O(N__19689),
            .I(N__19680));
    Odrv12 I__4310 (
            .O(N__19686),
            .I(RX_DATA_2));
    Odrv12 I__4309 (
            .O(N__19683),
            .I(RX_DATA_2));
    Odrv4 I__4308 (
            .O(N__19680),
            .I(RX_DATA_2));
    CascadeMux I__4307 (
            .O(N__19673),
            .I(N__19669));
    InMux I__4306 (
            .O(N__19672),
            .I(N__19666));
    InMux I__4305 (
            .O(N__19669),
            .I(N__19663));
    LocalMux I__4304 (
            .O(N__19666),
            .I(\transmit_module.X_DELTA_PATTERN_0 ));
    LocalMux I__4303 (
            .O(N__19663),
            .I(\transmit_module.X_DELTA_PATTERN_0 ));
    InMux I__4302 (
            .O(N__19658),
            .I(N__19655));
    LocalMux I__4301 (
            .O(N__19655),
            .I(\transmit_module.X_DELTA_PATTERN_10 ));
    InMux I__4300 (
            .O(N__19652),
            .I(N__19649));
    LocalMux I__4299 (
            .O(N__19649),
            .I(\transmit_module.X_DELTA_PATTERN_15 ));
    InMux I__4298 (
            .O(N__19646),
            .I(N__19643));
    LocalMux I__4297 (
            .O(N__19643),
            .I(\transmit_module.X_DELTA_PATTERN_14 ));
    InMux I__4296 (
            .O(N__19640),
            .I(N__19637));
    LocalMux I__4295 (
            .O(N__19637),
            .I(\transmit_module.X_DELTA_PATTERN_13 ));
    InMux I__4294 (
            .O(N__19634),
            .I(N__19631));
    LocalMux I__4293 (
            .O(N__19631),
            .I(\transmit_module.X_DELTA_PATTERN_12 ));
    InMux I__4292 (
            .O(N__19628),
            .I(N__19625));
    LocalMux I__4291 (
            .O(N__19625),
            .I(\transmit_module.X_DELTA_PATTERN_11 ));
    InMux I__4290 (
            .O(N__19622),
            .I(N__19619));
    LocalMux I__4289 (
            .O(N__19619),
            .I(\transmit_module.X_DELTA_PATTERN_9 ));
    InMux I__4288 (
            .O(N__19616),
            .I(N__19613));
    LocalMux I__4287 (
            .O(N__19613),
            .I(\transmit_module.X_DELTA_PATTERN_8 ));
    InMux I__4286 (
            .O(N__19610),
            .I(N__19607));
    LocalMux I__4285 (
            .O(N__19607),
            .I(N__19604));
    Odrv12 I__4284 (
            .O(N__19604),
            .I(\transmit_module.Y_DELTA_PATTERN_1 ));
    CascadeMux I__4283 (
            .O(N__19601),
            .I(N__19598));
    InMux I__4282 (
            .O(N__19598),
            .I(N__19595));
    LocalMux I__4281 (
            .O(N__19595),
            .I(N__19592));
    Span4Mux_h I__4280 (
            .O(N__19592),
            .I(N__19588));
    InMux I__4279 (
            .O(N__19591),
            .I(N__19585));
    Odrv4 I__4278 (
            .O(N__19588),
            .I(\transmit_module.n108 ));
    LocalMux I__4277 (
            .O(N__19585),
            .I(\transmit_module.n108 ));
    InMux I__4276 (
            .O(N__19580),
            .I(N__19577));
    LocalMux I__4275 (
            .O(N__19577),
            .I(N__19573));
    InMux I__4274 (
            .O(N__19576),
            .I(N__19570));
    Odrv4 I__4273 (
            .O(N__19573),
            .I(\transmit_module.n139 ));
    LocalMux I__4272 (
            .O(N__19570),
            .I(\transmit_module.n139 ));
    CascadeMux I__4271 (
            .O(N__19565),
            .I(N__19561));
    CascadeMux I__4270 (
            .O(N__19564),
            .I(N__19558));
    CascadeBuf I__4269 (
            .O(N__19561),
            .I(N__19555));
    CascadeBuf I__4268 (
            .O(N__19558),
            .I(N__19552));
    CascadeMux I__4267 (
            .O(N__19555),
            .I(N__19549));
    CascadeMux I__4266 (
            .O(N__19552),
            .I(N__19546));
    CascadeBuf I__4265 (
            .O(N__19549),
            .I(N__19543));
    CascadeBuf I__4264 (
            .O(N__19546),
            .I(N__19540));
    CascadeMux I__4263 (
            .O(N__19543),
            .I(N__19537));
    CascadeMux I__4262 (
            .O(N__19540),
            .I(N__19534));
    CascadeBuf I__4261 (
            .O(N__19537),
            .I(N__19531));
    CascadeBuf I__4260 (
            .O(N__19534),
            .I(N__19528));
    CascadeMux I__4259 (
            .O(N__19531),
            .I(N__19525));
    CascadeMux I__4258 (
            .O(N__19528),
            .I(N__19522));
    CascadeBuf I__4257 (
            .O(N__19525),
            .I(N__19519));
    CascadeBuf I__4256 (
            .O(N__19522),
            .I(N__19516));
    CascadeMux I__4255 (
            .O(N__19519),
            .I(N__19513));
    CascadeMux I__4254 (
            .O(N__19516),
            .I(N__19510));
    CascadeBuf I__4253 (
            .O(N__19513),
            .I(N__19507));
    CascadeBuf I__4252 (
            .O(N__19510),
            .I(N__19504));
    CascadeMux I__4251 (
            .O(N__19507),
            .I(N__19501));
    CascadeMux I__4250 (
            .O(N__19504),
            .I(N__19498));
    CascadeBuf I__4249 (
            .O(N__19501),
            .I(N__19495));
    CascadeBuf I__4248 (
            .O(N__19498),
            .I(N__19492));
    CascadeMux I__4247 (
            .O(N__19495),
            .I(N__19489));
    CascadeMux I__4246 (
            .O(N__19492),
            .I(N__19486));
    CascadeBuf I__4245 (
            .O(N__19489),
            .I(N__19483));
    CascadeBuf I__4244 (
            .O(N__19486),
            .I(N__19480));
    CascadeMux I__4243 (
            .O(N__19483),
            .I(N__19477));
    CascadeMux I__4242 (
            .O(N__19480),
            .I(N__19474));
    CascadeBuf I__4241 (
            .O(N__19477),
            .I(N__19471));
    CascadeBuf I__4240 (
            .O(N__19474),
            .I(N__19468));
    CascadeMux I__4239 (
            .O(N__19471),
            .I(N__19465));
    CascadeMux I__4238 (
            .O(N__19468),
            .I(N__19462));
    CascadeBuf I__4237 (
            .O(N__19465),
            .I(N__19459));
    CascadeBuf I__4236 (
            .O(N__19462),
            .I(N__19456));
    CascadeMux I__4235 (
            .O(N__19459),
            .I(N__19453));
    CascadeMux I__4234 (
            .O(N__19456),
            .I(N__19450));
    CascadeBuf I__4233 (
            .O(N__19453),
            .I(N__19447));
    CascadeBuf I__4232 (
            .O(N__19450),
            .I(N__19444));
    CascadeMux I__4231 (
            .O(N__19447),
            .I(N__19441));
    CascadeMux I__4230 (
            .O(N__19444),
            .I(N__19438));
    CascadeBuf I__4229 (
            .O(N__19441),
            .I(N__19435));
    CascadeBuf I__4228 (
            .O(N__19438),
            .I(N__19432));
    CascadeMux I__4227 (
            .O(N__19435),
            .I(N__19429));
    CascadeMux I__4226 (
            .O(N__19432),
            .I(N__19426));
    CascadeBuf I__4225 (
            .O(N__19429),
            .I(N__19423));
    CascadeBuf I__4224 (
            .O(N__19426),
            .I(N__19420));
    CascadeMux I__4223 (
            .O(N__19423),
            .I(N__19417));
    CascadeMux I__4222 (
            .O(N__19420),
            .I(N__19414));
    CascadeBuf I__4221 (
            .O(N__19417),
            .I(N__19411));
    CascadeBuf I__4220 (
            .O(N__19414),
            .I(N__19408));
    CascadeMux I__4219 (
            .O(N__19411),
            .I(N__19405));
    CascadeMux I__4218 (
            .O(N__19408),
            .I(N__19402));
    CascadeBuf I__4217 (
            .O(N__19405),
            .I(N__19399));
    CascadeBuf I__4216 (
            .O(N__19402),
            .I(N__19396));
    CascadeMux I__4215 (
            .O(N__19399),
            .I(N__19393));
    CascadeMux I__4214 (
            .O(N__19396),
            .I(N__19390));
    CascadeBuf I__4213 (
            .O(N__19393),
            .I(N__19387));
    CascadeBuf I__4212 (
            .O(N__19390),
            .I(N__19384));
    CascadeMux I__4211 (
            .O(N__19387),
            .I(N__19381));
    CascadeMux I__4210 (
            .O(N__19384),
            .I(N__19378));
    InMux I__4209 (
            .O(N__19381),
            .I(N__19375));
    InMux I__4208 (
            .O(N__19378),
            .I(N__19372));
    LocalMux I__4207 (
            .O(N__19375),
            .I(N__19369));
    LocalMux I__4206 (
            .O(N__19372),
            .I(N__19366));
    Span4Mux_h I__4205 (
            .O(N__19369),
            .I(N__19363));
    Span4Mux_v I__4204 (
            .O(N__19366),
            .I(N__19360));
    Span4Mux_h I__4203 (
            .O(N__19363),
            .I(N__19357));
    Sp12to4 I__4202 (
            .O(N__19360),
            .I(N__19354));
    Sp12to4 I__4201 (
            .O(N__19357),
            .I(N__19351));
    Span12Mux_h I__4200 (
            .O(N__19354),
            .I(N__19346));
    Span12Mux_s5_v I__4199 (
            .O(N__19351),
            .I(N__19346));
    Odrv12 I__4198 (
            .O(N__19346),
            .I(n20));
    InMux I__4197 (
            .O(N__19343),
            .I(N__19340));
    LocalMux I__4196 (
            .O(N__19340),
            .I(N__19337));
    Odrv4 I__4195 (
            .O(N__19337),
            .I(\transmit_module.ADDR_Y_COMPONENT_7 ));
    InMux I__4194 (
            .O(N__19334),
            .I(N__19329));
    InMux I__4193 (
            .O(N__19333),
            .I(N__19325));
    InMux I__4192 (
            .O(N__19332),
            .I(N__19322));
    LocalMux I__4191 (
            .O(N__19329),
            .I(N__19319));
    CascadeMux I__4190 (
            .O(N__19328),
            .I(N__19316));
    LocalMux I__4189 (
            .O(N__19325),
            .I(N__19311));
    LocalMux I__4188 (
            .O(N__19322),
            .I(N__19311));
    Span4Mux_v I__4187 (
            .O(N__19319),
            .I(N__19308));
    InMux I__4186 (
            .O(N__19316),
            .I(N__19305));
    Odrv12 I__4185 (
            .O(N__19311),
            .I(\transmit_module.TX_ADDR_7 ));
    Odrv4 I__4184 (
            .O(N__19308),
            .I(\transmit_module.TX_ADDR_7 ));
    LocalMux I__4183 (
            .O(N__19305),
            .I(\transmit_module.TX_ADDR_7 ));
    InMux I__4182 (
            .O(N__19298),
            .I(N__19295));
    LocalMux I__4181 (
            .O(N__19295),
            .I(N__19291));
    InMux I__4180 (
            .O(N__19294),
            .I(N__19288));
    Odrv12 I__4179 (
            .O(N__19291),
            .I(\transmit_module.n109 ));
    LocalMux I__4178 (
            .O(N__19288),
            .I(\transmit_module.n109 ));
    InMux I__4177 (
            .O(N__19283),
            .I(N__19280));
    LocalMux I__4176 (
            .O(N__19280),
            .I(\transmit_module.ADDR_Y_COMPONENT_6 ));
    InMux I__4175 (
            .O(N__19277),
            .I(N__19274));
    LocalMux I__4174 (
            .O(N__19274),
            .I(N__19269));
    InMux I__4173 (
            .O(N__19273),
            .I(N__19266));
    InMux I__4172 (
            .O(N__19272),
            .I(N__19263));
    Span4Mux_v I__4171 (
            .O(N__19269),
            .I(N__19255));
    LocalMux I__4170 (
            .O(N__19266),
            .I(N__19255));
    LocalMux I__4169 (
            .O(N__19263),
            .I(N__19255));
    CascadeMux I__4168 (
            .O(N__19262),
            .I(N__19252));
    Span4Mux_v I__4167 (
            .O(N__19255),
            .I(N__19249));
    InMux I__4166 (
            .O(N__19252),
            .I(N__19246));
    Odrv4 I__4165 (
            .O(N__19249),
            .I(\transmit_module.TX_ADDR_6 ));
    LocalMux I__4164 (
            .O(N__19246),
            .I(\transmit_module.TX_ADDR_6 ));
    InMux I__4163 (
            .O(N__19241),
            .I(N__19238));
    LocalMux I__4162 (
            .O(N__19238),
            .I(N__19234));
    InMux I__4161 (
            .O(N__19237),
            .I(N__19231));
    Odrv12 I__4160 (
            .O(N__19234),
            .I(\transmit_module.n110 ));
    LocalMux I__4159 (
            .O(N__19231),
            .I(\transmit_module.n110 ));
    InMux I__4158 (
            .O(N__19226),
            .I(N__19223));
    LocalMux I__4157 (
            .O(N__19223),
            .I(N__19220));
    Odrv4 I__4156 (
            .O(N__19220),
            .I(\transmit_module.ADDR_Y_COMPONENT_2 ));
    InMux I__4155 (
            .O(N__19217),
            .I(N__19212));
    InMux I__4154 (
            .O(N__19216),
            .I(N__19209));
    CascadeMux I__4153 (
            .O(N__19215),
            .I(N__19205));
    LocalMux I__4152 (
            .O(N__19212),
            .I(N__19200));
    LocalMux I__4151 (
            .O(N__19209),
            .I(N__19200));
    InMux I__4150 (
            .O(N__19208),
            .I(N__19197));
    InMux I__4149 (
            .O(N__19205),
            .I(N__19194));
    Odrv12 I__4148 (
            .O(N__19200),
            .I(\transmit_module.TX_ADDR_2 ));
    LocalMux I__4147 (
            .O(N__19197),
            .I(\transmit_module.TX_ADDR_2 ));
    LocalMux I__4146 (
            .O(N__19194),
            .I(\transmit_module.TX_ADDR_2 ));
    InMux I__4145 (
            .O(N__19187),
            .I(N__19184));
    LocalMux I__4144 (
            .O(N__19184),
            .I(N__19181));
    Odrv4 I__4143 (
            .O(N__19181),
            .I(\transmit_module.ADDR_Y_COMPONENT_9 ));
    InMux I__4142 (
            .O(N__19178),
            .I(N__19174));
    InMux I__4141 (
            .O(N__19177),
            .I(N__19171));
    LocalMux I__4140 (
            .O(N__19174),
            .I(N__19164));
    LocalMux I__4139 (
            .O(N__19171),
            .I(N__19164));
    InMux I__4138 (
            .O(N__19170),
            .I(N__19161));
    CascadeMux I__4137 (
            .O(N__19169),
            .I(N__19158));
    Span4Mux_v I__4136 (
            .O(N__19164),
            .I(N__19155));
    LocalMux I__4135 (
            .O(N__19161),
            .I(N__19152));
    InMux I__4134 (
            .O(N__19158),
            .I(N__19149));
    Odrv4 I__4133 (
            .O(N__19155),
            .I(\transmit_module.TX_ADDR_9 ));
    Odrv12 I__4132 (
            .O(N__19152),
            .I(\transmit_module.TX_ADDR_9 ));
    LocalMux I__4131 (
            .O(N__19149),
            .I(\transmit_module.TX_ADDR_9 ));
    InMux I__4130 (
            .O(N__19142),
            .I(N__19139));
    LocalMux I__4129 (
            .O(N__19139),
            .I(N__19136));
    Span4Mux_h I__4128 (
            .O(N__19136),
            .I(N__19133));
    Odrv4 I__4127 (
            .O(N__19133),
            .I(\transmit_module.n107 ));
    CascadeMux I__4126 (
            .O(N__19130),
            .I(\transmit_module.n107_cascade_ ));
    InMux I__4125 (
            .O(N__19127),
            .I(N__19124));
    LocalMux I__4124 (
            .O(N__19124),
            .I(N__19120));
    InMux I__4123 (
            .O(N__19123),
            .I(N__19117));
    Odrv12 I__4122 (
            .O(N__19120),
            .I(\transmit_module.n138 ));
    LocalMux I__4121 (
            .O(N__19117),
            .I(\transmit_module.n138 ));
    CascadeMux I__4120 (
            .O(N__19112),
            .I(N__19109));
    CascadeBuf I__4119 (
            .O(N__19109),
            .I(N__19105));
    CascadeMux I__4118 (
            .O(N__19108),
            .I(N__19102));
    CascadeMux I__4117 (
            .O(N__19105),
            .I(N__19099));
    CascadeBuf I__4116 (
            .O(N__19102),
            .I(N__19096));
    CascadeBuf I__4115 (
            .O(N__19099),
            .I(N__19093));
    CascadeMux I__4114 (
            .O(N__19096),
            .I(N__19090));
    CascadeMux I__4113 (
            .O(N__19093),
            .I(N__19087));
    CascadeBuf I__4112 (
            .O(N__19090),
            .I(N__19084));
    CascadeBuf I__4111 (
            .O(N__19087),
            .I(N__19081));
    CascadeMux I__4110 (
            .O(N__19084),
            .I(N__19078));
    CascadeMux I__4109 (
            .O(N__19081),
            .I(N__19075));
    CascadeBuf I__4108 (
            .O(N__19078),
            .I(N__19072));
    CascadeBuf I__4107 (
            .O(N__19075),
            .I(N__19069));
    CascadeMux I__4106 (
            .O(N__19072),
            .I(N__19066));
    CascadeMux I__4105 (
            .O(N__19069),
            .I(N__19063));
    CascadeBuf I__4104 (
            .O(N__19066),
            .I(N__19060));
    CascadeBuf I__4103 (
            .O(N__19063),
            .I(N__19057));
    CascadeMux I__4102 (
            .O(N__19060),
            .I(N__19054));
    CascadeMux I__4101 (
            .O(N__19057),
            .I(N__19051));
    CascadeBuf I__4100 (
            .O(N__19054),
            .I(N__19048));
    CascadeBuf I__4099 (
            .O(N__19051),
            .I(N__19045));
    CascadeMux I__4098 (
            .O(N__19048),
            .I(N__19042));
    CascadeMux I__4097 (
            .O(N__19045),
            .I(N__19039));
    CascadeBuf I__4096 (
            .O(N__19042),
            .I(N__19036));
    CascadeBuf I__4095 (
            .O(N__19039),
            .I(N__19033));
    CascadeMux I__4094 (
            .O(N__19036),
            .I(N__19030));
    CascadeMux I__4093 (
            .O(N__19033),
            .I(N__19027));
    CascadeBuf I__4092 (
            .O(N__19030),
            .I(N__19024));
    CascadeBuf I__4091 (
            .O(N__19027),
            .I(N__19021));
    CascadeMux I__4090 (
            .O(N__19024),
            .I(N__19018));
    CascadeMux I__4089 (
            .O(N__19021),
            .I(N__19015));
    CascadeBuf I__4088 (
            .O(N__19018),
            .I(N__19012));
    CascadeBuf I__4087 (
            .O(N__19015),
            .I(N__19009));
    CascadeMux I__4086 (
            .O(N__19012),
            .I(N__19006));
    CascadeMux I__4085 (
            .O(N__19009),
            .I(N__19003));
    CascadeBuf I__4084 (
            .O(N__19006),
            .I(N__19000));
    CascadeBuf I__4083 (
            .O(N__19003),
            .I(N__18997));
    CascadeMux I__4082 (
            .O(N__19000),
            .I(N__18994));
    CascadeMux I__4081 (
            .O(N__18997),
            .I(N__18991));
    CascadeBuf I__4080 (
            .O(N__18994),
            .I(N__18988));
    CascadeBuf I__4079 (
            .O(N__18991),
            .I(N__18985));
    CascadeMux I__4078 (
            .O(N__18988),
            .I(N__18982));
    CascadeMux I__4077 (
            .O(N__18985),
            .I(N__18979));
    CascadeBuf I__4076 (
            .O(N__18982),
            .I(N__18976));
    CascadeBuf I__4075 (
            .O(N__18979),
            .I(N__18973));
    CascadeMux I__4074 (
            .O(N__18976),
            .I(N__18970));
    CascadeMux I__4073 (
            .O(N__18973),
            .I(N__18967));
    CascadeBuf I__4072 (
            .O(N__18970),
            .I(N__18964));
    CascadeBuf I__4071 (
            .O(N__18967),
            .I(N__18961));
    CascadeMux I__4070 (
            .O(N__18964),
            .I(N__18958));
    CascadeMux I__4069 (
            .O(N__18961),
            .I(N__18955));
    CascadeBuf I__4068 (
            .O(N__18958),
            .I(N__18952));
    CascadeBuf I__4067 (
            .O(N__18955),
            .I(N__18949));
    CascadeMux I__4066 (
            .O(N__18952),
            .I(N__18946));
    CascadeMux I__4065 (
            .O(N__18949),
            .I(N__18943));
    CascadeBuf I__4064 (
            .O(N__18946),
            .I(N__18940));
    CascadeBuf I__4063 (
            .O(N__18943),
            .I(N__18937));
    CascadeMux I__4062 (
            .O(N__18940),
            .I(N__18934));
    CascadeMux I__4061 (
            .O(N__18937),
            .I(N__18931));
    CascadeBuf I__4060 (
            .O(N__18934),
            .I(N__18928));
    InMux I__4059 (
            .O(N__18931),
            .I(N__18925));
    CascadeMux I__4058 (
            .O(N__18928),
            .I(N__18922));
    LocalMux I__4057 (
            .O(N__18925),
            .I(N__18919));
    InMux I__4056 (
            .O(N__18922),
            .I(N__18916));
    Span4Mux_v I__4055 (
            .O(N__18919),
            .I(N__18913));
    LocalMux I__4054 (
            .O(N__18916),
            .I(N__18910));
    Span4Mux_v I__4053 (
            .O(N__18913),
            .I(N__18907));
    Span12Mux_h I__4052 (
            .O(N__18910),
            .I(N__18904));
    Span4Mux_v I__4051 (
            .O(N__18907),
            .I(N__18901));
    Span12Mux_v I__4050 (
            .O(N__18904),
            .I(N__18898));
    Span4Mux_h I__4049 (
            .O(N__18901),
            .I(N__18895));
    Odrv12 I__4048 (
            .O(N__18898),
            .I(n19));
    Odrv4 I__4047 (
            .O(N__18895),
            .I(n19));
    InMux I__4046 (
            .O(N__18890),
            .I(N__18886));
    InMux I__4045 (
            .O(N__18889),
            .I(N__18883));
    LocalMux I__4044 (
            .O(N__18886),
            .I(N__18880));
    LocalMux I__4043 (
            .O(N__18883),
            .I(N__18877));
    Span12Mux_s2_v I__4042 (
            .O(N__18880),
            .I(N__18874));
    Odrv12 I__4041 (
            .O(N__18877),
            .I(\transmit_module.n114 ));
    Odrv12 I__4040 (
            .O(N__18874),
            .I(\transmit_module.n114 ));
    InMux I__4039 (
            .O(N__18869),
            .I(N__18866));
    LocalMux I__4038 (
            .O(N__18866),
            .I(N__18863));
    Span12Mux_s6_v I__4037 (
            .O(N__18863),
            .I(N__18860));
    Span12Mux_v I__4036 (
            .O(N__18860),
            .I(N__18857));
    Odrv12 I__4035 (
            .O(N__18857),
            .I(\transmit_module.n145 ));
    CascadeMux I__4034 (
            .O(N__18854),
            .I(N__18850));
    CascadeMux I__4033 (
            .O(N__18853),
            .I(N__18847));
    CascadeBuf I__4032 (
            .O(N__18850),
            .I(N__18844));
    CascadeBuf I__4031 (
            .O(N__18847),
            .I(N__18841));
    CascadeMux I__4030 (
            .O(N__18844),
            .I(N__18838));
    CascadeMux I__4029 (
            .O(N__18841),
            .I(N__18835));
    CascadeBuf I__4028 (
            .O(N__18838),
            .I(N__18832));
    CascadeBuf I__4027 (
            .O(N__18835),
            .I(N__18829));
    CascadeMux I__4026 (
            .O(N__18832),
            .I(N__18826));
    CascadeMux I__4025 (
            .O(N__18829),
            .I(N__18823));
    CascadeBuf I__4024 (
            .O(N__18826),
            .I(N__18820));
    CascadeBuf I__4023 (
            .O(N__18823),
            .I(N__18817));
    CascadeMux I__4022 (
            .O(N__18820),
            .I(N__18814));
    CascadeMux I__4021 (
            .O(N__18817),
            .I(N__18811));
    CascadeBuf I__4020 (
            .O(N__18814),
            .I(N__18808));
    CascadeBuf I__4019 (
            .O(N__18811),
            .I(N__18805));
    CascadeMux I__4018 (
            .O(N__18808),
            .I(N__18802));
    CascadeMux I__4017 (
            .O(N__18805),
            .I(N__18799));
    CascadeBuf I__4016 (
            .O(N__18802),
            .I(N__18796));
    CascadeBuf I__4015 (
            .O(N__18799),
            .I(N__18793));
    CascadeMux I__4014 (
            .O(N__18796),
            .I(N__18790));
    CascadeMux I__4013 (
            .O(N__18793),
            .I(N__18787));
    CascadeBuf I__4012 (
            .O(N__18790),
            .I(N__18784));
    CascadeBuf I__4011 (
            .O(N__18787),
            .I(N__18781));
    CascadeMux I__4010 (
            .O(N__18784),
            .I(N__18778));
    CascadeMux I__4009 (
            .O(N__18781),
            .I(N__18775));
    CascadeBuf I__4008 (
            .O(N__18778),
            .I(N__18772));
    CascadeBuf I__4007 (
            .O(N__18775),
            .I(N__18769));
    CascadeMux I__4006 (
            .O(N__18772),
            .I(N__18766));
    CascadeMux I__4005 (
            .O(N__18769),
            .I(N__18763));
    CascadeBuf I__4004 (
            .O(N__18766),
            .I(N__18760));
    CascadeBuf I__4003 (
            .O(N__18763),
            .I(N__18757));
    CascadeMux I__4002 (
            .O(N__18760),
            .I(N__18754));
    CascadeMux I__4001 (
            .O(N__18757),
            .I(N__18751));
    CascadeBuf I__4000 (
            .O(N__18754),
            .I(N__18748));
    CascadeBuf I__3999 (
            .O(N__18751),
            .I(N__18745));
    CascadeMux I__3998 (
            .O(N__18748),
            .I(N__18742));
    CascadeMux I__3997 (
            .O(N__18745),
            .I(N__18739));
    CascadeBuf I__3996 (
            .O(N__18742),
            .I(N__18736));
    CascadeBuf I__3995 (
            .O(N__18739),
            .I(N__18733));
    CascadeMux I__3994 (
            .O(N__18736),
            .I(N__18730));
    CascadeMux I__3993 (
            .O(N__18733),
            .I(N__18727));
    CascadeBuf I__3992 (
            .O(N__18730),
            .I(N__18724));
    CascadeBuf I__3991 (
            .O(N__18727),
            .I(N__18721));
    CascadeMux I__3990 (
            .O(N__18724),
            .I(N__18718));
    CascadeMux I__3989 (
            .O(N__18721),
            .I(N__18715));
    CascadeBuf I__3988 (
            .O(N__18718),
            .I(N__18712));
    CascadeBuf I__3987 (
            .O(N__18715),
            .I(N__18709));
    CascadeMux I__3986 (
            .O(N__18712),
            .I(N__18706));
    CascadeMux I__3985 (
            .O(N__18709),
            .I(N__18703));
    CascadeBuf I__3984 (
            .O(N__18706),
            .I(N__18700));
    CascadeBuf I__3983 (
            .O(N__18703),
            .I(N__18697));
    CascadeMux I__3982 (
            .O(N__18700),
            .I(N__18694));
    CascadeMux I__3981 (
            .O(N__18697),
            .I(N__18691));
    CascadeBuf I__3980 (
            .O(N__18694),
            .I(N__18688));
    CascadeBuf I__3979 (
            .O(N__18691),
            .I(N__18685));
    CascadeMux I__3978 (
            .O(N__18688),
            .I(N__18682));
    CascadeMux I__3977 (
            .O(N__18685),
            .I(N__18679));
    CascadeBuf I__3976 (
            .O(N__18682),
            .I(N__18676));
    CascadeBuf I__3975 (
            .O(N__18679),
            .I(N__18673));
    CascadeMux I__3974 (
            .O(N__18676),
            .I(N__18670));
    CascadeMux I__3973 (
            .O(N__18673),
            .I(N__18667));
    InMux I__3972 (
            .O(N__18670),
            .I(N__18664));
    InMux I__3971 (
            .O(N__18667),
            .I(N__18661));
    LocalMux I__3970 (
            .O(N__18664),
            .I(N__18658));
    LocalMux I__3969 (
            .O(N__18661),
            .I(N__18655));
    Span4Mux_h I__3968 (
            .O(N__18658),
            .I(N__18652));
    Span4Mux_h I__3967 (
            .O(N__18655),
            .I(N__18649));
    Span4Mux_h I__3966 (
            .O(N__18652),
            .I(N__18644));
    Span4Mux_h I__3965 (
            .O(N__18649),
            .I(N__18644));
    Odrv4 I__3964 (
            .O(N__18644),
            .I(n26));
    InMux I__3963 (
            .O(N__18641),
            .I(N__18638));
    LocalMux I__3962 (
            .O(N__18638),
            .I(N__18635));
    Span4Mux_v I__3961 (
            .O(N__18635),
            .I(N__18632));
    Span4Mux_v I__3960 (
            .O(N__18632),
            .I(N__18629));
    Odrv4 I__3959 (
            .O(N__18629),
            .I(\tvp_video_buffer.BUFFER_1_4 ));
    InMux I__3958 (
            .O(N__18626),
            .I(N__18623));
    LocalMux I__3957 (
            .O(N__18623),
            .I(\transmit_module.Y_DELTA_PATTERN_17 ));
    InMux I__3956 (
            .O(N__18620),
            .I(N__18617));
    LocalMux I__3955 (
            .O(N__18617),
            .I(N__18614));
    Span4Mux_h I__3954 (
            .O(N__18614),
            .I(N__18611));
    Span4Mux_h I__3953 (
            .O(N__18611),
            .I(N__18608));
    Odrv4 I__3952 (
            .O(N__18608),
            .I(\transmit_module.Y_DELTA_PATTERN_20 ));
    InMux I__3951 (
            .O(N__18605),
            .I(N__18602));
    LocalMux I__3950 (
            .O(N__18602),
            .I(\transmit_module.Y_DELTA_PATTERN_19 ));
    InMux I__3949 (
            .O(N__18599),
            .I(N__18596));
    LocalMux I__3948 (
            .O(N__18596),
            .I(\transmit_module.Y_DELTA_PATTERN_18 ));
    InMux I__3947 (
            .O(N__18593),
            .I(N__18590));
    LocalMux I__3946 (
            .O(N__18590),
            .I(N__18587));
    Odrv4 I__3945 (
            .O(N__18587),
            .I(\transmit_module.ADDR_Y_COMPONENT_13 ));
    InMux I__3944 (
            .O(N__18584),
            .I(N__18581));
    LocalMux I__3943 (
            .O(N__18581),
            .I(\transmit_module.ADDR_Y_COMPONENT_12 ));
    InMux I__3942 (
            .O(N__18578),
            .I(N__18575));
    LocalMux I__3941 (
            .O(N__18575),
            .I(N__18572));
    Odrv4 I__3940 (
            .O(N__18572),
            .I(\transmit_module.ADDR_Y_COMPONENT_11 ));
    InMux I__3939 (
            .O(N__18569),
            .I(N__18565));
    InMux I__3938 (
            .O(N__18568),
            .I(N__18562));
    LocalMux I__3937 (
            .O(N__18565),
            .I(N__18553));
    LocalMux I__3936 (
            .O(N__18562),
            .I(N__18553));
    InMux I__3935 (
            .O(N__18561),
            .I(N__18550));
    InMux I__3934 (
            .O(N__18560),
            .I(N__18547));
    InMux I__3933 (
            .O(N__18559),
            .I(N__18544));
    InMux I__3932 (
            .O(N__18558),
            .I(N__18541));
    Span4Mux_v I__3931 (
            .O(N__18553),
            .I(N__18533));
    LocalMux I__3930 (
            .O(N__18550),
            .I(N__18533));
    LocalMux I__3929 (
            .O(N__18547),
            .I(N__18533));
    LocalMux I__3928 (
            .O(N__18544),
            .I(N__18529));
    LocalMux I__3927 (
            .O(N__18541),
            .I(N__18526));
    InMux I__3926 (
            .O(N__18540),
            .I(N__18523));
    Span4Mux_v I__3925 (
            .O(N__18533),
            .I(N__18520));
    InMux I__3924 (
            .O(N__18532),
            .I(N__18517));
    Span4Mux_v I__3923 (
            .O(N__18529),
            .I(N__18514));
    Span4Mux_s2_v I__3922 (
            .O(N__18526),
            .I(N__18509));
    LocalMux I__3921 (
            .O(N__18523),
            .I(N__18509));
    Span4Mux_v I__3920 (
            .O(N__18520),
            .I(N__18504));
    LocalMux I__3919 (
            .O(N__18517),
            .I(N__18504));
    Span4Mux_v I__3918 (
            .O(N__18514),
            .I(N__18501));
    Span4Mux_v I__3917 (
            .O(N__18509),
            .I(N__18498));
    Span4Mux_v I__3916 (
            .O(N__18504),
            .I(N__18495));
    Sp12to4 I__3915 (
            .O(N__18501),
            .I(N__18492));
    Span4Mux_h I__3914 (
            .O(N__18498),
            .I(N__18489));
    Span4Mux_h I__3913 (
            .O(N__18495),
            .I(N__18486));
    Span12Mux_h I__3912 (
            .O(N__18492),
            .I(N__18483));
    Span4Mux_h I__3911 (
            .O(N__18489),
            .I(N__18480));
    Span4Mux_h I__3910 (
            .O(N__18486),
            .I(N__18477));
    Odrv12 I__3909 (
            .O(N__18483),
            .I(RX_DATA_6));
    Odrv4 I__3908 (
            .O(N__18480),
            .I(RX_DATA_6));
    Odrv4 I__3907 (
            .O(N__18477),
            .I(RX_DATA_6));
    IoInMux I__3906 (
            .O(N__18470),
            .I(N__18467));
    LocalMux I__3905 (
            .O(N__18467),
            .I(N__18464));
    IoSpan4Mux I__3904 (
            .O(N__18464),
            .I(N__18461));
    Span4Mux_s3_h I__3903 (
            .O(N__18461),
            .I(N__18458));
    Sp12to4 I__3902 (
            .O(N__18458),
            .I(N__18455));
    Span12Mux_v I__3901 (
            .O(N__18455),
            .I(N__18451));
    InMux I__3900 (
            .O(N__18454),
            .I(N__18448));
    Span12Mux_h I__3899 (
            .O(N__18451),
            .I(N__18445));
    LocalMux I__3898 (
            .O(N__18448),
            .I(N__18442));
    Odrv12 I__3897 (
            .O(N__18445),
            .I(DEBUG_c_6_c));
    Odrv12 I__3896 (
            .O(N__18442),
            .I(DEBUG_c_6_c));
    InMux I__3895 (
            .O(N__18437),
            .I(N__18434));
    LocalMux I__3894 (
            .O(N__18434),
            .I(\tvp_video_buffer.BUFFER_0_8 ));
    InMux I__3893 (
            .O(N__18431),
            .I(N__18428));
    LocalMux I__3892 (
            .O(N__18428),
            .I(\tvp_video_buffer.BUFFER_1_8 ));
    InMux I__3891 (
            .O(N__18425),
            .I(N__18422));
    LocalMux I__3890 (
            .O(N__18422),
            .I(N__18419));
    Span4Mux_v I__3889 (
            .O(N__18419),
            .I(N__18415));
    InMux I__3888 (
            .O(N__18418),
            .I(N__18412));
    Odrv4 I__3887 (
            .O(N__18415),
            .I(\transmit_module.n141 ));
    LocalMux I__3886 (
            .O(N__18412),
            .I(\transmit_module.n141 ));
    CEMux I__3885 (
            .O(N__18407),
            .I(N__18403));
    CEMux I__3884 (
            .O(N__18406),
            .I(N__18399));
    LocalMux I__3883 (
            .O(N__18403),
            .I(N__18396));
    CEMux I__3882 (
            .O(N__18402),
            .I(N__18393));
    LocalMux I__3881 (
            .O(N__18399),
            .I(N__18388));
    Span4Mux_h I__3880 (
            .O(N__18396),
            .I(N__18383));
    LocalMux I__3879 (
            .O(N__18393),
            .I(N__18383));
    CEMux I__3878 (
            .O(N__18392),
            .I(N__18379));
    CEMux I__3877 (
            .O(N__18391),
            .I(N__18376));
    Span4Mux_h I__3876 (
            .O(N__18388),
            .I(N__18371));
    Span4Mux_v I__3875 (
            .O(N__18383),
            .I(N__18371));
    SRMux I__3874 (
            .O(N__18382),
            .I(N__18368));
    LocalMux I__3873 (
            .O(N__18379),
            .I(N__18365));
    LocalMux I__3872 (
            .O(N__18376),
            .I(N__18362));
    Span4Mux_h I__3871 (
            .O(N__18371),
            .I(N__18357));
    LocalMux I__3870 (
            .O(N__18368),
            .I(N__18357));
    Span4Mux_v I__3869 (
            .O(N__18365),
            .I(N__18354));
    Span4Mux_v I__3868 (
            .O(N__18362),
            .I(N__18349));
    Span4Mux_h I__3867 (
            .O(N__18357),
            .I(N__18349));
    Span4Mux_h I__3866 (
            .O(N__18354),
            .I(N__18346));
    Span4Mux_h I__3865 (
            .O(N__18349),
            .I(N__18343));
    Odrv4 I__3864 (
            .O(N__18346),
            .I(\transmit_module.n2167 ));
    Odrv4 I__3863 (
            .O(N__18343),
            .I(\transmit_module.n2167 ));
    InMux I__3862 (
            .O(N__18338),
            .I(N__18335));
    LocalMux I__3861 (
            .O(N__18335),
            .I(N__18332));
    Span4Mux_v I__3860 (
            .O(N__18332),
            .I(N__18328));
    InMux I__3859 (
            .O(N__18331),
            .I(N__18325));
    Odrv4 I__3858 (
            .O(N__18328),
            .I(\transmit_module.n140 ));
    LocalMux I__3857 (
            .O(N__18325),
            .I(\transmit_module.n140 ));
    InMux I__3856 (
            .O(N__18320),
            .I(N__18317));
    LocalMux I__3855 (
            .O(N__18317),
            .I(\transmit_module.n130 ));
    CascadeMux I__3854 (
            .O(N__18314),
            .I(\transmit_module.n145_cascade_ ));
    InMux I__3853 (
            .O(N__18311),
            .I(N__18308));
    LocalMux I__3852 (
            .O(N__18308),
            .I(N__18305));
    Span4Mux_h I__3851 (
            .O(N__18305),
            .I(N__18302));
    Odrv4 I__3850 (
            .O(N__18302),
            .I(\transmit_module.Y_DELTA_PATTERN_16 ));
    InMux I__3849 (
            .O(N__18299),
            .I(N__18296));
    LocalMux I__3848 (
            .O(N__18296),
            .I(N__18292));
    InMux I__3847 (
            .O(N__18295),
            .I(N__18289));
    Span4Mux_h I__3846 (
            .O(N__18292),
            .I(N__18283));
    LocalMux I__3845 (
            .O(N__18289),
            .I(N__18283));
    CascadeMux I__3844 (
            .O(N__18288),
            .I(N__18279));
    Span4Mux_v I__3843 (
            .O(N__18283),
            .I(N__18276));
    InMux I__3842 (
            .O(N__18282),
            .I(N__18273));
    InMux I__3841 (
            .O(N__18279),
            .I(N__18270));
    Odrv4 I__3840 (
            .O(N__18276),
            .I(\transmit_module.TX_ADDR_1 ));
    LocalMux I__3839 (
            .O(N__18273),
            .I(\transmit_module.TX_ADDR_1 ));
    LocalMux I__3838 (
            .O(N__18270),
            .I(\transmit_module.TX_ADDR_1 ));
    InMux I__3837 (
            .O(N__18263),
            .I(N__18260));
    LocalMux I__3836 (
            .O(N__18260),
            .I(\transmit_module.ADDR_Y_COMPONENT_1 ));
    InMux I__3835 (
            .O(N__18257),
            .I(N__18254));
    LocalMux I__3834 (
            .O(N__18254),
            .I(N__18251));
    Span12Mux_v I__3833 (
            .O(N__18251),
            .I(N__18248));
    Odrv12 I__3832 (
            .O(N__18248),
            .I(\transmit_module.n128 ));
    InMux I__3831 (
            .O(N__18245),
            .I(N__18242));
    LocalMux I__3830 (
            .O(N__18242),
            .I(N__18239));
    Span4Mux_v I__3829 (
            .O(N__18239),
            .I(N__18235));
    InMux I__3828 (
            .O(N__18238),
            .I(N__18232));
    Span4Mux_v I__3827 (
            .O(N__18235),
            .I(N__18229));
    LocalMux I__3826 (
            .O(N__18232),
            .I(N__18226));
    Span4Mux_h I__3825 (
            .O(N__18229),
            .I(N__18223));
    Odrv12 I__3824 (
            .O(N__18226),
            .I(\transmit_module.n143 ));
    Odrv4 I__3823 (
            .O(N__18223),
            .I(\transmit_module.n143 ));
    SRMux I__3822 (
            .O(N__18218),
            .I(N__18214));
    SRMux I__3821 (
            .O(N__18217),
            .I(N__18209));
    LocalMux I__3820 (
            .O(N__18214),
            .I(N__18204));
    SRMux I__3819 (
            .O(N__18213),
            .I(N__18201));
    SRMux I__3818 (
            .O(N__18212),
            .I(N__18198));
    LocalMux I__3817 (
            .O(N__18209),
            .I(N__18193));
    SRMux I__3816 (
            .O(N__18208),
            .I(N__18190));
    SRMux I__3815 (
            .O(N__18207),
            .I(N__18187));
    Span4Mux_s1_v I__3814 (
            .O(N__18204),
            .I(N__18178));
    LocalMux I__3813 (
            .O(N__18201),
            .I(N__18178));
    LocalMux I__3812 (
            .O(N__18198),
            .I(N__18178));
    SRMux I__3811 (
            .O(N__18197),
            .I(N__18175));
    SRMux I__3810 (
            .O(N__18196),
            .I(N__18172));
    Span4Mux_s1_v I__3809 (
            .O(N__18193),
            .I(N__18163));
    LocalMux I__3808 (
            .O(N__18190),
            .I(N__18163));
    LocalMux I__3807 (
            .O(N__18187),
            .I(N__18163));
    SRMux I__3806 (
            .O(N__18186),
            .I(N__18160));
    SRMux I__3805 (
            .O(N__18185),
            .I(N__18157));
    Span4Mux_v I__3804 (
            .O(N__18178),
            .I(N__18148));
    LocalMux I__3803 (
            .O(N__18175),
            .I(N__18148));
    LocalMux I__3802 (
            .O(N__18172),
            .I(N__18148));
    SRMux I__3801 (
            .O(N__18171),
            .I(N__18145));
    SRMux I__3800 (
            .O(N__18170),
            .I(N__18142));
    Span4Mux_v I__3799 (
            .O(N__18163),
            .I(N__18133));
    LocalMux I__3798 (
            .O(N__18160),
            .I(N__18133));
    LocalMux I__3797 (
            .O(N__18157),
            .I(N__18133));
    SRMux I__3796 (
            .O(N__18156),
            .I(N__18130));
    SRMux I__3795 (
            .O(N__18155),
            .I(N__18127));
    Span4Mux_v I__3794 (
            .O(N__18148),
            .I(N__18117));
    LocalMux I__3793 (
            .O(N__18145),
            .I(N__18117));
    LocalMux I__3792 (
            .O(N__18142),
            .I(N__18117));
    SRMux I__3791 (
            .O(N__18141),
            .I(N__18114));
    SRMux I__3790 (
            .O(N__18140),
            .I(N__18111));
    Span4Mux_v I__3789 (
            .O(N__18133),
            .I(N__18102));
    LocalMux I__3788 (
            .O(N__18130),
            .I(N__18102));
    LocalMux I__3787 (
            .O(N__18127),
            .I(N__18102));
    SRMux I__3786 (
            .O(N__18126),
            .I(N__18099));
    SRMux I__3785 (
            .O(N__18125),
            .I(N__18096));
    SRMux I__3784 (
            .O(N__18124),
            .I(N__18090));
    Span4Mux_v I__3783 (
            .O(N__18117),
            .I(N__18085));
    LocalMux I__3782 (
            .O(N__18114),
            .I(N__18080));
    LocalMux I__3781 (
            .O(N__18111),
            .I(N__18080));
    SRMux I__3780 (
            .O(N__18110),
            .I(N__18077));
    SRMux I__3779 (
            .O(N__18109),
            .I(N__18074));
    Span4Mux_v I__3778 (
            .O(N__18102),
            .I(N__18063));
    LocalMux I__3777 (
            .O(N__18099),
            .I(N__18063));
    LocalMux I__3776 (
            .O(N__18096),
            .I(N__18063));
    SRMux I__3775 (
            .O(N__18095),
            .I(N__18060));
    SRMux I__3774 (
            .O(N__18094),
            .I(N__18057));
    SRMux I__3773 (
            .O(N__18093),
            .I(N__18054));
    LocalMux I__3772 (
            .O(N__18090),
            .I(N__18047));
    SRMux I__3771 (
            .O(N__18089),
            .I(N__18044));
    SRMux I__3770 (
            .O(N__18088),
            .I(N__18041));
    Span4Mux_v I__3769 (
            .O(N__18085),
            .I(N__18038));
    Span4Mux_v I__3768 (
            .O(N__18080),
            .I(N__18031));
    LocalMux I__3767 (
            .O(N__18077),
            .I(N__18031));
    LocalMux I__3766 (
            .O(N__18074),
            .I(N__18031));
    SRMux I__3765 (
            .O(N__18073),
            .I(N__18028));
    SRMux I__3764 (
            .O(N__18072),
            .I(N__18025));
    IoInMux I__3763 (
            .O(N__18071),
            .I(N__18022));
    IoInMux I__3762 (
            .O(N__18070),
            .I(N__18019));
    Span4Mux_v I__3761 (
            .O(N__18063),
            .I(N__18012));
    LocalMux I__3760 (
            .O(N__18060),
            .I(N__18012));
    LocalMux I__3759 (
            .O(N__18057),
            .I(N__18012));
    LocalMux I__3758 (
            .O(N__18054),
            .I(N__18009));
    SRMux I__3757 (
            .O(N__18053),
            .I(N__18006));
    SRMux I__3756 (
            .O(N__18052),
            .I(N__18003));
    SRMux I__3755 (
            .O(N__18051),
            .I(N__18000));
    SRMux I__3754 (
            .O(N__18050),
            .I(N__17997));
    Span4Mux_s2_v I__3753 (
            .O(N__18047),
            .I(N__17990));
    LocalMux I__3752 (
            .O(N__18044),
            .I(N__17990));
    LocalMux I__3751 (
            .O(N__18041),
            .I(N__17990));
    Span4Mux_v I__3750 (
            .O(N__18038),
            .I(N__17981));
    Span4Mux_v I__3749 (
            .O(N__18031),
            .I(N__17981));
    LocalMux I__3748 (
            .O(N__18028),
            .I(N__17981));
    LocalMux I__3747 (
            .O(N__18025),
            .I(N__17981));
    LocalMux I__3746 (
            .O(N__18022),
            .I(N__17976));
    LocalMux I__3745 (
            .O(N__18019),
            .I(N__17976));
    Span4Mux_v I__3744 (
            .O(N__18012),
            .I(N__17973));
    Span4Mux_s2_v I__3743 (
            .O(N__18009),
            .I(N__17966));
    LocalMux I__3742 (
            .O(N__18006),
            .I(N__17966));
    LocalMux I__3741 (
            .O(N__18003),
            .I(N__17966));
    LocalMux I__3740 (
            .O(N__18000),
            .I(N__17961));
    LocalMux I__3739 (
            .O(N__17997),
            .I(N__17961));
    Span4Mux_v I__3738 (
            .O(N__17990),
            .I(N__17956));
    Span4Mux_v I__3737 (
            .O(N__17981),
            .I(N__17956));
    IoSpan4Mux I__3736 (
            .O(N__17976),
            .I(N__17953));
    Span4Mux_h I__3735 (
            .O(N__17973),
            .I(N__17950));
    Span4Mux_v I__3734 (
            .O(N__17966),
            .I(N__17945));
    Span4Mux_v I__3733 (
            .O(N__17961),
            .I(N__17945));
    Span4Mux_h I__3732 (
            .O(N__17956),
            .I(N__17942));
    Span4Mux_s2_v I__3731 (
            .O(N__17953),
            .I(N__17939));
    Span4Mux_v I__3730 (
            .O(N__17950),
            .I(N__17934));
    Span4Mux_h I__3729 (
            .O(N__17945),
            .I(N__17934));
    Span4Mux_h I__3728 (
            .O(N__17942),
            .I(N__17929));
    Span4Mux_v I__3727 (
            .O(N__17939),
            .I(N__17929));
    Odrv4 I__3726 (
            .O(N__17934),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__3725 (
            .O(N__17929),
            .I(CONSTANT_ONE_NET));
    InMux I__3724 (
            .O(N__17924),
            .I(N__17921));
    LocalMux I__3723 (
            .O(N__17921),
            .I(N__17917));
    InMux I__3722 (
            .O(N__17920),
            .I(N__17914));
    Span4Mux_s3_v I__3721 (
            .O(N__17917),
            .I(N__17908));
    LocalMux I__3720 (
            .O(N__17914),
            .I(N__17905));
    InMux I__3719 (
            .O(N__17913),
            .I(N__17902));
    InMux I__3718 (
            .O(N__17912),
            .I(N__17899));
    InMux I__3717 (
            .O(N__17911),
            .I(N__17896));
    Span4Mux_h I__3716 (
            .O(N__17908),
            .I(N__17893));
    Span4Mux_v I__3715 (
            .O(N__17905),
            .I(N__17887));
    LocalMux I__3714 (
            .O(N__17902),
            .I(N__17887));
    LocalMux I__3713 (
            .O(N__17899),
            .I(N__17883));
    LocalMux I__3712 (
            .O(N__17896),
            .I(N__17879));
    Sp12to4 I__3711 (
            .O(N__17893),
            .I(N__17876));
    InMux I__3710 (
            .O(N__17892),
            .I(N__17873));
    Span4Mux_v I__3709 (
            .O(N__17887),
            .I(N__17870));
    InMux I__3708 (
            .O(N__17886),
            .I(N__17867));
    Span4Mux_v I__3707 (
            .O(N__17883),
            .I(N__17864));
    InMux I__3706 (
            .O(N__17882),
            .I(N__17861));
    Span12Mux_s9_h I__3705 (
            .O(N__17879),
            .I(N__17858));
    Span12Mux_h I__3704 (
            .O(N__17876),
            .I(N__17855));
    LocalMux I__3703 (
            .O(N__17873),
            .I(N__17852));
    Span4Mux_v I__3702 (
            .O(N__17870),
            .I(N__17847));
    LocalMux I__3701 (
            .O(N__17867),
            .I(N__17847));
    Span4Mux_v I__3700 (
            .O(N__17864),
            .I(N__17842));
    LocalMux I__3699 (
            .O(N__17861),
            .I(N__17842));
    Span12Mux_v I__3698 (
            .O(N__17858),
            .I(N__17839));
    Span12Mux_v I__3697 (
            .O(N__17855),
            .I(N__17834));
    Span12Mux_s10_h I__3696 (
            .O(N__17852),
            .I(N__17834));
    Span4Mux_v I__3695 (
            .O(N__17847),
            .I(N__17831));
    Span4Mux_h I__3694 (
            .O(N__17842),
            .I(N__17828));
    Span12Mux_v I__3693 (
            .O(N__17839),
            .I(N__17821));
    Span12Mux_v I__3692 (
            .O(N__17834),
            .I(N__17821));
    Sp12to4 I__3691 (
            .O(N__17831),
            .I(N__17821));
    Span4Mux_h I__3690 (
            .O(N__17828),
            .I(N__17818));
    Odrv12 I__3689 (
            .O(N__17821),
            .I(RX_DATA_3));
    Odrv4 I__3688 (
            .O(N__17818),
            .I(RX_DATA_3));
    InMux I__3687 (
            .O(N__17813),
            .I(N__17810));
    LocalMux I__3686 (
            .O(N__17810),
            .I(\tvp_video_buffer.BUFFER_0_5 ));
    InMux I__3685 (
            .O(N__17807),
            .I(N__17804));
    LocalMux I__3684 (
            .O(N__17804),
            .I(\tvp_video_buffer.BUFFER_1_5 ));
    InMux I__3683 (
            .O(N__17801),
            .I(N__17798));
    LocalMux I__3682 (
            .O(N__17798),
            .I(\tvp_video_buffer.BUFFER_0_6 ));
    InMux I__3681 (
            .O(N__17795),
            .I(N__17792));
    LocalMux I__3680 (
            .O(N__17792),
            .I(\tvp_video_buffer.BUFFER_1_6 ));
    InMux I__3679 (
            .O(N__17789),
            .I(N__17785));
    InMux I__3678 (
            .O(N__17788),
            .I(N__17782));
    LocalMux I__3677 (
            .O(N__17785),
            .I(N__17779));
    LocalMux I__3676 (
            .O(N__17782),
            .I(N__17776));
    Span4Mux_h I__3675 (
            .O(N__17779),
            .I(N__17771));
    Span4Mux_v I__3674 (
            .O(N__17776),
            .I(N__17766));
    InMux I__3673 (
            .O(N__17775),
            .I(N__17763));
    InMux I__3672 (
            .O(N__17774),
            .I(N__17758));
    Sp12to4 I__3671 (
            .O(N__17771),
            .I(N__17755));
    InMux I__3670 (
            .O(N__17770),
            .I(N__17752));
    InMux I__3669 (
            .O(N__17769),
            .I(N__17749));
    Span4Mux_v I__3668 (
            .O(N__17766),
            .I(N__17744));
    LocalMux I__3667 (
            .O(N__17763),
            .I(N__17744));
    InMux I__3666 (
            .O(N__17762),
            .I(N__17741));
    InMux I__3665 (
            .O(N__17761),
            .I(N__17738));
    LocalMux I__3664 (
            .O(N__17758),
            .I(N__17735));
    Span12Mux_v I__3663 (
            .O(N__17755),
            .I(N__17732));
    LocalMux I__3662 (
            .O(N__17752),
            .I(N__17729));
    LocalMux I__3661 (
            .O(N__17749),
            .I(N__17726));
    Sp12to4 I__3660 (
            .O(N__17744),
            .I(N__17719));
    LocalMux I__3659 (
            .O(N__17741),
            .I(N__17719));
    LocalMux I__3658 (
            .O(N__17738),
            .I(N__17719));
    Span4Mux_h I__3657 (
            .O(N__17735),
            .I(N__17716));
    Span12Mux_v I__3656 (
            .O(N__17732),
            .I(N__17713));
    Span12Mux_h I__3655 (
            .O(N__17729),
            .I(N__17708));
    Span12Mux_h I__3654 (
            .O(N__17726),
            .I(N__17708));
    Span12Mux_v I__3653 (
            .O(N__17719),
            .I(N__17705));
    Span4Mux_h I__3652 (
            .O(N__17716),
            .I(N__17702));
    Odrv12 I__3651 (
            .O(N__17713),
            .I(RX_DATA_4));
    Odrv12 I__3650 (
            .O(N__17708),
            .I(RX_DATA_4));
    Odrv12 I__3649 (
            .O(N__17705),
            .I(RX_DATA_4));
    Odrv4 I__3648 (
            .O(N__17702),
            .I(RX_DATA_4));
    InMux I__3647 (
            .O(N__17693),
            .I(N__17690));
    LocalMux I__3646 (
            .O(N__17690),
            .I(\tvp_video_buffer.BUFFER_1_7 ));
    InMux I__3645 (
            .O(N__17687),
            .I(N__17684));
    LocalMux I__3644 (
            .O(N__17684),
            .I(N__17681));
    Span4Mux_v I__3643 (
            .O(N__17681),
            .I(N__17678));
    Span4Mux_v I__3642 (
            .O(N__17678),
            .I(N__17674));
    InMux I__3641 (
            .O(N__17677),
            .I(N__17668));
    Span4Mux_v I__3640 (
            .O(N__17674),
            .I(N__17665));
    InMux I__3639 (
            .O(N__17673),
            .I(N__17662));
    InMux I__3638 (
            .O(N__17672),
            .I(N__17659));
    InMux I__3637 (
            .O(N__17671),
            .I(N__17655));
    LocalMux I__3636 (
            .O(N__17668),
            .I(N__17651));
    Span4Mux_v I__3635 (
            .O(N__17665),
            .I(N__17646));
    LocalMux I__3634 (
            .O(N__17662),
            .I(N__17646));
    LocalMux I__3633 (
            .O(N__17659),
            .I(N__17642));
    InMux I__3632 (
            .O(N__17658),
            .I(N__17639));
    LocalMux I__3631 (
            .O(N__17655),
            .I(N__17636));
    InMux I__3630 (
            .O(N__17654),
            .I(N__17633));
    Span4Mux_s2_v I__3629 (
            .O(N__17651),
            .I(N__17630));
    Span4Mux_v I__3628 (
            .O(N__17646),
            .I(N__17627));
    InMux I__3627 (
            .O(N__17645),
            .I(N__17624));
    Sp12to4 I__3626 (
            .O(N__17642),
            .I(N__17621));
    LocalMux I__3625 (
            .O(N__17639),
            .I(N__17618));
    Span4Mux_v I__3624 (
            .O(N__17636),
            .I(N__17615));
    LocalMux I__3623 (
            .O(N__17633),
            .I(N__17612));
    Span4Mux_v I__3622 (
            .O(N__17630),
            .I(N__17605));
    Span4Mux_v I__3621 (
            .O(N__17627),
            .I(N__17605));
    LocalMux I__3620 (
            .O(N__17624),
            .I(N__17605));
    Span12Mux_v I__3619 (
            .O(N__17621),
            .I(N__17600));
    Sp12to4 I__3618 (
            .O(N__17618),
            .I(N__17600));
    Span4Mux_v I__3617 (
            .O(N__17615),
            .I(N__17597));
    Sp12to4 I__3616 (
            .O(N__17612),
            .I(N__17594));
    Span4Mux_h I__3615 (
            .O(N__17605),
            .I(N__17591));
    Span12Mux_v I__3614 (
            .O(N__17600),
            .I(N__17584));
    Sp12to4 I__3613 (
            .O(N__17597),
            .I(N__17584));
    Span12Mux_s7_v I__3612 (
            .O(N__17594),
            .I(N__17584));
    Span4Mux_h I__3611 (
            .O(N__17591),
            .I(N__17581));
    Odrv12 I__3610 (
            .O(N__17584),
            .I(RX_DATA_5));
    Odrv4 I__3609 (
            .O(N__17581),
            .I(RX_DATA_5));
    InMux I__3608 (
            .O(N__17576),
            .I(N__17573));
    LocalMux I__3607 (
            .O(N__17573),
            .I(N__17570));
    Odrv4 I__3606 (
            .O(N__17570),
            .I(\transmit_module.n121 ));
    InMux I__3605 (
            .O(N__17567),
            .I(N__17564));
    LocalMux I__3604 (
            .O(N__17564),
            .I(N__17561));
    Odrv4 I__3603 (
            .O(N__17561),
            .I(\transmit_module.n119 ));
    CEMux I__3602 (
            .O(N__17558),
            .I(N__17555));
    LocalMux I__3601 (
            .O(N__17555),
            .I(N__17552));
    Odrv4 I__3600 (
            .O(N__17552),
            .I(\transmit_module.n2057 ));
    InMux I__3599 (
            .O(N__17549),
            .I(N__17546));
    LocalMux I__3598 (
            .O(N__17546),
            .I(N__17543));
    Odrv12 I__3597 (
            .O(N__17543),
            .I(\transmit_module.n124 ));
    InMux I__3596 (
            .O(N__17540),
            .I(N__17537));
    LocalMux I__3595 (
            .O(N__17537),
            .I(N__17534));
    Odrv12 I__3594 (
            .O(N__17534),
            .I(\transmit_module.n126 ));
    InMux I__3593 (
            .O(N__17531),
            .I(N__17528));
    LocalMux I__3592 (
            .O(N__17528),
            .I(N__17525));
    Odrv12 I__3591 (
            .O(N__17525),
            .I(\transmit_module.n123 ));
    InMux I__3590 (
            .O(N__17522),
            .I(N__17519));
    LocalMux I__3589 (
            .O(N__17519),
            .I(N__17516));
    Odrv12 I__3588 (
            .O(N__17516),
            .I(\transmit_module.n125 ));
    CascadeMux I__3587 (
            .O(N__17513),
            .I(N__17510));
    CascadeBuf I__3586 (
            .O(N__17510),
            .I(N__17506));
    CascadeMux I__3585 (
            .O(N__17509),
            .I(N__17503));
    CascadeMux I__3584 (
            .O(N__17506),
            .I(N__17500));
    CascadeBuf I__3583 (
            .O(N__17503),
            .I(N__17497));
    CascadeBuf I__3582 (
            .O(N__17500),
            .I(N__17494));
    CascadeMux I__3581 (
            .O(N__17497),
            .I(N__17491));
    CascadeMux I__3580 (
            .O(N__17494),
            .I(N__17488));
    CascadeBuf I__3579 (
            .O(N__17491),
            .I(N__17485));
    CascadeBuf I__3578 (
            .O(N__17488),
            .I(N__17482));
    CascadeMux I__3577 (
            .O(N__17485),
            .I(N__17479));
    CascadeMux I__3576 (
            .O(N__17482),
            .I(N__17476));
    CascadeBuf I__3575 (
            .O(N__17479),
            .I(N__17473));
    CascadeBuf I__3574 (
            .O(N__17476),
            .I(N__17470));
    CascadeMux I__3573 (
            .O(N__17473),
            .I(N__17467));
    CascadeMux I__3572 (
            .O(N__17470),
            .I(N__17464));
    CascadeBuf I__3571 (
            .O(N__17467),
            .I(N__17461));
    CascadeBuf I__3570 (
            .O(N__17464),
            .I(N__17458));
    CascadeMux I__3569 (
            .O(N__17461),
            .I(N__17455));
    CascadeMux I__3568 (
            .O(N__17458),
            .I(N__17452));
    CascadeBuf I__3567 (
            .O(N__17455),
            .I(N__17449));
    CascadeBuf I__3566 (
            .O(N__17452),
            .I(N__17446));
    CascadeMux I__3565 (
            .O(N__17449),
            .I(N__17443));
    CascadeMux I__3564 (
            .O(N__17446),
            .I(N__17440));
    CascadeBuf I__3563 (
            .O(N__17443),
            .I(N__17437));
    CascadeBuf I__3562 (
            .O(N__17440),
            .I(N__17434));
    CascadeMux I__3561 (
            .O(N__17437),
            .I(N__17431));
    CascadeMux I__3560 (
            .O(N__17434),
            .I(N__17428));
    CascadeBuf I__3559 (
            .O(N__17431),
            .I(N__17425));
    CascadeBuf I__3558 (
            .O(N__17428),
            .I(N__17422));
    CascadeMux I__3557 (
            .O(N__17425),
            .I(N__17419));
    CascadeMux I__3556 (
            .O(N__17422),
            .I(N__17416));
    CascadeBuf I__3555 (
            .O(N__17419),
            .I(N__17413));
    CascadeBuf I__3554 (
            .O(N__17416),
            .I(N__17410));
    CascadeMux I__3553 (
            .O(N__17413),
            .I(N__17407));
    CascadeMux I__3552 (
            .O(N__17410),
            .I(N__17404));
    CascadeBuf I__3551 (
            .O(N__17407),
            .I(N__17401));
    CascadeBuf I__3550 (
            .O(N__17404),
            .I(N__17398));
    CascadeMux I__3549 (
            .O(N__17401),
            .I(N__17395));
    CascadeMux I__3548 (
            .O(N__17398),
            .I(N__17392));
    CascadeBuf I__3547 (
            .O(N__17395),
            .I(N__17389));
    CascadeBuf I__3546 (
            .O(N__17392),
            .I(N__17386));
    CascadeMux I__3545 (
            .O(N__17389),
            .I(N__17383));
    CascadeMux I__3544 (
            .O(N__17386),
            .I(N__17380));
    CascadeBuf I__3543 (
            .O(N__17383),
            .I(N__17377));
    CascadeBuf I__3542 (
            .O(N__17380),
            .I(N__17374));
    CascadeMux I__3541 (
            .O(N__17377),
            .I(N__17371));
    CascadeMux I__3540 (
            .O(N__17374),
            .I(N__17368));
    CascadeBuf I__3539 (
            .O(N__17371),
            .I(N__17365));
    CascadeBuf I__3538 (
            .O(N__17368),
            .I(N__17362));
    CascadeMux I__3537 (
            .O(N__17365),
            .I(N__17359));
    CascadeMux I__3536 (
            .O(N__17362),
            .I(N__17356));
    CascadeBuf I__3535 (
            .O(N__17359),
            .I(N__17353));
    CascadeBuf I__3534 (
            .O(N__17356),
            .I(N__17350));
    CascadeMux I__3533 (
            .O(N__17353),
            .I(N__17347));
    CascadeMux I__3532 (
            .O(N__17350),
            .I(N__17344));
    CascadeBuf I__3531 (
            .O(N__17347),
            .I(N__17341));
    CascadeBuf I__3530 (
            .O(N__17344),
            .I(N__17338));
    CascadeMux I__3529 (
            .O(N__17341),
            .I(N__17335));
    CascadeMux I__3528 (
            .O(N__17338),
            .I(N__17332));
    CascadeBuf I__3527 (
            .O(N__17335),
            .I(N__17329));
    InMux I__3526 (
            .O(N__17332),
            .I(N__17326));
    CascadeMux I__3525 (
            .O(N__17329),
            .I(N__17323));
    LocalMux I__3524 (
            .O(N__17326),
            .I(N__17320));
    InMux I__3523 (
            .O(N__17323),
            .I(N__17317));
    Span4Mux_v I__3522 (
            .O(N__17320),
            .I(N__17314));
    LocalMux I__3521 (
            .O(N__17317),
            .I(N__17311));
    Span4Mux_v I__3520 (
            .O(N__17314),
            .I(N__17308));
    Span4Mux_v I__3519 (
            .O(N__17311),
            .I(N__17305));
    Span4Mux_v I__3518 (
            .O(N__17308),
            .I(N__17302));
    Span4Mux_v I__3517 (
            .O(N__17305),
            .I(N__17299));
    Span4Mux_h I__3516 (
            .O(N__17302),
            .I(N__17296));
    Span4Mux_v I__3515 (
            .O(N__17299),
            .I(N__17293));
    Span4Mux_h I__3514 (
            .O(N__17296),
            .I(N__17288));
    Span4Mux_h I__3513 (
            .O(N__17293),
            .I(N__17288));
    Odrv4 I__3512 (
            .O(N__17288),
            .I(n22));
    InMux I__3511 (
            .O(N__17285),
            .I(N__17282));
    LocalMux I__3510 (
            .O(N__17282),
            .I(N__17279));
    Odrv12 I__3509 (
            .O(N__17279),
            .I(\transmit_module.ADDR_Y_COMPONENT_8 ));
    InMux I__3508 (
            .O(N__17276),
            .I(N__17273));
    LocalMux I__3507 (
            .O(N__17273),
            .I(N__17268));
    InMux I__3506 (
            .O(N__17272),
            .I(N__17265));
    CascadeMux I__3505 (
            .O(N__17271),
            .I(N__17261));
    Span4Mux_v I__3504 (
            .O(N__17268),
            .I(N__17256));
    LocalMux I__3503 (
            .O(N__17265),
            .I(N__17256));
    InMux I__3502 (
            .O(N__17264),
            .I(N__17251));
    InMux I__3501 (
            .O(N__17261),
            .I(N__17251));
    Odrv4 I__3500 (
            .O(N__17256),
            .I(\transmit_module.TX_ADDR_8 ));
    LocalMux I__3499 (
            .O(N__17251),
            .I(\transmit_module.TX_ADDR_8 ));
    CascadeMux I__3498 (
            .O(N__17246),
            .I(N__17242));
    CascadeMux I__3497 (
            .O(N__17245),
            .I(N__17239));
    CascadeBuf I__3496 (
            .O(N__17242),
            .I(N__17236));
    CascadeBuf I__3495 (
            .O(N__17239),
            .I(N__17233));
    CascadeMux I__3494 (
            .O(N__17236),
            .I(N__17230));
    CascadeMux I__3493 (
            .O(N__17233),
            .I(N__17227));
    CascadeBuf I__3492 (
            .O(N__17230),
            .I(N__17224));
    CascadeBuf I__3491 (
            .O(N__17227),
            .I(N__17221));
    CascadeMux I__3490 (
            .O(N__17224),
            .I(N__17218));
    CascadeMux I__3489 (
            .O(N__17221),
            .I(N__17215));
    CascadeBuf I__3488 (
            .O(N__17218),
            .I(N__17212));
    CascadeBuf I__3487 (
            .O(N__17215),
            .I(N__17209));
    CascadeMux I__3486 (
            .O(N__17212),
            .I(N__17206));
    CascadeMux I__3485 (
            .O(N__17209),
            .I(N__17203));
    CascadeBuf I__3484 (
            .O(N__17206),
            .I(N__17200));
    CascadeBuf I__3483 (
            .O(N__17203),
            .I(N__17197));
    CascadeMux I__3482 (
            .O(N__17200),
            .I(N__17194));
    CascadeMux I__3481 (
            .O(N__17197),
            .I(N__17191));
    CascadeBuf I__3480 (
            .O(N__17194),
            .I(N__17188));
    CascadeBuf I__3479 (
            .O(N__17191),
            .I(N__17185));
    CascadeMux I__3478 (
            .O(N__17188),
            .I(N__17182));
    CascadeMux I__3477 (
            .O(N__17185),
            .I(N__17179));
    CascadeBuf I__3476 (
            .O(N__17182),
            .I(N__17176));
    CascadeBuf I__3475 (
            .O(N__17179),
            .I(N__17173));
    CascadeMux I__3474 (
            .O(N__17176),
            .I(N__17170));
    CascadeMux I__3473 (
            .O(N__17173),
            .I(N__17167));
    CascadeBuf I__3472 (
            .O(N__17170),
            .I(N__17164));
    CascadeBuf I__3471 (
            .O(N__17167),
            .I(N__17161));
    CascadeMux I__3470 (
            .O(N__17164),
            .I(N__17158));
    CascadeMux I__3469 (
            .O(N__17161),
            .I(N__17155));
    CascadeBuf I__3468 (
            .O(N__17158),
            .I(N__17152));
    CascadeBuf I__3467 (
            .O(N__17155),
            .I(N__17149));
    CascadeMux I__3466 (
            .O(N__17152),
            .I(N__17146));
    CascadeMux I__3465 (
            .O(N__17149),
            .I(N__17143));
    CascadeBuf I__3464 (
            .O(N__17146),
            .I(N__17140));
    CascadeBuf I__3463 (
            .O(N__17143),
            .I(N__17137));
    CascadeMux I__3462 (
            .O(N__17140),
            .I(N__17134));
    CascadeMux I__3461 (
            .O(N__17137),
            .I(N__17131));
    CascadeBuf I__3460 (
            .O(N__17134),
            .I(N__17128));
    CascadeBuf I__3459 (
            .O(N__17131),
            .I(N__17125));
    CascadeMux I__3458 (
            .O(N__17128),
            .I(N__17122));
    CascadeMux I__3457 (
            .O(N__17125),
            .I(N__17119));
    CascadeBuf I__3456 (
            .O(N__17122),
            .I(N__17116));
    CascadeBuf I__3455 (
            .O(N__17119),
            .I(N__17113));
    CascadeMux I__3454 (
            .O(N__17116),
            .I(N__17110));
    CascadeMux I__3453 (
            .O(N__17113),
            .I(N__17107));
    CascadeBuf I__3452 (
            .O(N__17110),
            .I(N__17104));
    CascadeBuf I__3451 (
            .O(N__17107),
            .I(N__17101));
    CascadeMux I__3450 (
            .O(N__17104),
            .I(N__17098));
    CascadeMux I__3449 (
            .O(N__17101),
            .I(N__17095));
    CascadeBuf I__3448 (
            .O(N__17098),
            .I(N__17092));
    CascadeBuf I__3447 (
            .O(N__17095),
            .I(N__17089));
    CascadeMux I__3446 (
            .O(N__17092),
            .I(N__17086));
    CascadeMux I__3445 (
            .O(N__17089),
            .I(N__17083));
    CascadeBuf I__3444 (
            .O(N__17086),
            .I(N__17080));
    CascadeBuf I__3443 (
            .O(N__17083),
            .I(N__17077));
    CascadeMux I__3442 (
            .O(N__17080),
            .I(N__17074));
    CascadeMux I__3441 (
            .O(N__17077),
            .I(N__17071));
    CascadeBuf I__3440 (
            .O(N__17074),
            .I(N__17068));
    CascadeBuf I__3439 (
            .O(N__17071),
            .I(N__17065));
    CascadeMux I__3438 (
            .O(N__17068),
            .I(N__17062));
    CascadeMux I__3437 (
            .O(N__17065),
            .I(N__17059));
    InMux I__3436 (
            .O(N__17062),
            .I(N__17056));
    InMux I__3435 (
            .O(N__17059),
            .I(N__17053));
    LocalMux I__3434 (
            .O(N__17056),
            .I(N__17050));
    LocalMux I__3433 (
            .O(N__17053),
            .I(N__17047));
    Sp12to4 I__3432 (
            .O(N__17050),
            .I(N__17044));
    Span4Mux_h I__3431 (
            .O(N__17047),
            .I(N__17041));
    Span12Mux_h I__3430 (
            .O(N__17044),
            .I(N__17038));
    Sp12to4 I__3429 (
            .O(N__17041),
            .I(N__17035));
    Span12Mux_v I__3428 (
            .O(N__17038),
            .I(N__17030));
    Span12Mux_v I__3427 (
            .O(N__17035),
            .I(N__17030));
    Odrv12 I__3426 (
            .O(N__17030),
            .I(n21));
    InMux I__3425 (
            .O(N__17027),
            .I(N__17024));
    LocalMux I__3424 (
            .O(N__17024),
            .I(\transmit_module.ADDR_Y_COMPONENT_5 ));
    InMux I__3423 (
            .O(N__17021),
            .I(N__17017));
    CascadeMux I__3422 (
            .O(N__17020),
            .I(N__17012));
    LocalMux I__3421 (
            .O(N__17017),
            .I(N__17009));
    InMux I__3420 (
            .O(N__17016),
            .I(N__17006));
    InMux I__3419 (
            .O(N__17015),
            .I(N__17003));
    InMux I__3418 (
            .O(N__17012),
            .I(N__17000));
    Odrv4 I__3417 (
            .O(N__17009),
            .I(\transmit_module.TX_ADDR_5 ));
    LocalMux I__3416 (
            .O(N__17006),
            .I(\transmit_module.TX_ADDR_5 ));
    LocalMux I__3415 (
            .O(N__17003),
            .I(\transmit_module.TX_ADDR_5 ));
    LocalMux I__3414 (
            .O(N__17000),
            .I(\transmit_module.TX_ADDR_5 ));
    InMux I__3413 (
            .O(N__16991),
            .I(N__16988));
    LocalMux I__3412 (
            .O(N__16988),
            .I(\transmit_module.n111 ));
    CascadeMux I__3411 (
            .O(N__16985),
            .I(\transmit_module.n111_cascade_ ));
    InMux I__3410 (
            .O(N__16982),
            .I(N__16979));
    LocalMux I__3409 (
            .O(N__16979),
            .I(\transmit_module.n142 ));
    CascadeMux I__3408 (
            .O(N__16976),
            .I(N__16973));
    CascadeBuf I__3407 (
            .O(N__16973),
            .I(N__16969));
    CascadeMux I__3406 (
            .O(N__16972),
            .I(N__16966));
    CascadeMux I__3405 (
            .O(N__16969),
            .I(N__16963));
    CascadeBuf I__3404 (
            .O(N__16966),
            .I(N__16960));
    CascadeBuf I__3403 (
            .O(N__16963),
            .I(N__16957));
    CascadeMux I__3402 (
            .O(N__16960),
            .I(N__16954));
    CascadeMux I__3401 (
            .O(N__16957),
            .I(N__16951));
    CascadeBuf I__3400 (
            .O(N__16954),
            .I(N__16948));
    CascadeBuf I__3399 (
            .O(N__16951),
            .I(N__16945));
    CascadeMux I__3398 (
            .O(N__16948),
            .I(N__16942));
    CascadeMux I__3397 (
            .O(N__16945),
            .I(N__16939));
    CascadeBuf I__3396 (
            .O(N__16942),
            .I(N__16936));
    CascadeBuf I__3395 (
            .O(N__16939),
            .I(N__16933));
    CascadeMux I__3394 (
            .O(N__16936),
            .I(N__16930));
    CascadeMux I__3393 (
            .O(N__16933),
            .I(N__16927));
    CascadeBuf I__3392 (
            .O(N__16930),
            .I(N__16924));
    CascadeBuf I__3391 (
            .O(N__16927),
            .I(N__16921));
    CascadeMux I__3390 (
            .O(N__16924),
            .I(N__16918));
    CascadeMux I__3389 (
            .O(N__16921),
            .I(N__16915));
    CascadeBuf I__3388 (
            .O(N__16918),
            .I(N__16912));
    CascadeBuf I__3387 (
            .O(N__16915),
            .I(N__16909));
    CascadeMux I__3386 (
            .O(N__16912),
            .I(N__16906));
    CascadeMux I__3385 (
            .O(N__16909),
            .I(N__16903));
    CascadeBuf I__3384 (
            .O(N__16906),
            .I(N__16900));
    CascadeBuf I__3383 (
            .O(N__16903),
            .I(N__16897));
    CascadeMux I__3382 (
            .O(N__16900),
            .I(N__16894));
    CascadeMux I__3381 (
            .O(N__16897),
            .I(N__16891));
    CascadeBuf I__3380 (
            .O(N__16894),
            .I(N__16888));
    CascadeBuf I__3379 (
            .O(N__16891),
            .I(N__16885));
    CascadeMux I__3378 (
            .O(N__16888),
            .I(N__16882));
    CascadeMux I__3377 (
            .O(N__16885),
            .I(N__16879));
    CascadeBuf I__3376 (
            .O(N__16882),
            .I(N__16876));
    CascadeBuf I__3375 (
            .O(N__16879),
            .I(N__16873));
    CascadeMux I__3374 (
            .O(N__16876),
            .I(N__16870));
    CascadeMux I__3373 (
            .O(N__16873),
            .I(N__16867));
    CascadeBuf I__3372 (
            .O(N__16870),
            .I(N__16864));
    CascadeBuf I__3371 (
            .O(N__16867),
            .I(N__16861));
    CascadeMux I__3370 (
            .O(N__16864),
            .I(N__16858));
    CascadeMux I__3369 (
            .O(N__16861),
            .I(N__16855));
    CascadeBuf I__3368 (
            .O(N__16858),
            .I(N__16852));
    CascadeBuf I__3367 (
            .O(N__16855),
            .I(N__16849));
    CascadeMux I__3366 (
            .O(N__16852),
            .I(N__16846));
    CascadeMux I__3365 (
            .O(N__16849),
            .I(N__16843));
    CascadeBuf I__3364 (
            .O(N__16846),
            .I(N__16840));
    CascadeBuf I__3363 (
            .O(N__16843),
            .I(N__16837));
    CascadeMux I__3362 (
            .O(N__16840),
            .I(N__16834));
    CascadeMux I__3361 (
            .O(N__16837),
            .I(N__16831));
    CascadeBuf I__3360 (
            .O(N__16834),
            .I(N__16828));
    CascadeBuf I__3359 (
            .O(N__16831),
            .I(N__16825));
    CascadeMux I__3358 (
            .O(N__16828),
            .I(N__16822));
    CascadeMux I__3357 (
            .O(N__16825),
            .I(N__16819));
    CascadeBuf I__3356 (
            .O(N__16822),
            .I(N__16816));
    CascadeBuf I__3355 (
            .O(N__16819),
            .I(N__16813));
    CascadeMux I__3354 (
            .O(N__16816),
            .I(N__16810));
    CascadeMux I__3353 (
            .O(N__16813),
            .I(N__16807));
    CascadeBuf I__3352 (
            .O(N__16810),
            .I(N__16804));
    CascadeBuf I__3351 (
            .O(N__16807),
            .I(N__16801));
    CascadeMux I__3350 (
            .O(N__16804),
            .I(N__16798));
    CascadeMux I__3349 (
            .O(N__16801),
            .I(N__16795));
    CascadeBuf I__3348 (
            .O(N__16798),
            .I(N__16792));
    InMux I__3347 (
            .O(N__16795),
            .I(N__16789));
    CascadeMux I__3346 (
            .O(N__16792),
            .I(N__16786));
    LocalMux I__3345 (
            .O(N__16789),
            .I(N__16783));
    InMux I__3344 (
            .O(N__16786),
            .I(N__16780));
    Span4Mux_v I__3343 (
            .O(N__16783),
            .I(N__16777));
    LocalMux I__3342 (
            .O(N__16780),
            .I(N__16774));
    Span4Mux_v I__3341 (
            .O(N__16777),
            .I(N__16771));
    Span4Mux_v I__3340 (
            .O(N__16774),
            .I(N__16768));
    Span4Mux_v I__3339 (
            .O(N__16771),
            .I(N__16765));
    Span4Mux_v I__3338 (
            .O(N__16768),
            .I(N__16762));
    Span4Mux_v I__3337 (
            .O(N__16765),
            .I(N__16759));
    Span4Mux_v I__3336 (
            .O(N__16762),
            .I(N__16756));
    Span4Mux_h I__3335 (
            .O(N__16759),
            .I(N__16753));
    Span4Mux_v I__3334 (
            .O(N__16756),
            .I(N__16750));
    Span4Mux_h I__3333 (
            .O(N__16753),
            .I(N__16745));
    Span4Mux_h I__3332 (
            .O(N__16750),
            .I(N__16745));
    Odrv4 I__3331 (
            .O(N__16745),
            .I(n23));
    InMux I__3330 (
            .O(N__16742),
            .I(N__16739));
    LocalMux I__3329 (
            .O(N__16739),
            .I(\transmit_module.video_signal_controller.VGA_VISIBLE_N_580 ));
    InMux I__3328 (
            .O(N__16736),
            .I(N__16732));
    InMux I__3327 (
            .O(N__16735),
            .I(N__16729));
    LocalMux I__3326 (
            .O(N__16732),
            .I(N__16726));
    LocalMux I__3325 (
            .O(N__16729),
            .I(\transmit_module.video_signal_controller.n3333 ));
    Odrv4 I__3324 (
            .O(N__16726),
            .I(\transmit_module.video_signal_controller.n3333 ));
    CascadeMux I__3323 (
            .O(N__16721),
            .I(N__16718));
    InMux I__3322 (
            .O(N__16718),
            .I(N__16713));
    InMux I__3321 (
            .O(N__16717),
            .I(N__16708));
    InMux I__3320 (
            .O(N__16716),
            .I(N__16705));
    LocalMux I__3319 (
            .O(N__16713),
            .I(N__16702));
    InMux I__3318 (
            .O(N__16712),
            .I(N__16697));
    InMux I__3317 (
            .O(N__16711),
            .I(N__16697));
    LocalMux I__3316 (
            .O(N__16708),
            .I(N__16694));
    LocalMux I__3315 (
            .O(N__16705),
            .I(\transmit_module.video_signal_controller.VGA_X_11 ));
    Odrv4 I__3314 (
            .O(N__16702),
            .I(\transmit_module.video_signal_controller.VGA_X_11 ));
    LocalMux I__3313 (
            .O(N__16697),
            .I(\transmit_module.video_signal_controller.VGA_X_11 ));
    Odrv4 I__3312 (
            .O(N__16694),
            .I(\transmit_module.video_signal_controller.VGA_X_11 ));
    InMux I__3311 (
            .O(N__16685),
            .I(N__16682));
    LocalMux I__3310 (
            .O(N__16682),
            .I(N__16679));
    Span4Mux_h I__3309 (
            .O(N__16679),
            .I(N__16676));
    Odrv4 I__3308 (
            .O(N__16676),
            .I(\transmit_module.video_signal_controller.n7 ));
    InMux I__3307 (
            .O(N__16673),
            .I(N__16670));
    LocalMux I__3306 (
            .O(N__16670),
            .I(\transmit_module.ADDR_Y_COMPONENT_10 ));
    InMux I__3305 (
            .O(N__16667),
            .I(N__16661));
    InMux I__3304 (
            .O(N__16666),
            .I(N__16658));
    InMux I__3303 (
            .O(N__16665),
            .I(N__16655));
    InMux I__3302 (
            .O(N__16664),
            .I(N__16652));
    LocalMux I__3301 (
            .O(N__16661),
            .I(\transmit_module.TX_ADDR_10 ));
    LocalMux I__3300 (
            .O(N__16658),
            .I(\transmit_module.TX_ADDR_10 ));
    LocalMux I__3299 (
            .O(N__16655),
            .I(\transmit_module.TX_ADDR_10 ));
    LocalMux I__3298 (
            .O(N__16652),
            .I(\transmit_module.TX_ADDR_10 ));
    InMux I__3297 (
            .O(N__16643),
            .I(N__16639));
    InMux I__3296 (
            .O(N__16642),
            .I(N__16636));
    LocalMux I__3295 (
            .O(N__16639),
            .I(N__16633));
    LocalMux I__3294 (
            .O(N__16636),
            .I(\transmit_module.n106 ));
    Odrv4 I__3293 (
            .O(N__16633),
            .I(\transmit_module.n106 ));
    InMux I__3292 (
            .O(N__16628),
            .I(N__16625));
    LocalMux I__3291 (
            .O(N__16625),
            .I(N__16622));
    Odrv4 I__3290 (
            .O(N__16622),
            .I(\transmit_module.n120 ));
    InMux I__3289 (
            .O(N__16619),
            .I(\transmit_module.n3110 ));
    InMux I__3288 (
            .O(N__16616),
            .I(bfn_15_14_0_));
    InMux I__3287 (
            .O(N__16613),
            .I(\transmit_module.n3112 ));
    InMux I__3286 (
            .O(N__16610),
            .I(N__16607));
    LocalMux I__3285 (
            .O(N__16607),
            .I(\transmit_module.n122 ));
    InMux I__3284 (
            .O(N__16604),
            .I(\transmit_module.n3113 ));
    InMux I__3283 (
            .O(N__16601),
            .I(\transmit_module.n3114 ));
    InMux I__3282 (
            .O(N__16598),
            .I(\transmit_module.n3115 ));
    InMux I__3281 (
            .O(N__16595),
            .I(\transmit_module.n3116 ));
    IoInMux I__3280 (
            .O(N__16592),
            .I(N__16589));
    LocalMux I__3279 (
            .O(N__16589),
            .I(N__16586));
    IoSpan4Mux I__3278 (
            .O(N__16586),
            .I(N__16583));
    Span4Mux_s2_h I__3277 (
            .O(N__16583),
            .I(N__16580));
    Sp12to4 I__3276 (
            .O(N__16580),
            .I(N__16577));
    Span12Mux_v I__3275 (
            .O(N__16577),
            .I(N__16573));
    InMux I__3274 (
            .O(N__16576),
            .I(N__16570));
    Span12Mux_h I__3273 (
            .O(N__16573),
            .I(N__16567));
    LocalMux I__3272 (
            .O(N__16570),
            .I(N__16564));
    Odrv12 I__3271 (
            .O(N__16567),
            .I(DEBUG_c_5_c));
    Odrv12 I__3270 (
            .O(N__16564),
            .I(DEBUG_c_5_c));
    InMux I__3269 (
            .O(N__16559),
            .I(N__16556));
    LocalMux I__3268 (
            .O(N__16556),
            .I(\tvp_video_buffer.BUFFER_0_7 ));
    InMux I__3267 (
            .O(N__16553),
            .I(N__16548));
    InMux I__3266 (
            .O(N__16552),
            .I(N__16545));
    InMux I__3265 (
            .O(N__16551),
            .I(N__16541));
    LocalMux I__3264 (
            .O(N__16548),
            .I(N__16536));
    LocalMux I__3263 (
            .O(N__16545),
            .I(N__16536));
    InMux I__3262 (
            .O(N__16544),
            .I(N__16533));
    LocalMux I__3261 (
            .O(N__16541),
            .I(\transmit_module.TX_ADDR_0 ));
    Odrv12 I__3260 (
            .O(N__16536),
            .I(\transmit_module.TX_ADDR_0 ));
    LocalMux I__3259 (
            .O(N__16533),
            .I(\transmit_module.TX_ADDR_0 ));
    InMux I__3258 (
            .O(N__16526),
            .I(N__16523));
    LocalMux I__3257 (
            .O(N__16523),
            .I(\transmit_module.n132 ));
    CascadeMux I__3256 (
            .O(N__16520),
            .I(N__16517));
    InMux I__3255 (
            .O(N__16517),
            .I(N__16514));
    LocalMux I__3254 (
            .O(N__16514),
            .I(\transmit_module.n131 ));
    InMux I__3253 (
            .O(N__16511),
            .I(\transmit_module.n3104 ));
    InMux I__3252 (
            .O(N__16508),
            .I(\transmit_module.n3105 ));
    InMux I__3251 (
            .O(N__16505),
            .I(N__16502));
    LocalMux I__3250 (
            .O(N__16502),
            .I(N__16498));
    InMux I__3249 (
            .O(N__16501),
            .I(N__16495));
    Span4Mux_v I__3248 (
            .O(N__16498),
            .I(N__16488));
    LocalMux I__3247 (
            .O(N__16495),
            .I(N__16488));
    InMux I__3246 (
            .O(N__16494),
            .I(N__16485));
    CascadeMux I__3245 (
            .O(N__16493),
            .I(N__16482));
    Sp12to4 I__3244 (
            .O(N__16488),
            .I(N__16477));
    LocalMux I__3243 (
            .O(N__16485),
            .I(N__16477));
    InMux I__3242 (
            .O(N__16482),
            .I(N__16474));
    Odrv12 I__3241 (
            .O(N__16477),
            .I(\transmit_module.TX_ADDR_3 ));
    LocalMux I__3240 (
            .O(N__16474),
            .I(\transmit_module.TX_ADDR_3 ));
    InMux I__3239 (
            .O(N__16469),
            .I(N__16466));
    LocalMux I__3238 (
            .O(N__16466),
            .I(N__16463));
    Span4Mux_v I__3237 (
            .O(N__16463),
            .I(N__16460));
    Odrv4 I__3236 (
            .O(N__16460),
            .I(\transmit_module.n129 ));
    InMux I__3235 (
            .O(N__16457),
            .I(\transmit_module.n3106 ));
    InMux I__3234 (
            .O(N__16454),
            .I(\transmit_module.n3107 ));
    InMux I__3233 (
            .O(N__16451),
            .I(N__16448));
    LocalMux I__3232 (
            .O(N__16448),
            .I(\transmit_module.n127 ));
    InMux I__3231 (
            .O(N__16445),
            .I(\transmit_module.n3108 ));
    InMux I__3230 (
            .O(N__16442),
            .I(\transmit_module.n3109 ));
    InMux I__3229 (
            .O(N__16439),
            .I(N__16436));
    LocalMux I__3228 (
            .O(N__16436),
            .I(N__16433));
    Span4Mux_v I__3227 (
            .O(N__16433),
            .I(N__16430));
    Odrv4 I__3226 (
            .O(N__16430),
            .I(\transmit_module.ADDR_Y_COMPONENT_0 ));
    InMux I__3225 (
            .O(N__16427),
            .I(N__16424));
    LocalMux I__3224 (
            .O(N__16424),
            .I(N__16418));
    InMux I__3223 (
            .O(N__16423),
            .I(N__16415));
    InMux I__3222 (
            .O(N__16422),
            .I(N__16410));
    InMux I__3221 (
            .O(N__16421),
            .I(N__16410));
    Odrv4 I__3220 (
            .O(N__16418),
            .I(\transmit_module.old_VGA_HS ));
    LocalMux I__3219 (
            .O(N__16415),
            .I(\transmit_module.old_VGA_HS ));
    LocalMux I__3218 (
            .O(N__16410),
            .I(\transmit_module.old_VGA_HS ));
    InMux I__3217 (
            .O(N__16403),
            .I(N__16400));
    LocalMux I__3216 (
            .O(N__16400),
            .I(N__16394));
    InMux I__3215 (
            .O(N__16399),
            .I(N__16391));
    InMux I__3214 (
            .O(N__16398),
            .I(N__16386));
    InMux I__3213 (
            .O(N__16397),
            .I(N__16386));
    Odrv4 I__3212 (
            .O(N__16394),
            .I(\transmit_module.VGA_VISIBLE_Y ));
    LocalMux I__3211 (
            .O(N__16391),
            .I(\transmit_module.VGA_VISIBLE_Y ));
    LocalMux I__3210 (
            .O(N__16386),
            .I(\transmit_module.VGA_VISIBLE_Y ));
    IoInMux I__3209 (
            .O(N__16379),
            .I(N__16376));
    LocalMux I__3208 (
            .O(N__16376),
            .I(N__16373));
    Span4Mux_s3_h I__3207 (
            .O(N__16373),
            .I(N__16370));
    Sp12to4 I__3206 (
            .O(N__16370),
            .I(N__16366));
    InMux I__3205 (
            .O(N__16369),
            .I(N__16363));
    Span12Mux_v I__3204 (
            .O(N__16366),
            .I(N__16356));
    LocalMux I__3203 (
            .O(N__16363),
            .I(N__16353));
    InMux I__3202 (
            .O(N__16362),
            .I(N__16348));
    InMux I__3201 (
            .O(N__16361),
            .I(N__16348));
    InMux I__3200 (
            .O(N__16360),
            .I(N__16343));
    InMux I__3199 (
            .O(N__16359),
            .I(N__16343));
    Odrv12 I__3198 (
            .O(N__16356),
            .I(ADV_HSYNC_c));
    Odrv4 I__3197 (
            .O(N__16353),
            .I(ADV_HSYNC_c));
    LocalMux I__3196 (
            .O(N__16348),
            .I(ADV_HSYNC_c));
    LocalMux I__3195 (
            .O(N__16343),
            .I(ADV_HSYNC_c));
    InMux I__3194 (
            .O(N__16334),
            .I(N__16331));
    LocalMux I__3193 (
            .O(N__16331),
            .I(N__16328));
    Odrv12 I__3192 (
            .O(N__16328),
            .I(\transmit_module.n137 ));
    CascadeMux I__3191 (
            .O(N__16325),
            .I(N__16322));
    CascadeBuf I__3190 (
            .O(N__16322),
            .I(N__16318));
    CascadeMux I__3189 (
            .O(N__16321),
            .I(N__16315));
    CascadeMux I__3188 (
            .O(N__16318),
            .I(N__16312));
    CascadeBuf I__3187 (
            .O(N__16315),
            .I(N__16309));
    CascadeBuf I__3186 (
            .O(N__16312),
            .I(N__16306));
    CascadeMux I__3185 (
            .O(N__16309),
            .I(N__16303));
    CascadeMux I__3184 (
            .O(N__16306),
            .I(N__16300));
    CascadeBuf I__3183 (
            .O(N__16303),
            .I(N__16297));
    CascadeBuf I__3182 (
            .O(N__16300),
            .I(N__16294));
    CascadeMux I__3181 (
            .O(N__16297),
            .I(N__16291));
    CascadeMux I__3180 (
            .O(N__16294),
            .I(N__16288));
    CascadeBuf I__3179 (
            .O(N__16291),
            .I(N__16285));
    CascadeBuf I__3178 (
            .O(N__16288),
            .I(N__16282));
    CascadeMux I__3177 (
            .O(N__16285),
            .I(N__16279));
    CascadeMux I__3176 (
            .O(N__16282),
            .I(N__16276));
    CascadeBuf I__3175 (
            .O(N__16279),
            .I(N__16273));
    CascadeBuf I__3174 (
            .O(N__16276),
            .I(N__16270));
    CascadeMux I__3173 (
            .O(N__16273),
            .I(N__16267));
    CascadeMux I__3172 (
            .O(N__16270),
            .I(N__16264));
    CascadeBuf I__3171 (
            .O(N__16267),
            .I(N__16261));
    CascadeBuf I__3170 (
            .O(N__16264),
            .I(N__16258));
    CascadeMux I__3169 (
            .O(N__16261),
            .I(N__16255));
    CascadeMux I__3168 (
            .O(N__16258),
            .I(N__16252));
    CascadeBuf I__3167 (
            .O(N__16255),
            .I(N__16249));
    CascadeBuf I__3166 (
            .O(N__16252),
            .I(N__16246));
    CascadeMux I__3165 (
            .O(N__16249),
            .I(N__16243));
    CascadeMux I__3164 (
            .O(N__16246),
            .I(N__16240));
    CascadeBuf I__3163 (
            .O(N__16243),
            .I(N__16237));
    CascadeBuf I__3162 (
            .O(N__16240),
            .I(N__16234));
    CascadeMux I__3161 (
            .O(N__16237),
            .I(N__16231));
    CascadeMux I__3160 (
            .O(N__16234),
            .I(N__16228));
    CascadeBuf I__3159 (
            .O(N__16231),
            .I(N__16225));
    CascadeBuf I__3158 (
            .O(N__16228),
            .I(N__16222));
    CascadeMux I__3157 (
            .O(N__16225),
            .I(N__16219));
    CascadeMux I__3156 (
            .O(N__16222),
            .I(N__16216));
    CascadeBuf I__3155 (
            .O(N__16219),
            .I(N__16213));
    CascadeBuf I__3154 (
            .O(N__16216),
            .I(N__16210));
    CascadeMux I__3153 (
            .O(N__16213),
            .I(N__16207));
    CascadeMux I__3152 (
            .O(N__16210),
            .I(N__16204));
    CascadeBuf I__3151 (
            .O(N__16207),
            .I(N__16201));
    CascadeBuf I__3150 (
            .O(N__16204),
            .I(N__16198));
    CascadeMux I__3149 (
            .O(N__16201),
            .I(N__16195));
    CascadeMux I__3148 (
            .O(N__16198),
            .I(N__16192));
    CascadeBuf I__3147 (
            .O(N__16195),
            .I(N__16189));
    CascadeBuf I__3146 (
            .O(N__16192),
            .I(N__16186));
    CascadeMux I__3145 (
            .O(N__16189),
            .I(N__16183));
    CascadeMux I__3144 (
            .O(N__16186),
            .I(N__16180));
    CascadeBuf I__3143 (
            .O(N__16183),
            .I(N__16177));
    CascadeBuf I__3142 (
            .O(N__16180),
            .I(N__16174));
    CascadeMux I__3141 (
            .O(N__16177),
            .I(N__16171));
    CascadeMux I__3140 (
            .O(N__16174),
            .I(N__16168));
    CascadeBuf I__3139 (
            .O(N__16171),
            .I(N__16165));
    CascadeBuf I__3138 (
            .O(N__16168),
            .I(N__16162));
    CascadeMux I__3137 (
            .O(N__16165),
            .I(N__16159));
    CascadeMux I__3136 (
            .O(N__16162),
            .I(N__16156));
    CascadeBuf I__3135 (
            .O(N__16159),
            .I(N__16153));
    CascadeBuf I__3134 (
            .O(N__16156),
            .I(N__16150));
    CascadeMux I__3133 (
            .O(N__16153),
            .I(N__16147));
    CascadeMux I__3132 (
            .O(N__16150),
            .I(N__16144));
    CascadeBuf I__3131 (
            .O(N__16147),
            .I(N__16141));
    InMux I__3130 (
            .O(N__16144),
            .I(N__16138));
    CascadeMux I__3129 (
            .O(N__16141),
            .I(N__16135));
    LocalMux I__3128 (
            .O(N__16138),
            .I(N__16132));
    InMux I__3127 (
            .O(N__16135),
            .I(N__16129));
    Span4Mux_v I__3126 (
            .O(N__16132),
            .I(N__16126));
    LocalMux I__3125 (
            .O(N__16129),
            .I(N__16123));
    Span4Mux_v I__3124 (
            .O(N__16126),
            .I(N__16120));
    Span4Mux_v I__3123 (
            .O(N__16123),
            .I(N__16117));
    Span4Mux_v I__3122 (
            .O(N__16120),
            .I(N__16114));
    Span4Mux_v I__3121 (
            .O(N__16117),
            .I(N__16111));
    Span4Mux_h I__3120 (
            .O(N__16114),
            .I(N__16108));
    Span4Mux_v I__3119 (
            .O(N__16111),
            .I(N__16105));
    Span4Mux_h I__3118 (
            .O(N__16108),
            .I(N__16100));
    Span4Mux_h I__3117 (
            .O(N__16105),
            .I(N__16100));
    Odrv4 I__3116 (
            .O(N__16100),
            .I(n18));
    InMux I__3115 (
            .O(N__16097),
            .I(N__16094));
    LocalMux I__3114 (
            .O(N__16094),
            .I(N__16090));
    InMux I__3113 (
            .O(N__16093),
            .I(N__16087));
    Odrv12 I__3112 (
            .O(N__16090),
            .I(\transmit_module.n116 ));
    LocalMux I__3111 (
            .O(N__16087),
            .I(\transmit_module.n116 ));
    InMux I__3110 (
            .O(N__16082),
            .I(N__16078));
    InMux I__3109 (
            .O(N__16081),
            .I(N__16075));
    LocalMux I__3108 (
            .O(N__16078),
            .I(N__16072));
    LocalMux I__3107 (
            .O(N__16075),
            .I(\transmit_module.n147 ));
    Odrv12 I__3106 (
            .O(N__16072),
            .I(\transmit_module.n147 ));
    CascadeMux I__3105 (
            .O(N__16067),
            .I(N__16063));
    CascadeMux I__3104 (
            .O(N__16066),
            .I(N__16060));
    CascadeBuf I__3103 (
            .O(N__16063),
            .I(N__16057));
    CascadeBuf I__3102 (
            .O(N__16060),
            .I(N__16054));
    CascadeMux I__3101 (
            .O(N__16057),
            .I(N__16051));
    CascadeMux I__3100 (
            .O(N__16054),
            .I(N__16048));
    CascadeBuf I__3099 (
            .O(N__16051),
            .I(N__16045));
    CascadeBuf I__3098 (
            .O(N__16048),
            .I(N__16042));
    CascadeMux I__3097 (
            .O(N__16045),
            .I(N__16039));
    CascadeMux I__3096 (
            .O(N__16042),
            .I(N__16036));
    CascadeBuf I__3095 (
            .O(N__16039),
            .I(N__16033));
    CascadeBuf I__3094 (
            .O(N__16036),
            .I(N__16030));
    CascadeMux I__3093 (
            .O(N__16033),
            .I(N__16027));
    CascadeMux I__3092 (
            .O(N__16030),
            .I(N__16024));
    CascadeBuf I__3091 (
            .O(N__16027),
            .I(N__16021));
    CascadeBuf I__3090 (
            .O(N__16024),
            .I(N__16018));
    CascadeMux I__3089 (
            .O(N__16021),
            .I(N__16015));
    CascadeMux I__3088 (
            .O(N__16018),
            .I(N__16012));
    CascadeBuf I__3087 (
            .O(N__16015),
            .I(N__16009));
    CascadeBuf I__3086 (
            .O(N__16012),
            .I(N__16006));
    CascadeMux I__3085 (
            .O(N__16009),
            .I(N__16003));
    CascadeMux I__3084 (
            .O(N__16006),
            .I(N__16000));
    CascadeBuf I__3083 (
            .O(N__16003),
            .I(N__15997));
    CascadeBuf I__3082 (
            .O(N__16000),
            .I(N__15994));
    CascadeMux I__3081 (
            .O(N__15997),
            .I(N__15991));
    CascadeMux I__3080 (
            .O(N__15994),
            .I(N__15988));
    CascadeBuf I__3079 (
            .O(N__15991),
            .I(N__15985));
    CascadeBuf I__3078 (
            .O(N__15988),
            .I(N__15982));
    CascadeMux I__3077 (
            .O(N__15985),
            .I(N__15979));
    CascadeMux I__3076 (
            .O(N__15982),
            .I(N__15976));
    CascadeBuf I__3075 (
            .O(N__15979),
            .I(N__15973));
    CascadeBuf I__3074 (
            .O(N__15976),
            .I(N__15970));
    CascadeMux I__3073 (
            .O(N__15973),
            .I(N__15967));
    CascadeMux I__3072 (
            .O(N__15970),
            .I(N__15964));
    CascadeBuf I__3071 (
            .O(N__15967),
            .I(N__15961));
    CascadeBuf I__3070 (
            .O(N__15964),
            .I(N__15958));
    CascadeMux I__3069 (
            .O(N__15961),
            .I(N__15955));
    CascadeMux I__3068 (
            .O(N__15958),
            .I(N__15952));
    CascadeBuf I__3067 (
            .O(N__15955),
            .I(N__15949));
    CascadeBuf I__3066 (
            .O(N__15952),
            .I(N__15946));
    CascadeMux I__3065 (
            .O(N__15949),
            .I(N__15943));
    CascadeMux I__3064 (
            .O(N__15946),
            .I(N__15940));
    CascadeBuf I__3063 (
            .O(N__15943),
            .I(N__15937));
    CascadeBuf I__3062 (
            .O(N__15940),
            .I(N__15934));
    CascadeMux I__3061 (
            .O(N__15937),
            .I(N__15931));
    CascadeMux I__3060 (
            .O(N__15934),
            .I(N__15928));
    CascadeBuf I__3059 (
            .O(N__15931),
            .I(N__15925));
    CascadeBuf I__3058 (
            .O(N__15928),
            .I(N__15922));
    CascadeMux I__3057 (
            .O(N__15925),
            .I(N__15919));
    CascadeMux I__3056 (
            .O(N__15922),
            .I(N__15916));
    CascadeBuf I__3055 (
            .O(N__15919),
            .I(N__15913));
    CascadeBuf I__3054 (
            .O(N__15916),
            .I(N__15910));
    CascadeMux I__3053 (
            .O(N__15913),
            .I(N__15907));
    CascadeMux I__3052 (
            .O(N__15910),
            .I(N__15904));
    CascadeBuf I__3051 (
            .O(N__15907),
            .I(N__15901));
    CascadeBuf I__3050 (
            .O(N__15904),
            .I(N__15898));
    CascadeMux I__3049 (
            .O(N__15901),
            .I(N__15895));
    CascadeMux I__3048 (
            .O(N__15898),
            .I(N__15892));
    CascadeBuf I__3047 (
            .O(N__15895),
            .I(N__15889));
    CascadeBuf I__3046 (
            .O(N__15892),
            .I(N__15886));
    CascadeMux I__3045 (
            .O(N__15889),
            .I(N__15883));
    CascadeMux I__3044 (
            .O(N__15886),
            .I(N__15880));
    InMux I__3043 (
            .O(N__15883),
            .I(N__15877));
    InMux I__3042 (
            .O(N__15880),
            .I(N__15874));
    LocalMux I__3041 (
            .O(N__15877),
            .I(N__15871));
    LocalMux I__3040 (
            .O(N__15874),
            .I(N__15868));
    Span4Mux_s2_v I__3039 (
            .O(N__15871),
            .I(N__15865));
    Span12Mux_s11_h I__3038 (
            .O(N__15868),
            .I(N__15862));
    Sp12to4 I__3037 (
            .O(N__15865),
            .I(N__15859));
    Span12Mux_v I__3036 (
            .O(N__15862),
            .I(N__15854));
    Span12Mux_v I__3035 (
            .O(N__15859),
            .I(N__15854));
    Odrv12 I__3034 (
            .O(N__15854),
            .I(n28));
    InMux I__3033 (
            .O(N__15851),
            .I(N__15847));
    InMux I__3032 (
            .O(N__15850),
            .I(N__15844));
    LocalMux I__3031 (
            .O(N__15847),
            .I(N__15841));
    LocalMux I__3030 (
            .O(N__15844),
            .I(N__15838));
    Span12Mux_v I__3029 (
            .O(N__15841),
            .I(N__15833));
    Span12Mux_s5_v I__3028 (
            .O(N__15838),
            .I(N__15833));
    Odrv12 I__3027 (
            .O(N__15833),
            .I(\transmit_module.n115 ));
    InMux I__3026 (
            .O(N__15830),
            .I(N__15827));
    LocalMux I__3025 (
            .O(N__15827),
            .I(N__15823));
    InMux I__3024 (
            .O(N__15826),
            .I(N__15820));
    Span12Mux_s10_v I__3023 (
            .O(N__15823),
            .I(N__15817));
    LocalMux I__3022 (
            .O(N__15820),
            .I(\transmit_module.n146 ));
    Odrv12 I__3021 (
            .O(N__15817),
            .I(\transmit_module.n146 ));
    CascadeMux I__3020 (
            .O(N__15812),
            .I(N__15808));
    CascadeMux I__3019 (
            .O(N__15811),
            .I(N__15805));
    CascadeBuf I__3018 (
            .O(N__15808),
            .I(N__15802));
    CascadeBuf I__3017 (
            .O(N__15805),
            .I(N__15799));
    CascadeMux I__3016 (
            .O(N__15802),
            .I(N__15796));
    CascadeMux I__3015 (
            .O(N__15799),
            .I(N__15793));
    CascadeBuf I__3014 (
            .O(N__15796),
            .I(N__15790));
    CascadeBuf I__3013 (
            .O(N__15793),
            .I(N__15787));
    CascadeMux I__3012 (
            .O(N__15790),
            .I(N__15784));
    CascadeMux I__3011 (
            .O(N__15787),
            .I(N__15781));
    CascadeBuf I__3010 (
            .O(N__15784),
            .I(N__15778));
    CascadeBuf I__3009 (
            .O(N__15781),
            .I(N__15775));
    CascadeMux I__3008 (
            .O(N__15778),
            .I(N__15772));
    CascadeMux I__3007 (
            .O(N__15775),
            .I(N__15769));
    CascadeBuf I__3006 (
            .O(N__15772),
            .I(N__15766));
    CascadeBuf I__3005 (
            .O(N__15769),
            .I(N__15763));
    CascadeMux I__3004 (
            .O(N__15766),
            .I(N__15760));
    CascadeMux I__3003 (
            .O(N__15763),
            .I(N__15757));
    CascadeBuf I__3002 (
            .O(N__15760),
            .I(N__15754));
    CascadeBuf I__3001 (
            .O(N__15757),
            .I(N__15751));
    CascadeMux I__3000 (
            .O(N__15754),
            .I(N__15748));
    CascadeMux I__2999 (
            .O(N__15751),
            .I(N__15745));
    CascadeBuf I__2998 (
            .O(N__15748),
            .I(N__15742));
    CascadeBuf I__2997 (
            .O(N__15745),
            .I(N__15739));
    CascadeMux I__2996 (
            .O(N__15742),
            .I(N__15736));
    CascadeMux I__2995 (
            .O(N__15739),
            .I(N__15733));
    CascadeBuf I__2994 (
            .O(N__15736),
            .I(N__15730));
    CascadeBuf I__2993 (
            .O(N__15733),
            .I(N__15727));
    CascadeMux I__2992 (
            .O(N__15730),
            .I(N__15724));
    CascadeMux I__2991 (
            .O(N__15727),
            .I(N__15721));
    CascadeBuf I__2990 (
            .O(N__15724),
            .I(N__15718));
    CascadeBuf I__2989 (
            .O(N__15721),
            .I(N__15715));
    CascadeMux I__2988 (
            .O(N__15718),
            .I(N__15712));
    CascadeMux I__2987 (
            .O(N__15715),
            .I(N__15709));
    CascadeBuf I__2986 (
            .O(N__15712),
            .I(N__15706));
    CascadeBuf I__2985 (
            .O(N__15709),
            .I(N__15703));
    CascadeMux I__2984 (
            .O(N__15706),
            .I(N__15700));
    CascadeMux I__2983 (
            .O(N__15703),
            .I(N__15697));
    CascadeBuf I__2982 (
            .O(N__15700),
            .I(N__15694));
    CascadeBuf I__2981 (
            .O(N__15697),
            .I(N__15691));
    CascadeMux I__2980 (
            .O(N__15694),
            .I(N__15688));
    CascadeMux I__2979 (
            .O(N__15691),
            .I(N__15685));
    CascadeBuf I__2978 (
            .O(N__15688),
            .I(N__15682));
    CascadeBuf I__2977 (
            .O(N__15685),
            .I(N__15679));
    CascadeMux I__2976 (
            .O(N__15682),
            .I(N__15676));
    CascadeMux I__2975 (
            .O(N__15679),
            .I(N__15673));
    CascadeBuf I__2974 (
            .O(N__15676),
            .I(N__15670));
    CascadeBuf I__2973 (
            .O(N__15673),
            .I(N__15667));
    CascadeMux I__2972 (
            .O(N__15670),
            .I(N__15664));
    CascadeMux I__2971 (
            .O(N__15667),
            .I(N__15661));
    CascadeBuf I__2970 (
            .O(N__15664),
            .I(N__15658));
    CascadeBuf I__2969 (
            .O(N__15661),
            .I(N__15655));
    CascadeMux I__2968 (
            .O(N__15658),
            .I(N__15652));
    CascadeMux I__2967 (
            .O(N__15655),
            .I(N__15649));
    CascadeBuf I__2966 (
            .O(N__15652),
            .I(N__15646));
    CascadeBuf I__2965 (
            .O(N__15649),
            .I(N__15643));
    CascadeMux I__2964 (
            .O(N__15646),
            .I(N__15640));
    CascadeMux I__2963 (
            .O(N__15643),
            .I(N__15637));
    CascadeBuf I__2962 (
            .O(N__15640),
            .I(N__15634));
    CascadeBuf I__2961 (
            .O(N__15637),
            .I(N__15631));
    CascadeMux I__2960 (
            .O(N__15634),
            .I(N__15628));
    CascadeMux I__2959 (
            .O(N__15631),
            .I(N__15625));
    InMux I__2958 (
            .O(N__15628),
            .I(N__15622));
    InMux I__2957 (
            .O(N__15625),
            .I(N__15619));
    LocalMux I__2956 (
            .O(N__15622),
            .I(N__15616));
    LocalMux I__2955 (
            .O(N__15619),
            .I(N__15613));
    Span12Mux_s9_h I__2954 (
            .O(N__15616),
            .I(N__15610));
    Span4Mux_h I__2953 (
            .O(N__15613),
            .I(N__15607));
    Odrv12 I__2952 (
            .O(N__15610),
            .I(n27));
    Odrv4 I__2951 (
            .O(N__15607),
            .I(n27));
    InMux I__2950 (
            .O(N__15602),
            .I(N__15598));
    IoInMux I__2949 (
            .O(N__15601),
            .I(N__15595));
    LocalMux I__2948 (
            .O(N__15598),
            .I(N__15592));
    LocalMux I__2947 (
            .O(N__15595),
            .I(N__15589));
    Span4Mux_h I__2946 (
            .O(N__15592),
            .I(N__15586));
    Span12Mux_s11_h I__2945 (
            .O(N__15589),
            .I(N__15583));
    Span4Mux_v I__2944 (
            .O(N__15586),
            .I(N__15580));
    Odrv12 I__2943 (
            .O(N__15583),
            .I(DEBUG_c_3_c));
    Odrv4 I__2942 (
            .O(N__15580),
            .I(DEBUG_c_3_c));
    IoInMux I__2941 (
            .O(N__15575),
            .I(N__15572));
    LocalMux I__2940 (
            .O(N__15572),
            .I(N__15569));
    IoSpan4Mux I__2939 (
            .O(N__15569),
            .I(N__15566));
    Span4Mux_s0_h I__2938 (
            .O(N__15566),
            .I(N__15562));
    InMux I__2937 (
            .O(N__15565),
            .I(N__15559));
    Sp12to4 I__2936 (
            .O(N__15562),
            .I(N__15556));
    LocalMux I__2935 (
            .O(N__15559),
            .I(N__15553));
    Span12Mux_s11_h I__2934 (
            .O(N__15556),
            .I(N__15550));
    Span4Mux_h I__2933 (
            .O(N__15553),
            .I(N__15547));
    Span12Mux_v I__2932 (
            .O(N__15550),
            .I(N__15544));
    Span4Mux_v I__2931 (
            .O(N__15547),
            .I(N__15541));
    Odrv12 I__2930 (
            .O(N__15544),
            .I(DEBUG_c_4_c));
    Odrv4 I__2929 (
            .O(N__15541),
            .I(DEBUG_c_4_c));
    CascadeMux I__2928 (
            .O(N__15536),
            .I(N__15533));
    InMux I__2927 (
            .O(N__15533),
            .I(N__15529));
    InMux I__2926 (
            .O(N__15532),
            .I(N__15524));
    LocalMux I__2925 (
            .O(N__15529),
            .I(N__15521));
    InMux I__2924 (
            .O(N__15528),
            .I(N__15518));
    InMux I__2923 (
            .O(N__15527),
            .I(N__15515));
    LocalMux I__2922 (
            .O(N__15524),
            .I(N__15510));
    Span4Mux_v I__2921 (
            .O(N__15521),
            .I(N__15510));
    LocalMux I__2920 (
            .O(N__15518),
            .I(\transmit_module.video_signal_controller.VGA_Y_4 ));
    LocalMux I__2919 (
            .O(N__15515),
            .I(\transmit_module.video_signal_controller.VGA_Y_4 ));
    Odrv4 I__2918 (
            .O(N__15510),
            .I(\transmit_module.video_signal_controller.VGA_Y_4 ));
    InMux I__2917 (
            .O(N__15503),
            .I(N__15500));
    LocalMux I__2916 (
            .O(N__15500),
            .I(\transmit_module.video_signal_controller.n3628 ));
    InMux I__2915 (
            .O(N__15497),
            .I(N__15493));
    CascadeMux I__2914 (
            .O(N__15496),
            .I(N__15489));
    LocalMux I__2913 (
            .O(N__15493),
            .I(N__15485));
    InMux I__2912 (
            .O(N__15492),
            .I(N__15482));
    InMux I__2911 (
            .O(N__15489),
            .I(N__15479));
    InMux I__2910 (
            .O(N__15488),
            .I(N__15476));
    Span4Mux_v I__2909 (
            .O(N__15485),
            .I(N__15469));
    LocalMux I__2908 (
            .O(N__15482),
            .I(N__15469));
    LocalMux I__2907 (
            .O(N__15479),
            .I(N__15469));
    LocalMux I__2906 (
            .O(N__15476),
            .I(\transmit_module.video_signal_controller.VGA_Y_9 ));
    Odrv4 I__2905 (
            .O(N__15469),
            .I(\transmit_module.video_signal_controller.VGA_Y_9 ));
    InMux I__2904 (
            .O(N__15464),
            .I(N__15461));
    LocalMux I__2903 (
            .O(N__15461),
            .I(N__15457));
    InMux I__2902 (
            .O(N__15460),
            .I(N__15454));
    Odrv4 I__2901 (
            .O(N__15457),
            .I(\transmit_module.video_signal_controller.n3331 ));
    LocalMux I__2900 (
            .O(N__15454),
            .I(\transmit_module.video_signal_controller.n3331 ));
    CascadeMux I__2899 (
            .O(N__15449),
            .I(\transmit_module.video_signal_controller.n7_adj_618_cascade_ ));
    InMux I__2898 (
            .O(N__15446),
            .I(N__15443));
    LocalMux I__2897 (
            .O(N__15443),
            .I(N__15440));
    Odrv4 I__2896 (
            .O(N__15440),
            .I(\transmit_module.video_signal_controller.n3622 ));
    CascadeMux I__2895 (
            .O(N__15437),
            .I(\transmit_module.video_signal_controller.VGA_VISIBLE_N_580_cascade_ ));
    InMux I__2894 (
            .O(N__15434),
            .I(N__15431));
    LocalMux I__2893 (
            .O(N__15431),
            .I(N__15426));
    InMux I__2892 (
            .O(N__15430),
            .I(N__15423));
    InMux I__2891 (
            .O(N__15429),
            .I(N__15420));
    Span4Mux_v I__2890 (
            .O(N__15426),
            .I(N__15415));
    LocalMux I__2889 (
            .O(N__15423),
            .I(N__15415));
    LocalMux I__2888 (
            .O(N__15420),
            .I(\transmit_module.video_signal_controller.VGA_Y_10 ));
    Odrv4 I__2887 (
            .O(N__15415),
            .I(\transmit_module.video_signal_controller.VGA_Y_10 ));
    InMux I__2886 (
            .O(N__15410),
            .I(N__15407));
    LocalMux I__2885 (
            .O(N__15407),
            .I(N__15404));
    Odrv4 I__2884 (
            .O(N__15404),
            .I(\transmit_module.video_signal_controller.n3477 ));
    CascadeMux I__2883 (
            .O(N__15401),
            .I(N__15398));
    InMux I__2882 (
            .O(N__15398),
            .I(N__15395));
    LocalMux I__2881 (
            .O(N__15395),
            .I(N__15392));
    Odrv4 I__2880 (
            .O(N__15392),
            .I(\transmit_module.video_signal_controller.n16 ));
    InMux I__2879 (
            .O(N__15389),
            .I(N__15386));
    LocalMux I__2878 (
            .O(N__15386),
            .I(N__15382));
    InMux I__2877 (
            .O(N__15385),
            .I(N__15378));
    Span4Mux_v I__2876 (
            .O(N__15382),
            .I(N__15374));
    InMux I__2875 (
            .O(N__15381),
            .I(N__15371));
    LocalMux I__2874 (
            .O(N__15378),
            .I(N__15368));
    InMux I__2873 (
            .O(N__15377),
            .I(N__15365));
    Odrv4 I__2872 (
            .O(N__15374),
            .I(\transmit_module.video_signal_controller.VGA_Y_2 ));
    LocalMux I__2871 (
            .O(N__15371),
            .I(\transmit_module.video_signal_controller.VGA_Y_2 ));
    Odrv12 I__2870 (
            .O(N__15368),
            .I(\transmit_module.video_signal_controller.VGA_Y_2 ));
    LocalMux I__2869 (
            .O(N__15365),
            .I(\transmit_module.video_signal_controller.VGA_Y_2 ));
    InMux I__2868 (
            .O(N__15356),
            .I(N__15353));
    LocalMux I__2867 (
            .O(N__15353),
            .I(N__15347));
    InMux I__2866 (
            .O(N__15352),
            .I(N__15342));
    InMux I__2865 (
            .O(N__15351),
            .I(N__15342));
    InMux I__2864 (
            .O(N__15350),
            .I(N__15339));
    Span4Mux_h I__2863 (
            .O(N__15347),
            .I(N__15334));
    LocalMux I__2862 (
            .O(N__15342),
            .I(N__15334));
    LocalMux I__2861 (
            .O(N__15339),
            .I(\transmit_module.video_signal_controller.VGA_X_8 ));
    Odrv4 I__2860 (
            .O(N__15334),
            .I(\transmit_module.video_signal_controller.VGA_X_8 ));
    InMux I__2859 (
            .O(N__15329),
            .I(N__15326));
    LocalMux I__2858 (
            .O(N__15326),
            .I(N__15323));
    Odrv4 I__2857 (
            .O(N__15323),
            .I(\transmit_module.video_signal_controller.n3471 ));
    CascadeMux I__2856 (
            .O(N__15320),
            .I(N__15317));
    InMux I__2855 (
            .O(N__15317),
            .I(N__15314));
    LocalMux I__2854 (
            .O(N__15314),
            .I(N__15311));
    Odrv4 I__2853 (
            .O(N__15311),
            .I(\transmit_module.video_signal_controller.n4_adj_617 ));
    InMux I__2852 (
            .O(N__15308),
            .I(N__15305));
    LocalMux I__2851 (
            .O(N__15305),
            .I(N__15301));
    InMux I__2850 (
            .O(N__15304),
            .I(N__15296));
    Span4Mux_h I__2849 (
            .O(N__15301),
            .I(N__15293));
    InMux I__2848 (
            .O(N__15300),
            .I(N__15290));
    InMux I__2847 (
            .O(N__15299),
            .I(N__15287));
    LocalMux I__2846 (
            .O(N__15296),
            .I(N__15284));
    Odrv4 I__2845 (
            .O(N__15293),
            .I(\transmit_module.video_signal_controller.VGA_X_6 ));
    LocalMux I__2844 (
            .O(N__15290),
            .I(\transmit_module.video_signal_controller.VGA_X_6 ));
    LocalMux I__2843 (
            .O(N__15287),
            .I(\transmit_module.video_signal_controller.VGA_X_6 ));
    Odrv4 I__2842 (
            .O(N__15284),
            .I(\transmit_module.video_signal_controller.VGA_X_6 ));
    InMux I__2841 (
            .O(N__15275),
            .I(N__15272));
    LocalMux I__2840 (
            .O(N__15272),
            .I(N__15269));
    Span4Mux_h I__2839 (
            .O(N__15269),
            .I(N__15265));
    InMux I__2838 (
            .O(N__15268),
            .I(N__15262));
    Odrv4 I__2837 (
            .O(N__15265),
            .I(\transmit_module.n144 ));
    LocalMux I__2836 (
            .O(N__15262),
            .I(\transmit_module.n144 ));
    CEMux I__2835 (
            .O(N__15257),
            .I(N__15245));
    CEMux I__2834 (
            .O(N__15256),
            .I(N__15241));
    CEMux I__2833 (
            .O(N__15255),
            .I(N__15237));
    CEMux I__2832 (
            .O(N__15254),
            .I(N__15234));
    CEMux I__2831 (
            .O(N__15253),
            .I(N__15231));
    CEMux I__2830 (
            .O(N__15252),
            .I(N__15228));
    CEMux I__2829 (
            .O(N__15251),
            .I(N__15225));
    CEMux I__2828 (
            .O(N__15250),
            .I(N__15222));
    CEMux I__2827 (
            .O(N__15249),
            .I(N__15216));
    CEMux I__2826 (
            .O(N__15248),
            .I(N__15213));
    LocalMux I__2825 (
            .O(N__15245),
            .I(N__15209));
    CEMux I__2824 (
            .O(N__15244),
            .I(N__15206));
    LocalMux I__2823 (
            .O(N__15241),
            .I(N__15203));
    CEMux I__2822 (
            .O(N__15240),
            .I(N__15200));
    LocalMux I__2821 (
            .O(N__15237),
            .I(N__15196));
    LocalMux I__2820 (
            .O(N__15234),
            .I(N__15191));
    LocalMux I__2819 (
            .O(N__15231),
            .I(N__15191));
    LocalMux I__2818 (
            .O(N__15228),
            .I(N__15188));
    LocalMux I__2817 (
            .O(N__15225),
            .I(N__15183));
    LocalMux I__2816 (
            .O(N__15222),
            .I(N__15183));
    CEMux I__2815 (
            .O(N__15221),
            .I(N__15180));
    CEMux I__2814 (
            .O(N__15220),
            .I(N__15177));
    CEMux I__2813 (
            .O(N__15219),
            .I(N__15174));
    LocalMux I__2812 (
            .O(N__15216),
            .I(N__15171));
    LocalMux I__2811 (
            .O(N__15213),
            .I(N__15168));
    CEMux I__2810 (
            .O(N__15212),
            .I(N__15165));
    Span4Mux_v I__2809 (
            .O(N__15209),
            .I(N__15161));
    LocalMux I__2808 (
            .O(N__15206),
            .I(N__15158));
    Span4Mux_v I__2807 (
            .O(N__15203),
            .I(N__15153));
    LocalMux I__2806 (
            .O(N__15200),
            .I(N__15153));
    CEMux I__2805 (
            .O(N__15199),
            .I(N__15150));
    Span4Mux_v I__2804 (
            .O(N__15196),
            .I(N__15147));
    Span4Mux_v I__2803 (
            .O(N__15191),
            .I(N__15142));
    Span4Mux_v I__2802 (
            .O(N__15188),
            .I(N__15142));
    Span4Mux_v I__2801 (
            .O(N__15183),
            .I(N__15135));
    LocalMux I__2800 (
            .O(N__15180),
            .I(N__15135));
    LocalMux I__2799 (
            .O(N__15177),
            .I(N__15135));
    LocalMux I__2798 (
            .O(N__15174),
            .I(N__15132));
    Span4Mux_h I__2797 (
            .O(N__15171),
            .I(N__15129));
    Span4Mux_h I__2796 (
            .O(N__15168),
            .I(N__15124));
    LocalMux I__2795 (
            .O(N__15165),
            .I(N__15124));
    CEMux I__2794 (
            .O(N__15164),
            .I(N__15121));
    Span4Mux_h I__2793 (
            .O(N__15161),
            .I(N__15112));
    Span4Mux_v I__2792 (
            .O(N__15158),
            .I(N__15112));
    Span4Mux_v I__2791 (
            .O(N__15153),
            .I(N__15112));
    LocalMux I__2790 (
            .O(N__15150),
            .I(N__15112));
    Span4Mux_h I__2789 (
            .O(N__15147),
            .I(N__15103));
    Span4Mux_v I__2788 (
            .O(N__15142),
            .I(N__15103));
    Span4Mux_h I__2787 (
            .O(N__15135),
            .I(N__15103));
    Span4Mux_v I__2786 (
            .O(N__15132),
            .I(N__15103));
    Span4Mux_v I__2785 (
            .O(N__15129),
            .I(N__15098));
    Span4Mux_h I__2784 (
            .O(N__15124),
            .I(N__15098));
    LocalMux I__2783 (
            .O(N__15121),
            .I(N__15095));
    Span4Mux_h I__2782 (
            .O(N__15112),
            .I(N__15092));
    Odrv4 I__2781 (
            .O(N__15103),
            .I(\transmit_module.n3636 ));
    Odrv4 I__2780 (
            .O(N__15098),
            .I(\transmit_module.n3636 ));
    Odrv12 I__2779 (
            .O(N__15095),
            .I(\transmit_module.n3636 ));
    Odrv4 I__2778 (
            .O(N__15092),
            .I(\transmit_module.n3636 ));
    InMux I__2777 (
            .O(N__15083),
            .I(N__15080));
    LocalMux I__2776 (
            .O(N__15080),
            .I(N__15077));
    Odrv4 I__2775 (
            .O(N__15077),
            .I(\transmit_module.video_signal_controller.n3412 ));
    InMux I__2774 (
            .O(N__15074),
            .I(N__15069));
    InMux I__2773 (
            .O(N__15073),
            .I(N__15066));
    InMux I__2772 (
            .O(N__15072),
            .I(N__15063));
    LocalMux I__2771 (
            .O(N__15069),
            .I(N__15060));
    LocalMux I__2770 (
            .O(N__15066),
            .I(\transmit_module.video_signal_controller.VGA_Y_8 ));
    LocalMux I__2769 (
            .O(N__15063),
            .I(\transmit_module.video_signal_controller.VGA_Y_8 ));
    Odrv4 I__2768 (
            .O(N__15060),
            .I(\transmit_module.video_signal_controller.VGA_Y_8 ));
    InMux I__2767 (
            .O(N__15053),
            .I(N__15049));
    InMux I__2766 (
            .O(N__15052),
            .I(N__15045));
    LocalMux I__2765 (
            .O(N__15049),
            .I(N__15042));
    InMux I__2764 (
            .O(N__15048),
            .I(N__15039));
    LocalMux I__2763 (
            .O(N__15045),
            .I(N__15036));
    Span4Mux_h I__2762 (
            .O(N__15042),
            .I(N__15033));
    LocalMux I__2761 (
            .O(N__15039),
            .I(\transmit_module.video_signal_controller.VGA_Y_7 ));
    Odrv4 I__2760 (
            .O(N__15036),
            .I(\transmit_module.video_signal_controller.VGA_Y_7 ));
    Odrv4 I__2759 (
            .O(N__15033),
            .I(\transmit_module.video_signal_controller.VGA_Y_7 ));
    InMux I__2758 (
            .O(N__15026),
            .I(N__15023));
    LocalMux I__2757 (
            .O(N__15023),
            .I(N__15020));
    Odrv4 I__2756 (
            .O(N__15020),
            .I(\transmit_module.video_signal_controller.n3626 ));
    CascadeMux I__2755 (
            .O(N__15017),
            .I(N__15013));
    InMux I__2754 (
            .O(N__15016),
            .I(N__15009));
    InMux I__2753 (
            .O(N__15013),
            .I(N__15006));
    InMux I__2752 (
            .O(N__15012),
            .I(N__15002));
    LocalMux I__2751 (
            .O(N__15009),
            .I(N__14997));
    LocalMux I__2750 (
            .O(N__15006),
            .I(N__14997));
    InMux I__2749 (
            .O(N__15005),
            .I(N__14994));
    LocalMux I__2748 (
            .O(N__15002),
            .I(\transmit_module.video_signal_controller.VGA_Y_6 ));
    Odrv4 I__2747 (
            .O(N__14997),
            .I(\transmit_module.video_signal_controller.VGA_Y_6 ));
    LocalMux I__2746 (
            .O(N__14994),
            .I(\transmit_module.video_signal_controller.VGA_Y_6 ));
    CascadeMux I__2745 (
            .O(N__14987),
            .I(\transmit_module.video_signal_controller.n3626_cascade_ ));
    InMux I__2744 (
            .O(N__14984),
            .I(N__14979));
    InMux I__2743 (
            .O(N__14983),
            .I(N__14976));
    InMux I__2742 (
            .O(N__14982),
            .I(N__14973));
    LocalMux I__2741 (
            .O(N__14979),
            .I(N__14970));
    LocalMux I__2740 (
            .O(N__14976),
            .I(\transmit_module.video_signal_controller.VGA_Y_11 ));
    LocalMux I__2739 (
            .O(N__14973),
            .I(\transmit_module.video_signal_controller.VGA_Y_11 ));
    Odrv4 I__2738 (
            .O(N__14970),
            .I(\transmit_module.video_signal_controller.VGA_Y_11 ));
    CascadeMux I__2737 (
            .O(N__14963),
            .I(\transmit_module.n137_cascade_ ));
    InMux I__2736 (
            .O(N__14960),
            .I(N__14956));
    InMux I__2735 (
            .O(N__14959),
            .I(N__14951));
    LocalMux I__2734 (
            .O(N__14956),
            .I(N__14948));
    InMux I__2733 (
            .O(N__14955),
            .I(N__14945));
    InMux I__2732 (
            .O(N__14954),
            .I(N__14942));
    LocalMux I__2731 (
            .O(N__14951),
            .I(N__14937));
    Span4Mux_v I__2730 (
            .O(N__14948),
            .I(N__14937));
    LocalMux I__2729 (
            .O(N__14945),
            .I(\transmit_module.video_signal_controller.VGA_Y_5 ));
    LocalMux I__2728 (
            .O(N__14942),
            .I(\transmit_module.video_signal_controller.VGA_Y_5 ));
    Odrv4 I__2727 (
            .O(N__14937),
            .I(\transmit_module.video_signal_controller.VGA_Y_5 ));
    InMux I__2726 (
            .O(N__14930),
            .I(N__14926));
    InMux I__2725 (
            .O(N__14929),
            .I(N__14923));
    LocalMux I__2724 (
            .O(N__14926),
            .I(N__14917));
    LocalMux I__2723 (
            .O(N__14923),
            .I(N__14917));
    InMux I__2722 (
            .O(N__14922),
            .I(N__14913));
    Span4Mux_v I__2721 (
            .O(N__14917),
            .I(N__14910));
    InMux I__2720 (
            .O(N__14916),
            .I(N__14907));
    LocalMux I__2719 (
            .O(N__14913),
            .I(\transmit_module.video_signal_controller.VGA_Y_3 ));
    Odrv4 I__2718 (
            .O(N__14910),
            .I(\transmit_module.video_signal_controller.VGA_Y_3 ));
    LocalMux I__2717 (
            .O(N__14907),
            .I(\transmit_module.video_signal_controller.VGA_Y_3 ));
    InMux I__2716 (
            .O(N__14900),
            .I(N__14897));
    LocalMux I__2715 (
            .O(N__14897),
            .I(N__14893));
    InMux I__2714 (
            .O(N__14896),
            .I(N__14888));
    Span4Mux_v I__2713 (
            .O(N__14893),
            .I(N__14885));
    InMux I__2712 (
            .O(N__14892),
            .I(N__14880));
    InMux I__2711 (
            .O(N__14891),
            .I(N__14880));
    LocalMux I__2710 (
            .O(N__14888),
            .I(\transmit_module.video_signal_controller.VGA_Y_1 ));
    Odrv4 I__2709 (
            .O(N__14885),
            .I(\transmit_module.video_signal_controller.VGA_Y_1 ));
    LocalMux I__2708 (
            .O(N__14880),
            .I(\transmit_module.video_signal_controller.VGA_Y_1 ));
    InMux I__2707 (
            .O(N__14873),
            .I(N__14869));
    InMux I__2706 (
            .O(N__14872),
            .I(N__14866));
    LocalMux I__2705 (
            .O(N__14869),
            .I(\transmit_module.video_signal_controller.VGA_Y_0 ));
    LocalMux I__2704 (
            .O(N__14866),
            .I(\transmit_module.video_signal_controller.VGA_Y_0 ));
    InMux I__2703 (
            .O(N__14861),
            .I(N__14858));
    LocalMux I__2702 (
            .O(N__14858),
            .I(N__14854));
    CascadeMux I__2701 (
            .O(N__14857),
            .I(N__14851));
    Span4Mux_v I__2700 (
            .O(N__14854),
            .I(N__14848));
    InMux I__2699 (
            .O(N__14851),
            .I(N__14845));
    Odrv4 I__2698 (
            .O(N__14848),
            .I(\transmit_module.n113 ));
    LocalMux I__2697 (
            .O(N__14845),
            .I(\transmit_module.n113 ));
    CascadeMux I__2696 (
            .O(N__14840),
            .I(\transmit_module.n142_cascade_ ));
    CascadeMux I__2695 (
            .O(N__14837),
            .I(N__14834));
    InMux I__2694 (
            .O(N__14834),
            .I(N__14831));
    LocalMux I__2693 (
            .O(N__14831),
            .I(N__14828));
    Odrv4 I__2692 (
            .O(N__14828),
            .I(\transmit_module.video_signal_controller.n45 ));
    InMux I__2691 (
            .O(N__14825),
            .I(N__14822));
    LocalMux I__2690 (
            .O(N__14822),
            .I(RX_TX_SYNC));
    InMux I__2689 (
            .O(N__14819),
            .I(N__14816));
    LocalMux I__2688 (
            .O(N__14816),
            .I(\sync_buffer.BUFFER_0_0 ));
    InMux I__2687 (
            .O(N__14813),
            .I(N__14807));
    InMux I__2686 (
            .O(N__14812),
            .I(N__14804));
    InMux I__2685 (
            .O(N__14811),
            .I(N__14800));
    InMux I__2684 (
            .O(N__14810),
            .I(N__14796));
    LocalMux I__2683 (
            .O(N__14807),
            .I(N__14791));
    LocalMux I__2682 (
            .O(N__14804),
            .I(N__14788));
    InMux I__2681 (
            .O(N__14803),
            .I(N__14785));
    LocalMux I__2680 (
            .O(N__14800),
            .I(N__14782));
    InMux I__2679 (
            .O(N__14799),
            .I(N__14779));
    LocalMux I__2678 (
            .O(N__14796),
            .I(N__14775));
    InMux I__2677 (
            .O(N__14795),
            .I(N__14772));
    InMux I__2676 (
            .O(N__14794),
            .I(N__14769));
    Span4Mux_v I__2675 (
            .O(N__14791),
            .I(N__14764));
    Span4Mux_v I__2674 (
            .O(N__14788),
            .I(N__14764));
    LocalMux I__2673 (
            .O(N__14785),
            .I(N__14757));
    Span4Mux_v I__2672 (
            .O(N__14782),
            .I(N__14757));
    LocalMux I__2671 (
            .O(N__14779),
            .I(N__14757));
    InMux I__2670 (
            .O(N__14778),
            .I(N__14754));
    Span4Mux_h I__2669 (
            .O(N__14775),
            .I(N__14747));
    LocalMux I__2668 (
            .O(N__14772),
            .I(N__14747));
    LocalMux I__2667 (
            .O(N__14769),
            .I(N__14747));
    Odrv4 I__2666 (
            .O(N__14764),
            .I(RX_ADDR_12));
    Odrv4 I__2665 (
            .O(N__14757),
            .I(RX_ADDR_12));
    LocalMux I__2664 (
            .O(N__14754),
            .I(RX_ADDR_12));
    Odrv4 I__2663 (
            .O(N__14747),
            .I(RX_ADDR_12));
    CascadeMux I__2662 (
            .O(N__14738),
            .I(N__14735));
    InMux I__2661 (
            .O(N__14735),
            .I(N__14726));
    CascadeMux I__2660 (
            .O(N__14734),
            .I(N__14723));
    CascadeMux I__2659 (
            .O(N__14733),
            .I(N__14719));
    CascadeMux I__2658 (
            .O(N__14732),
            .I(N__14715));
    CascadeMux I__2657 (
            .O(N__14731),
            .I(N__14711));
    CascadeMux I__2656 (
            .O(N__14730),
            .I(N__14708));
    CascadeMux I__2655 (
            .O(N__14729),
            .I(N__14705));
    LocalMux I__2654 (
            .O(N__14726),
            .I(N__14702));
    InMux I__2653 (
            .O(N__14723),
            .I(N__14687));
    InMux I__2652 (
            .O(N__14722),
            .I(N__14687));
    InMux I__2651 (
            .O(N__14719),
            .I(N__14687));
    InMux I__2650 (
            .O(N__14718),
            .I(N__14687));
    InMux I__2649 (
            .O(N__14715),
            .I(N__14687));
    InMux I__2648 (
            .O(N__14714),
            .I(N__14687));
    InMux I__2647 (
            .O(N__14711),
            .I(N__14687));
    InMux I__2646 (
            .O(N__14708),
            .I(N__14684));
    InMux I__2645 (
            .O(N__14705),
            .I(N__14681));
    Span4Mux_v I__2644 (
            .O(N__14702),
            .I(N__14676));
    LocalMux I__2643 (
            .O(N__14687),
            .I(N__14676));
    LocalMux I__2642 (
            .O(N__14684),
            .I(N__14670));
    LocalMux I__2641 (
            .O(N__14681),
            .I(N__14670));
    Span4Mux_v I__2640 (
            .O(N__14676),
            .I(N__14665));
    InMux I__2639 (
            .O(N__14675),
            .I(N__14662));
    Span4Mux_v I__2638 (
            .O(N__14670),
            .I(N__14659));
    CascadeMux I__2637 (
            .O(N__14669),
            .I(N__14656));
    InMux I__2636 (
            .O(N__14668),
            .I(N__14650));
    Span4Mux_v I__2635 (
            .O(N__14665),
            .I(N__14644));
    LocalMux I__2634 (
            .O(N__14662),
            .I(N__14644));
    Sp12to4 I__2633 (
            .O(N__14659),
            .I(N__14640));
    InMux I__2632 (
            .O(N__14656),
            .I(N__14637));
    InMux I__2631 (
            .O(N__14655),
            .I(N__14634));
    InMux I__2630 (
            .O(N__14654),
            .I(N__14631));
    InMux I__2629 (
            .O(N__14653),
            .I(N__14628));
    LocalMux I__2628 (
            .O(N__14650),
            .I(N__14625));
    InMux I__2627 (
            .O(N__14649),
            .I(N__14622));
    Span4Mux_v I__2626 (
            .O(N__14644),
            .I(N__14617));
    InMux I__2625 (
            .O(N__14643),
            .I(N__14614));
    Span12Mux_v I__2624 (
            .O(N__14640),
            .I(N__14603));
    LocalMux I__2623 (
            .O(N__14637),
            .I(N__14603));
    LocalMux I__2622 (
            .O(N__14634),
            .I(N__14603));
    LocalMux I__2621 (
            .O(N__14631),
            .I(N__14603));
    LocalMux I__2620 (
            .O(N__14628),
            .I(N__14603));
    Span4Mux_h I__2619 (
            .O(N__14625),
            .I(N__14600));
    LocalMux I__2618 (
            .O(N__14622),
            .I(N__14597));
    InMux I__2617 (
            .O(N__14621),
            .I(N__14594));
    InMux I__2616 (
            .O(N__14620),
            .I(N__14591));
    Odrv4 I__2615 (
            .O(N__14617),
            .I(RX_WE));
    LocalMux I__2614 (
            .O(N__14614),
            .I(RX_WE));
    Odrv12 I__2613 (
            .O(N__14603),
            .I(RX_WE));
    Odrv4 I__2612 (
            .O(N__14600),
            .I(RX_WE));
    Odrv4 I__2611 (
            .O(N__14597),
            .I(RX_WE));
    LocalMux I__2610 (
            .O(N__14594),
            .I(RX_WE));
    LocalMux I__2609 (
            .O(N__14591),
            .I(RX_WE));
    CascadeMux I__2608 (
            .O(N__14576),
            .I(N__14570));
    CascadeMux I__2607 (
            .O(N__14575),
            .I(N__14567));
    CascadeMux I__2606 (
            .O(N__14574),
            .I(N__14562));
    CascadeMux I__2605 (
            .O(N__14573),
            .I(N__14557));
    InMux I__2604 (
            .O(N__14570),
            .I(N__14554));
    InMux I__2603 (
            .O(N__14567),
            .I(N__14551));
    CascadeMux I__2602 (
            .O(N__14566),
            .I(N__14548));
    CascadeMux I__2601 (
            .O(N__14565),
            .I(N__14545));
    InMux I__2600 (
            .O(N__14562),
            .I(N__14542));
    CascadeMux I__2599 (
            .O(N__14561),
            .I(N__14539));
    CascadeMux I__2598 (
            .O(N__14560),
            .I(N__14536));
    InMux I__2597 (
            .O(N__14557),
            .I(N__14533));
    LocalMux I__2596 (
            .O(N__14554),
            .I(N__14529));
    LocalMux I__2595 (
            .O(N__14551),
            .I(N__14526));
    InMux I__2594 (
            .O(N__14548),
            .I(N__14523));
    InMux I__2593 (
            .O(N__14545),
            .I(N__14520));
    LocalMux I__2592 (
            .O(N__14542),
            .I(N__14517));
    InMux I__2591 (
            .O(N__14539),
            .I(N__14514));
    InMux I__2590 (
            .O(N__14536),
            .I(N__14511));
    LocalMux I__2589 (
            .O(N__14533),
            .I(N__14508));
    InMux I__2588 (
            .O(N__14532),
            .I(N__14505));
    Span4Mux_v I__2587 (
            .O(N__14529),
            .I(N__14500));
    Span4Mux_v I__2586 (
            .O(N__14526),
            .I(N__14500));
    LocalMux I__2585 (
            .O(N__14523),
            .I(N__14493));
    LocalMux I__2584 (
            .O(N__14520),
            .I(N__14493));
    Span4Mux_v I__2583 (
            .O(N__14517),
            .I(N__14493));
    LocalMux I__2582 (
            .O(N__14514),
            .I(N__14490));
    LocalMux I__2581 (
            .O(N__14511),
            .I(N__14485));
    Span4Mux_h I__2580 (
            .O(N__14508),
            .I(N__14485));
    LocalMux I__2579 (
            .O(N__14505),
            .I(RX_ADDR_13));
    Odrv4 I__2578 (
            .O(N__14500),
            .I(RX_ADDR_13));
    Odrv4 I__2577 (
            .O(N__14493),
            .I(RX_ADDR_13));
    Odrv4 I__2576 (
            .O(N__14490),
            .I(RX_ADDR_13));
    Odrv4 I__2575 (
            .O(N__14485),
            .I(RX_ADDR_13));
    InMux I__2574 (
            .O(N__14474),
            .I(N__14468));
    InMux I__2573 (
            .O(N__14473),
            .I(N__14464));
    InMux I__2572 (
            .O(N__14472),
            .I(N__14461));
    InMux I__2571 (
            .O(N__14471),
            .I(N__14457));
    LocalMux I__2570 (
            .O(N__14468),
            .I(N__14452));
    InMux I__2569 (
            .O(N__14467),
            .I(N__14449));
    LocalMux I__2568 (
            .O(N__14464),
            .I(N__14446));
    LocalMux I__2567 (
            .O(N__14461),
            .I(N__14443));
    InMux I__2566 (
            .O(N__14460),
            .I(N__14440));
    LocalMux I__2565 (
            .O(N__14457),
            .I(N__14437));
    InMux I__2564 (
            .O(N__14456),
            .I(N__14434));
    InMux I__2563 (
            .O(N__14455),
            .I(N__14431));
    Span4Mux_h I__2562 (
            .O(N__14452),
            .I(N__14423));
    LocalMux I__2561 (
            .O(N__14449),
            .I(N__14423));
    Span4Mux_h I__2560 (
            .O(N__14446),
            .I(N__14423));
    Span4Mux_v I__2559 (
            .O(N__14443),
            .I(N__14414));
    LocalMux I__2558 (
            .O(N__14440),
            .I(N__14414));
    Span4Mux_v I__2557 (
            .O(N__14437),
            .I(N__14414));
    LocalMux I__2556 (
            .O(N__14434),
            .I(N__14414));
    LocalMux I__2555 (
            .O(N__14431),
            .I(N__14411));
    InMux I__2554 (
            .O(N__14430),
            .I(N__14408));
    Odrv4 I__2553 (
            .O(N__14423),
            .I(RX_ADDR_11));
    Odrv4 I__2552 (
            .O(N__14414),
            .I(RX_ADDR_11));
    Odrv4 I__2551 (
            .O(N__14411),
            .I(RX_ADDR_11));
    LocalMux I__2550 (
            .O(N__14408),
            .I(RX_ADDR_11));
    SRMux I__2549 (
            .O(N__14399),
            .I(N__14396));
    LocalMux I__2548 (
            .O(N__14396),
            .I(N__14390));
    SRMux I__2547 (
            .O(N__14395),
            .I(N__14387));
    SRMux I__2546 (
            .O(N__14394),
            .I(N__14384));
    SRMux I__2545 (
            .O(N__14393),
            .I(N__14381));
    Span4Mux_v I__2544 (
            .O(N__14390),
            .I(N__14376));
    LocalMux I__2543 (
            .O(N__14387),
            .I(N__14376));
    LocalMux I__2542 (
            .O(N__14384),
            .I(N__14371));
    LocalMux I__2541 (
            .O(N__14381),
            .I(N__14371));
    Span4Mux_v I__2540 (
            .O(N__14376),
            .I(N__14366));
    Span4Mux_v I__2539 (
            .O(N__14371),
            .I(N__14366));
    Sp12to4 I__2538 (
            .O(N__14366),
            .I(N__14363));
    Odrv12 I__2537 (
            .O(N__14363),
            .I(\line_buffer.n532 ));
    InMux I__2536 (
            .O(N__14360),
            .I(N__14357));
    LocalMux I__2535 (
            .O(N__14357),
            .I(N__14354));
    Span4Mux_v I__2534 (
            .O(N__14354),
            .I(N__14351));
    Odrv4 I__2533 (
            .O(N__14351),
            .I(\tvp_video_buffer.BUFFER_1_3 ));
    InMux I__2532 (
            .O(N__14348),
            .I(N__14343));
    InMux I__2531 (
            .O(N__14347),
            .I(N__14340));
    InMux I__2530 (
            .O(N__14346),
            .I(N__14336));
    LocalMux I__2529 (
            .O(N__14343),
            .I(N__14331));
    LocalMux I__2528 (
            .O(N__14340),
            .I(N__14328));
    InMux I__2527 (
            .O(N__14339),
            .I(N__14324));
    LocalMux I__2526 (
            .O(N__14336),
            .I(N__14321));
    InMux I__2525 (
            .O(N__14335),
            .I(N__14318));
    InMux I__2524 (
            .O(N__14334),
            .I(N__14315));
    Span4Mux_v I__2523 (
            .O(N__14331),
            .I(N__14312));
    Span4Mux_v I__2522 (
            .O(N__14328),
            .I(N__14309));
    InMux I__2521 (
            .O(N__14327),
            .I(N__14306));
    LocalMux I__2520 (
            .O(N__14324),
            .I(N__14302));
    Span12Mux_s9_v I__2519 (
            .O(N__14321),
            .I(N__14295));
    LocalMux I__2518 (
            .O(N__14318),
            .I(N__14295));
    LocalMux I__2517 (
            .O(N__14315),
            .I(N__14295));
    Span4Mux_v I__2516 (
            .O(N__14312),
            .I(N__14290));
    Span4Mux_v I__2515 (
            .O(N__14309),
            .I(N__14290));
    LocalMux I__2514 (
            .O(N__14306),
            .I(N__14287));
    InMux I__2513 (
            .O(N__14305),
            .I(N__14284));
    Span12Mux_s10_v I__2512 (
            .O(N__14302),
            .I(N__14279));
    Span12Mux_v I__2511 (
            .O(N__14295),
            .I(N__14279));
    Sp12to4 I__2510 (
            .O(N__14290),
            .I(N__14272));
    Span12Mux_h I__2509 (
            .O(N__14287),
            .I(N__14272));
    LocalMux I__2508 (
            .O(N__14284),
            .I(N__14272));
    Odrv12 I__2507 (
            .O(N__14279),
            .I(RX_DATA_1));
    Odrv12 I__2506 (
            .O(N__14272),
            .I(RX_DATA_1));
    InMux I__2505 (
            .O(N__14267),
            .I(N__14264));
    LocalMux I__2504 (
            .O(N__14264),
            .I(N__14261));
    Odrv4 I__2503 (
            .O(N__14261),
            .I(\sync_buffer.BUFFER_1_0 ));
    InMux I__2502 (
            .O(N__14258),
            .I(N__14255));
    LocalMux I__2501 (
            .O(N__14255),
            .I(RX_TX_SYNC_BUFF));
    SRMux I__2500 (
            .O(N__14252),
            .I(N__14249));
    LocalMux I__2499 (
            .O(N__14249),
            .I(N__14243));
    SRMux I__2498 (
            .O(N__14248),
            .I(N__14240));
    CEMux I__2497 (
            .O(N__14247),
            .I(N__14236));
    CEMux I__2496 (
            .O(N__14246),
            .I(N__14233));
    Span4Mux_v I__2495 (
            .O(N__14243),
            .I(N__14228));
    LocalMux I__2494 (
            .O(N__14240),
            .I(N__14228));
    InMux I__2493 (
            .O(N__14239),
            .I(N__14225));
    LocalMux I__2492 (
            .O(N__14236),
            .I(N__14222));
    LocalMux I__2491 (
            .O(N__14233),
            .I(N__14217));
    Span4Mux_h I__2490 (
            .O(N__14228),
            .I(N__14217));
    LocalMux I__2489 (
            .O(N__14225),
            .I(N__14214));
    Odrv12 I__2488 (
            .O(N__14222),
            .I(\transmit_module.video_signal_controller.n2036 ));
    Odrv4 I__2487 (
            .O(N__14217),
            .I(\transmit_module.video_signal_controller.n2036 ));
    Odrv4 I__2486 (
            .O(N__14214),
            .I(\transmit_module.video_signal_controller.n2036 ));
    SRMux I__2485 (
            .O(N__14207),
            .I(N__14204));
    LocalMux I__2484 (
            .O(N__14204),
            .I(N__14200));
    SRMux I__2483 (
            .O(N__14203),
            .I(N__14197));
    Span4Mux_h I__2482 (
            .O(N__14200),
            .I(N__14194));
    LocalMux I__2481 (
            .O(N__14197),
            .I(N__14191));
    Odrv4 I__2480 (
            .O(N__14194),
            .I(\transmit_module.video_signal_controller.n2378 ));
    Odrv12 I__2479 (
            .O(N__14191),
            .I(\transmit_module.video_signal_controller.n2378 ));
    CascadeMux I__2478 (
            .O(N__14186),
            .I(\transmit_module.video_signal_controller.n49_cascade_ ));
    SRMux I__2477 (
            .O(N__14183),
            .I(N__14179));
    SRMux I__2476 (
            .O(N__14182),
            .I(N__14176));
    LocalMux I__2475 (
            .O(N__14179),
            .I(N__14169));
    LocalMux I__2474 (
            .O(N__14176),
            .I(N__14169));
    SRMux I__2473 (
            .O(N__14175),
            .I(N__14166));
    SRMux I__2472 (
            .O(N__14174),
            .I(N__14163));
    Span4Mux_v I__2471 (
            .O(N__14169),
            .I(N__14156));
    LocalMux I__2470 (
            .O(N__14166),
            .I(N__14156));
    LocalMux I__2469 (
            .O(N__14163),
            .I(N__14156));
    Span4Mux_v I__2468 (
            .O(N__14156),
            .I(N__14153));
    Span4Mux_h I__2467 (
            .O(N__14153),
            .I(N__14150));
    Span4Mux_h I__2466 (
            .O(N__14150),
            .I(N__14147));
    Span4Mux_h I__2465 (
            .O(N__14147),
            .I(N__14144));
    Odrv4 I__2464 (
            .O(N__14144),
            .I(\line_buffer.n468 ));
    CascadeMux I__2463 (
            .O(N__14141),
            .I(N__14138));
    CascadeBuf I__2462 (
            .O(N__14138),
            .I(N__14135));
    CascadeMux I__2461 (
            .O(N__14135),
            .I(N__14132));
    CascadeBuf I__2460 (
            .O(N__14132),
            .I(N__14128));
    CascadeMux I__2459 (
            .O(N__14131),
            .I(N__14125));
    CascadeMux I__2458 (
            .O(N__14128),
            .I(N__14122));
    CascadeBuf I__2457 (
            .O(N__14125),
            .I(N__14119));
    CascadeBuf I__2456 (
            .O(N__14122),
            .I(N__14116));
    CascadeMux I__2455 (
            .O(N__14119),
            .I(N__14113));
    CascadeMux I__2454 (
            .O(N__14116),
            .I(N__14110));
    CascadeBuf I__2453 (
            .O(N__14113),
            .I(N__14107));
    CascadeBuf I__2452 (
            .O(N__14110),
            .I(N__14104));
    CascadeMux I__2451 (
            .O(N__14107),
            .I(N__14101));
    CascadeMux I__2450 (
            .O(N__14104),
            .I(N__14098));
    CascadeBuf I__2449 (
            .O(N__14101),
            .I(N__14095));
    CascadeBuf I__2448 (
            .O(N__14098),
            .I(N__14092));
    CascadeMux I__2447 (
            .O(N__14095),
            .I(N__14089));
    CascadeMux I__2446 (
            .O(N__14092),
            .I(N__14086));
    CascadeBuf I__2445 (
            .O(N__14089),
            .I(N__14083));
    CascadeBuf I__2444 (
            .O(N__14086),
            .I(N__14080));
    CascadeMux I__2443 (
            .O(N__14083),
            .I(N__14077));
    CascadeMux I__2442 (
            .O(N__14080),
            .I(N__14074));
    CascadeBuf I__2441 (
            .O(N__14077),
            .I(N__14071));
    CascadeBuf I__2440 (
            .O(N__14074),
            .I(N__14068));
    CascadeMux I__2439 (
            .O(N__14071),
            .I(N__14065));
    CascadeMux I__2438 (
            .O(N__14068),
            .I(N__14062));
    CascadeBuf I__2437 (
            .O(N__14065),
            .I(N__14059));
    CascadeBuf I__2436 (
            .O(N__14062),
            .I(N__14056));
    CascadeMux I__2435 (
            .O(N__14059),
            .I(N__14053));
    CascadeMux I__2434 (
            .O(N__14056),
            .I(N__14050));
    CascadeBuf I__2433 (
            .O(N__14053),
            .I(N__14047));
    CascadeBuf I__2432 (
            .O(N__14050),
            .I(N__14044));
    CascadeMux I__2431 (
            .O(N__14047),
            .I(N__14041));
    CascadeMux I__2430 (
            .O(N__14044),
            .I(N__14038));
    CascadeBuf I__2429 (
            .O(N__14041),
            .I(N__14035));
    CascadeBuf I__2428 (
            .O(N__14038),
            .I(N__14032));
    CascadeMux I__2427 (
            .O(N__14035),
            .I(N__14029));
    CascadeMux I__2426 (
            .O(N__14032),
            .I(N__14026));
    CascadeBuf I__2425 (
            .O(N__14029),
            .I(N__14023));
    CascadeBuf I__2424 (
            .O(N__14026),
            .I(N__14020));
    CascadeMux I__2423 (
            .O(N__14023),
            .I(N__14017));
    CascadeMux I__2422 (
            .O(N__14020),
            .I(N__14014));
    CascadeBuf I__2421 (
            .O(N__14017),
            .I(N__14011));
    CascadeBuf I__2420 (
            .O(N__14014),
            .I(N__14008));
    CascadeMux I__2419 (
            .O(N__14011),
            .I(N__14005));
    CascadeMux I__2418 (
            .O(N__14008),
            .I(N__14002));
    CascadeBuf I__2417 (
            .O(N__14005),
            .I(N__13999));
    CascadeBuf I__2416 (
            .O(N__14002),
            .I(N__13996));
    CascadeMux I__2415 (
            .O(N__13999),
            .I(N__13993));
    CascadeMux I__2414 (
            .O(N__13996),
            .I(N__13990));
    CascadeBuf I__2413 (
            .O(N__13993),
            .I(N__13987));
    CascadeBuf I__2412 (
            .O(N__13990),
            .I(N__13984));
    CascadeMux I__2411 (
            .O(N__13987),
            .I(N__13981));
    CascadeMux I__2410 (
            .O(N__13984),
            .I(N__13978));
    CascadeBuf I__2409 (
            .O(N__13981),
            .I(N__13975));
    CascadeBuf I__2408 (
            .O(N__13978),
            .I(N__13972));
    CascadeMux I__2407 (
            .O(N__13975),
            .I(N__13969));
    CascadeMux I__2406 (
            .O(N__13972),
            .I(N__13966));
    CascadeBuf I__2405 (
            .O(N__13969),
            .I(N__13963));
    InMux I__2404 (
            .O(N__13966),
            .I(N__13960));
    CascadeMux I__2403 (
            .O(N__13963),
            .I(N__13957));
    LocalMux I__2402 (
            .O(N__13960),
            .I(N__13954));
    CascadeBuf I__2401 (
            .O(N__13957),
            .I(N__13951));
    Span4Mux_v I__2400 (
            .O(N__13954),
            .I(N__13948));
    CascadeMux I__2399 (
            .O(N__13951),
            .I(N__13945));
    Span4Mux_v I__2398 (
            .O(N__13948),
            .I(N__13942));
    InMux I__2397 (
            .O(N__13945),
            .I(N__13939));
    Span4Mux_h I__2396 (
            .O(N__13942),
            .I(N__13936));
    LocalMux I__2395 (
            .O(N__13939),
            .I(N__13933));
    Span4Mux_h I__2394 (
            .O(N__13936),
            .I(N__13930));
    Span4Mux_v I__2393 (
            .O(N__13933),
            .I(N__13927));
    Span4Mux_h I__2392 (
            .O(N__13930),
            .I(N__13922));
    Span4Mux_h I__2391 (
            .O(N__13927),
            .I(N__13922));
    Sp12to4 I__2390 (
            .O(N__13922),
            .I(N__13919));
    Odrv12 I__2389 (
            .O(N__13919),
            .I(n25));
    InMux I__2388 (
            .O(N__13916),
            .I(N__13913));
    LocalMux I__2387 (
            .O(N__13913),
            .I(\transmit_module.ADDR_Y_COMPONENT_3 ));
    InMux I__2386 (
            .O(N__13910),
            .I(N__13907));
    LocalMux I__2385 (
            .O(N__13907),
            .I(N__13904));
    Span4Mux_h I__2384 (
            .O(N__13904),
            .I(N__13901));
    Odrv4 I__2383 (
            .O(N__13901),
            .I(\tvp_video_buffer.BUFFER_0_4 ));
    CascadeMux I__2382 (
            .O(N__13898),
            .I(N__13895));
    InMux I__2381 (
            .O(N__13895),
            .I(N__13892));
    LocalMux I__2380 (
            .O(N__13892),
            .I(N__13886));
    InMux I__2379 (
            .O(N__13891),
            .I(N__13883));
    InMux I__2378 (
            .O(N__13890),
            .I(N__13880));
    InMux I__2377 (
            .O(N__13889),
            .I(N__13877));
    Odrv4 I__2376 (
            .O(N__13886),
            .I(\receive_module.rx_counter.Y_4 ));
    LocalMux I__2375 (
            .O(N__13883),
            .I(\receive_module.rx_counter.Y_4 ));
    LocalMux I__2374 (
            .O(N__13880),
            .I(\receive_module.rx_counter.Y_4 ));
    LocalMux I__2373 (
            .O(N__13877),
            .I(\receive_module.rx_counter.Y_4 ));
    InMux I__2372 (
            .O(N__13868),
            .I(N__13864));
    InMux I__2371 (
            .O(N__13867),
            .I(N__13859));
    LocalMux I__2370 (
            .O(N__13864),
            .I(N__13856));
    InMux I__2369 (
            .O(N__13863),
            .I(N__13853));
    InMux I__2368 (
            .O(N__13862),
            .I(N__13850));
    LocalMux I__2367 (
            .O(N__13859),
            .I(\receive_module.rx_counter.Y_7 ));
    Odrv4 I__2366 (
            .O(N__13856),
            .I(\receive_module.rx_counter.Y_7 ));
    LocalMux I__2365 (
            .O(N__13853),
            .I(\receive_module.rx_counter.Y_7 ));
    LocalMux I__2364 (
            .O(N__13850),
            .I(\receive_module.rx_counter.Y_7 ));
    CascadeMux I__2363 (
            .O(N__13841),
            .I(N__13835));
    InMux I__2362 (
            .O(N__13840),
            .I(N__13832));
    InMux I__2361 (
            .O(N__13839),
            .I(N__13829));
    InMux I__2360 (
            .O(N__13838),
            .I(N__13826));
    InMux I__2359 (
            .O(N__13835),
            .I(N__13823));
    LocalMux I__2358 (
            .O(N__13832),
            .I(\receive_module.rx_counter.Y_1 ));
    LocalMux I__2357 (
            .O(N__13829),
            .I(\receive_module.rx_counter.Y_1 ));
    LocalMux I__2356 (
            .O(N__13826),
            .I(\receive_module.rx_counter.Y_1 ));
    LocalMux I__2355 (
            .O(N__13823),
            .I(\receive_module.rx_counter.Y_1 ));
    InMux I__2354 (
            .O(N__13814),
            .I(N__13808));
    InMux I__2353 (
            .O(N__13813),
            .I(N__13805));
    InMux I__2352 (
            .O(N__13812),
            .I(N__13800));
    InMux I__2351 (
            .O(N__13811),
            .I(N__13800));
    LocalMux I__2350 (
            .O(N__13808),
            .I(\receive_module.rx_counter.Y_3 ));
    LocalMux I__2349 (
            .O(N__13805),
            .I(\receive_module.rx_counter.Y_3 ));
    LocalMux I__2348 (
            .O(N__13800),
            .I(\receive_module.rx_counter.Y_3 ));
    CascadeMux I__2347 (
            .O(N__13793),
            .I(N__13790));
    InMux I__2346 (
            .O(N__13790),
            .I(N__13784));
    InMux I__2345 (
            .O(N__13789),
            .I(N__13781));
    InMux I__2344 (
            .O(N__13788),
            .I(N__13776));
    InMux I__2343 (
            .O(N__13787),
            .I(N__13776));
    LocalMux I__2342 (
            .O(N__13784),
            .I(\receive_module.rx_counter.Y_2 ));
    LocalMux I__2341 (
            .O(N__13781),
            .I(\receive_module.rx_counter.Y_2 ));
    LocalMux I__2340 (
            .O(N__13776),
            .I(\receive_module.rx_counter.Y_2 ));
    CascadeMux I__2339 (
            .O(N__13769),
            .I(N__13765));
    InMux I__2338 (
            .O(N__13768),
            .I(N__13758));
    InMux I__2337 (
            .O(N__13765),
            .I(N__13758));
    InMux I__2336 (
            .O(N__13764),
            .I(N__13755));
    InMux I__2335 (
            .O(N__13763),
            .I(N__13752));
    LocalMux I__2334 (
            .O(N__13758),
            .I(N__13747));
    LocalMux I__2333 (
            .O(N__13755),
            .I(N__13747));
    LocalMux I__2332 (
            .O(N__13752),
            .I(\receive_module.rx_counter.Y_8 ));
    Odrv4 I__2331 (
            .O(N__13747),
            .I(\receive_module.rx_counter.Y_8 ));
    InMux I__2330 (
            .O(N__13742),
            .I(N__13739));
    LocalMux I__2329 (
            .O(N__13739),
            .I(\receive_module.rx_counter.n10_adj_610 ));
    InMux I__2328 (
            .O(N__13736),
            .I(N__13728));
    InMux I__2327 (
            .O(N__13735),
            .I(N__13728));
    InMux I__2326 (
            .O(N__13734),
            .I(N__13725));
    InMux I__2325 (
            .O(N__13733),
            .I(N__13722));
    LocalMux I__2324 (
            .O(N__13728),
            .I(N__13719));
    LocalMux I__2323 (
            .O(N__13725),
            .I(\receive_module.rx_counter.Y_0 ));
    LocalMux I__2322 (
            .O(N__13722),
            .I(\receive_module.rx_counter.Y_0 ));
    Odrv4 I__2321 (
            .O(N__13719),
            .I(\receive_module.rx_counter.Y_0 ));
    CascadeMux I__2320 (
            .O(N__13712),
            .I(\receive_module.rx_counter.n14_cascade_ ));
    InMux I__2319 (
            .O(N__13709),
            .I(N__13705));
    InMux I__2318 (
            .O(N__13708),
            .I(N__13702));
    LocalMux I__2317 (
            .O(N__13705),
            .I(\receive_module.rx_counter.n3633 ));
    LocalMux I__2316 (
            .O(N__13702),
            .I(\receive_module.rx_counter.n3633 ));
    CascadeMux I__2315 (
            .O(N__13697),
            .I(\transmit_module.video_signal_controller.n2947_cascade_ ));
    CascadeMux I__2314 (
            .O(N__13694),
            .I(N__13691));
    InMux I__2313 (
            .O(N__13691),
            .I(N__13688));
    LocalMux I__2312 (
            .O(N__13688),
            .I(N__13685));
    Span12Mux_v I__2311 (
            .O(N__13685),
            .I(N__13682));
    Span12Mux_h I__2310 (
            .O(N__13682),
            .I(N__13679));
    Odrv12 I__2309 (
            .O(N__13679),
            .I(\line_buffer.n522 ));
    InMux I__2308 (
            .O(N__13676),
            .I(N__13673));
    LocalMux I__2307 (
            .O(N__13673),
            .I(N__13670));
    Span4Mux_v I__2306 (
            .O(N__13670),
            .I(N__13667));
    Span4Mux_h I__2305 (
            .O(N__13667),
            .I(N__13664));
    Odrv4 I__2304 (
            .O(N__13664),
            .I(\line_buffer.n530 ));
    CascadeMux I__2303 (
            .O(N__13661),
            .I(N__13658));
    InMux I__2302 (
            .O(N__13658),
            .I(N__13652));
    InMux I__2301 (
            .O(N__13657),
            .I(N__13649));
    InMux I__2300 (
            .O(N__13656),
            .I(N__13646));
    InMux I__2299 (
            .O(N__13655),
            .I(N__13643));
    LocalMux I__2298 (
            .O(N__13652),
            .I(\transmit_module.video_signal_controller.VGA_X_3 ));
    LocalMux I__2297 (
            .O(N__13649),
            .I(\transmit_module.video_signal_controller.VGA_X_3 ));
    LocalMux I__2296 (
            .O(N__13646),
            .I(\transmit_module.video_signal_controller.VGA_X_3 ));
    LocalMux I__2295 (
            .O(N__13643),
            .I(\transmit_module.video_signal_controller.VGA_X_3 ));
    InMux I__2294 (
            .O(N__13634),
            .I(N__13628));
    InMux I__2293 (
            .O(N__13633),
            .I(N__13625));
    InMux I__2292 (
            .O(N__13632),
            .I(N__13622));
    InMux I__2291 (
            .O(N__13631),
            .I(N__13619));
    LocalMux I__2290 (
            .O(N__13628),
            .I(\transmit_module.video_signal_controller.VGA_X_5 ));
    LocalMux I__2289 (
            .O(N__13625),
            .I(\transmit_module.video_signal_controller.VGA_X_5 ));
    LocalMux I__2288 (
            .O(N__13622),
            .I(\transmit_module.video_signal_controller.VGA_X_5 ));
    LocalMux I__2287 (
            .O(N__13619),
            .I(\transmit_module.video_signal_controller.VGA_X_5 ));
    InMux I__2286 (
            .O(N__13610),
            .I(N__13607));
    LocalMux I__2285 (
            .O(N__13607),
            .I(\transmit_module.video_signal_controller.n18 ));
    InMux I__2284 (
            .O(N__13604),
            .I(N__13599));
    CascadeMux I__2283 (
            .O(N__13603),
            .I(N__13596));
    InMux I__2282 (
            .O(N__13602),
            .I(N__13592));
    LocalMux I__2281 (
            .O(N__13599),
            .I(N__13589));
    InMux I__2280 (
            .O(N__13596),
            .I(N__13584));
    InMux I__2279 (
            .O(N__13595),
            .I(N__13584));
    LocalMux I__2278 (
            .O(N__13592),
            .I(\transmit_module.video_signal_controller.VGA_X_9 ));
    Odrv4 I__2277 (
            .O(N__13589),
            .I(\transmit_module.video_signal_controller.VGA_X_9 ));
    LocalMux I__2276 (
            .O(N__13584),
            .I(\transmit_module.video_signal_controller.VGA_X_9 ));
    InMux I__2275 (
            .O(N__13577),
            .I(N__13574));
    LocalMux I__2274 (
            .O(N__13574),
            .I(N__13569));
    InMux I__2273 (
            .O(N__13573),
            .I(N__13565));
    InMux I__2272 (
            .O(N__13572),
            .I(N__13562));
    Span4Mux_v I__2271 (
            .O(N__13569),
            .I(N__13559));
    InMux I__2270 (
            .O(N__13568),
            .I(N__13556));
    LocalMux I__2269 (
            .O(N__13565),
            .I(\transmit_module.video_signal_controller.VGA_X_10 ));
    LocalMux I__2268 (
            .O(N__13562),
            .I(\transmit_module.video_signal_controller.VGA_X_10 ));
    Odrv4 I__2267 (
            .O(N__13559),
            .I(\transmit_module.video_signal_controller.VGA_X_10 ));
    LocalMux I__2266 (
            .O(N__13556),
            .I(\transmit_module.video_signal_controller.VGA_X_10 ));
    InMux I__2265 (
            .O(N__13547),
            .I(N__13544));
    LocalMux I__2264 (
            .O(N__13544),
            .I(\transmit_module.video_signal_controller.n4 ));
    InMux I__2263 (
            .O(N__13541),
            .I(N__13535));
    InMux I__2262 (
            .O(N__13540),
            .I(N__13532));
    InMux I__2261 (
            .O(N__13539),
            .I(N__13529));
    InMux I__2260 (
            .O(N__13538),
            .I(N__13526));
    LocalMux I__2259 (
            .O(N__13535),
            .I(\transmit_module.video_signal_controller.VGA_X_7 ));
    LocalMux I__2258 (
            .O(N__13532),
            .I(\transmit_module.video_signal_controller.VGA_X_7 ));
    LocalMux I__2257 (
            .O(N__13529),
            .I(\transmit_module.video_signal_controller.VGA_X_7 ));
    LocalMux I__2256 (
            .O(N__13526),
            .I(\transmit_module.video_signal_controller.VGA_X_7 ));
    CascadeMux I__2255 (
            .O(N__13517),
            .I(\transmit_module.video_signal_controller.n3625_cascade_ ));
    InMux I__2254 (
            .O(N__13514),
            .I(N__13508));
    InMux I__2253 (
            .O(N__13513),
            .I(N__13503));
    InMux I__2252 (
            .O(N__13512),
            .I(N__13503));
    InMux I__2251 (
            .O(N__13511),
            .I(N__13500));
    LocalMux I__2250 (
            .O(N__13508),
            .I(\transmit_module.video_signal_controller.VGA_X_4 ));
    LocalMux I__2249 (
            .O(N__13503),
            .I(\transmit_module.video_signal_controller.VGA_X_4 ));
    LocalMux I__2248 (
            .O(N__13500),
            .I(\transmit_module.video_signal_controller.VGA_X_4 ));
    SRMux I__2247 (
            .O(N__13493),
            .I(N__13490));
    LocalMux I__2246 (
            .O(N__13490),
            .I(N__13487));
    Span4Mux_h I__2245 (
            .O(N__13487),
            .I(N__13481));
    SRMux I__2244 (
            .O(N__13486),
            .I(N__13478));
    SRMux I__2243 (
            .O(N__13485),
            .I(N__13475));
    SRMux I__2242 (
            .O(N__13484),
            .I(N__13472));
    Span4Mux_v I__2241 (
            .O(N__13481),
            .I(N__13467));
    LocalMux I__2240 (
            .O(N__13478),
            .I(N__13467));
    LocalMux I__2239 (
            .O(N__13475),
            .I(N__13464));
    LocalMux I__2238 (
            .O(N__13472),
            .I(N__13461));
    Span4Mux_v I__2237 (
            .O(N__13467),
            .I(N__13456));
    Span4Mux_h I__2236 (
            .O(N__13464),
            .I(N__13456));
    Span4Mux_h I__2235 (
            .O(N__13461),
            .I(N__13453));
    Span4Mux_h I__2234 (
            .O(N__13456),
            .I(N__13448));
    Span4Mux_h I__2233 (
            .O(N__13453),
            .I(N__13448));
    Odrv4 I__2232 (
            .O(N__13448),
            .I(\line_buffer.n597 ));
    InMux I__2231 (
            .O(N__13445),
            .I(N__13442));
    LocalMux I__2230 (
            .O(N__13442),
            .I(N__13439));
    Span4Mux_v I__2229 (
            .O(N__13439),
            .I(N__13436));
    Span4Mux_v I__2228 (
            .O(N__13436),
            .I(N__13433));
    Span4Mux_h I__2227 (
            .O(N__13433),
            .I(N__13430));
    Odrv4 I__2226 (
            .O(N__13430),
            .I(\line_buffer.n594 ));
    InMux I__2225 (
            .O(N__13427),
            .I(N__13424));
    LocalMux I__2224 (
            .O(N__13424),
            .I(N__13421));
    Span4Mux_v I__2223 (
            .O(N__13421),
            .I(N__13418));
    Span4Mux_h I__2222 (
            .O(N__13418),
            .I(N__13415));
    Odrv4 I__2221 (
            .O(N__13415),
            .I(\line_buffer.n586 ));
    InMux I__2220 (
            .O(N__13412),
            .I(N__13409));
    LocalMux I__2219 (
            .O(N__13409),
            .I(\line_buffer.n3591 ));
    InMux I__2218 (
            .O(N__13406),
            .I(\transmit_module.video_signal_controller.n3145 ));
    InMux I__2217 (
            .O(N__13403),
            .I(\transmit_module.video_signal_controller.n3146 ));
    SRMux I__2216 (
            .O(N__13400),
            .I(N__13396));
    SRMux I__2215 (
            .O(N__13399),
            .I(N__13393));
    LocalMux I__2214 (
            .O(N__13396),
            .I(N__13389));
    LocalMux I__2213 (
            .O(N__13393),
            .I(N__13386));
    SRMux I__2212 (
            .O(N__13392),
            .I(N__13383));
    Span4Mux_v I__2211 (
            .O(N__13389),
            .I(N__13380));
    Span4Mux_h I__2210 (
            .O(N__13386),
            .I(N__13375));
    LocalMux I__2209 (
            .O(N__13383),
            .I(N__13375));
    Span4Mux_v I__2208 (
            .O(N__13380),
            .I(N__13371));
    Span4Mux_v I__2207 (
            .O(N__13375),
            .I(N__13368));
    SRMux I__2206 (
            .O(N__13374),
            .I(N__13365));
    Span4Mux_v I__2205 (
            .O(N__13371),
            .I(N__13358));
    Span4Mux_h I__2204 (
            .O(N__13368),
            .I(N__13358));
    LocalMux I__2203 (
            .O(N__13365),
            .I(N__13358));
    Span4Mux_h I__2202 (
            .O(N__13358),
            .I(N__13355));
    Sp12to4 I__2201 (
            .O(N__13355),
            .I(N__13352));
    Odrv12 I__2200 (
            .O(N__13352),
            .I(\line_buffer.n564 ));
    InMux I__2199 (
            .O(N__13349),
            .I(N__13346));
    LocalMux I__2198 (
            .O(N__13346),
            .I(\transmit_module.video_signal_controller.n3624 ));
    InMux I__2197 (
            .O(N__13343),
            .I(N__13337));
    CascadeMux I__2196 (
            .O(N__13342),
            .I(N__13334));
    InMux I__2195 (
            .O(N__13341),
            .I(N__13331));
    InMux I__2194 (
            .O(N__13340),
            .I(N__13328));
    LocalMux I__2193 (
            .O(N__13337),
            .I(N__13325));
    InMux I__2192 (
            .O(N__13334),
            .I(N__13322));
    LocalMux I__2191 (
            .O(N__13331),
            .I(\transmit_module.video_signal_controller.VGA_X_2 ));
    LocalMux I__2190 (
            .O(N__13328),
            .I(\transmit_module.video_signal_controller.VGA_X_2 ));
    Odrv4 I__2189 (
            .O(N__13325),
            .I(\transmit_module.video_signal_controller.VGA_X_2 ));
    LocalMux I__2188 (
            .O(N__13322),
            .I(\transmit_module.video_signal_controller.VGA_X_2 ));
    InMux I__2187 (
            .O(N__13313),
            .I(N__13307));
    InMux I__2186 (
            .O(N__13312),
            .I(N__13304));
    InMux I__2185 (
            .O(N__13311),
            .I(N__13299));
    InMux I__2184 (
            .O(N__13310),
            .I(N__13299));
    LocalMux I__2183 (
            .O(N__13307),
            .I(\transmit_module.video_signal_controller.VGA_X_1 ));
    LocalMux I__2182 (
            .O(N__13304),
            .I(\transmit_module.video_signal_controller.VGA_X_1 ));
    LocalMux I__2181 (
            .O(N__13299),
            .I(\transmit_module.video_signal_controller.VGA_X_1 ));
    InMux I__2180 (
            .O(N__13292),
            .I(N__13287));
    InMux I__2179 (
            .O(N__13291),
            .I(N__13284));
    InMux I__2178 (
            .O(N__13290),
            .I(N__13281));
    LocalMux I__2177 (
            .O(N__13287),
            .I(\transmit_module.video_signal_controller.VGA_X_0 ));
    LocalMux I__2176 (
            .O(N__13284),
            .I(\transmit_module.video_signal_controller.VGA_X_0 ));
    LocalMux I__2175 (
            .O(N__13281),
            .I(\transmit_module.video_signal_controller.VGA_X_0 ));
    CascadeMux I__2174 (
            .O(N__13274),
            .I(N__13271));
    InMux I__2173 (
            .O(N__13271),
            .I(N__13265));
    InMux I__2172 (
            .O(N__13270),
            .I(N__13265));
    LocalMux I__2171 (
            .O(N__13265),
            .I(N__13262));
    Odrv4 I__2170 (
            .O(N__13262),
            .I(\transmit_module.video_signal_controller.n2001 ));
    CascadeMux I__2169 (
            .O(N__13259),
            .I(\transmit_module.video_signal_controller.n2917_cascade_ ));
    InMux I__2168 (
            .O(N__13256),
            .I(N__13250));
    InMux I__2167 (
            .O(N__13255),
            .I(N__13250));
    LocalMux I__2166 (
            .O(N__13250),
            .I(\transmit_module.video_signal_controller.n3313 ));
    InMux I__2165 (
            .O(N__13247),
            .I(\transmit_module.video_signal_controller.n3136 ));
    InMux I__2164 (
            .O(N__13244),
            .I(\transmit_module.video_signal_controller.n3137 ));
    InMux I__2163 (
            .O(N__13241),
            .I(\transmit_module.video_signal_controller.n3138 ));
    InMux I__2162 (
            .O(N__13238),
            .I(\transmit_module.video_signal_controller.n3139 ));
    InMux I__2161 (
            .O(N__13235),
            .I(\transmit_module.video_signal_controller.n3140 ));
    InMux I__2160 (
            .O(N__13232),
            .I(\transmit_module.video_signal_controller.n3141 ));
    InMux I__2159 (
            .O(N__13229),
            .I(\transmit_module.video_signal_controller.n3142 ));
    InMux I__2158 (
            .O(N__13226),
            .I(bfn_13_13_0_));
    InMux I__2157 (
            .O(N__13223),
            .I(\transmit_module.video_signal_controller.n3144 ));
    InMux I__2156 (
            .O(N__13220),
            .I(\receive_module.rx_counter.n3118 ));
    InMux I__2155 (
            .O(N__13217),
            .I(\receive_module.rx_counter.n3119 ));
    InMux I__2154 (
            .O(N__13214),
            .I(\receive_module.rx_counter.n3120 ));
    InMux I__2153 (
            .O(N__13211),
            .I(N__13206));
    InMux I__2152 (
            .O(N__13210),
            .I(N__13201));
    InMux I__2151 (
            .O(N__13209),
            .I(N__13201));
    LocalMux I__2150 (
            .O(N__13206),
            .I(\receive_module.rx_counter.Y_5 ));
    LocalMux I__2149 (
            .O(N__13201),
            .I(\receive_module.rx_counter.Y_5 ));
    InMux I__2148 (
            .O(N__13196),
            .I(\receive_module.rx_counter.n3121 ));
    InMux I__2147 (
            .O(N__13193),
            .I(N__13188));
    InMux I__2146 (
            .O(N__13192),
            .I(N__13185));
    InMux I__2145 (
            .O(N__13191),
            .I(N__13182));
    LocalMux I__2144 (
            .O(N__13188),
            .I(\receive_module.rx_counter.Y_6 ));
    LocalMux I__2143 (
            .O(N__13185),
            .I(\receive_module.rx_counter.Y_6 ));
    LocalMux I__2142 (
            .O(N__13182),
            .I(\receive_module.rx_counter.Y_6 ));
    InMux I__2141 (
            .O(N__13175),
            .I(\receive_module.rx_counter.n3122 ));
    InMux I__2140 (
            .O(N__13172),
            .I(\receive_module.rx_counter.n3123 ));
    InMux I__2139 (
            .O(N__13169),
            .I(bfn_13_10_0_));
    CEMux I__2138 (
            .O(N__13166),
            .I(N__13162));
    CEMux I__2137 (
            .O(N__13165),
            .I(N__13159));
    LocalMux I__2136 (
            .O(N__13162),
            .I(N__13156));
    LocalMux I__2135 (
            .O(N__13159),
            .I(N__13153));
    Odrv4 I__2134 (
            .O(N__13156),
            .I(\receive_module.rx_counter.n2063 ));
    Odrv4 I__2133 (
            .O(N__13153),
            .I(\receive_module.rx_counter.n2063 ));
    InMux I__2132 (
            .O(N__13148),
            .I(N__13145));
    LocalMux I__2131 (
            .O(N__13145),
            .I(\receive_module.n134 ));
    InMux I__2130 (
            .O(N__13142),
            .I(N__13138));
    InMux I__2129 (
            .O(N__13141),
            .I(N__13135));
    LocalMux I__2128 (
            .O(N__13138),
            .I(N__13130));
    LocalMux I__2127 (
            .O(N__13135),
            .I(N__13130));
    Span4Mux_v I__2126 (
            .O(N__13130),
            .I(N__13126));
    InMux I__2125 (
            .O(N__13129),
            .I(N__13123));
    Span4Mux_v I__2124 (
            .O(N__13126),
            .I(N__13111));
    LocalMux I__2123 (
            .O(N__13123),
            .I(N__13111));
    InMux I__2122 (
            .O(N__13122),
            .I(N__13096));
    InMux I__2121 (
            .O(N__13121),
            .I(N__13096));
    InMux I__2120 (
            .O(N__13120),
            .I(N__13096));
    InMux I__2119 (
            .O(N__13119),
            .I(N__13096));
    InMux I__2118 (
            .O(N__13118),
            .I(N__13096));
    InMux I__2117 (
            .O(N__13117),
            .I(N__13096));
    InMux I__2116 (
            .O(N__13116),
            .I(N__13096));
    Span4Mux_v I__2115 (
            .O(N__13111),
            .I(N__13090));
    LocalMux I__2114 (
            .O(N__13096),
            .I(N__13090));
    InMux I__2113 (
            .O(N__13095),
            .I(N__13083));
    Span4Mux_v I__2112 (
            .O(N__13090),
            .I(N__13080));
    InMux I__2111 (
            .O(N__13089),
            .I(N__13077));
    InMux I__2110 (
            .O(N__13088),
            .I(N__13074));
    InMux I__2109 (
            .O(N__13087),
            .I(N__13069));
    InMux I__2108 (
            .O(N__13086),
            .I(N__13069));
    LocalMux I__2107 (
            .O(N__13083),
            .I(N__13064));
    Span4Mux_v I__2106 (
            .O(N__13080),
            .I(N__13059));
    LocalMux I__2105 (
            .O(N__13077),
            .I(N__13059));
    LocalMux I__2104 (
            .O(N__13074),
            .I(N__13054));
    LocalMux I__2103 (
            .O(N__13069),
            .I(N__13054));
    InMux I__2102 (
            .O(N__13068),
            .I(N__13049));
    InMux I__2101 (
            .O(N__13067),
            .I(N__13049));
    Odrv4 I__2100 (
            .O(N__13064),
            .I(TVP_VSYNC_buff));
    Odrv4 I__2099 (
            .O(N__13059),
            .I(TVP_VSYNC_buff));
    Odrv4 I__2098 (
            .O(N__13054),
            .I(TVP_VSYNC_buff));
    LocalMux I__2097 (
            .O(N__13049),
            .I(TVP_VSYNC_buff));
    CascadeMux I__2096 (
            .O(N__13040),
            .I(N__13037));
    CascadeBuf I__2095 (
            .O(N__13037),
            .I(N__13033));
    CascadeMux I__2094 (
            .O(N__13036),
            .I(N__13030));
    CascadeMux I__2093 (
            .O(N__13033),
            .I(N__13027));
    CascadeBuf I__2092 (
            .O(N__13030),
            .I(N__13024));
    CascadeBuf I__2091 (
            .O(N__13027),
            .I(N__13021));
    CascadeMux I__2090 (
            .O(N__13024),
            .I(N__13018));
    CascadeMux I__2089 (
            .O(N__13021),
            .I(N__13015));
    CascadeBuf I__2088 (
            .O(N__13018),
            .I(N__13012));
    CascadeBuf I__2087 (
            .O(N__13015),
            .I(N__13009));
    CascadeMux I__2086 (
            .O(N__13012),
            .I(N__13006));
    CascadeMux I__2085 (
            .O(N__13009),
            .I(N__13003));
    CascadeBuf I__2084 (
            .O(N__13006),
            .I(N__13000));
    CascadeBuf I__2083 (
            .O(N__13003),
            .I(N__12997));
    CascadeMux I__2082 (
            .O(N__13000),
            .I(N__12994));
    CascadeMux I__2081 (
            .O(N__12997),
            .I(N__12991));
    CascadeBuf I__2080 (
            .O(N__12994),
            .I(N__12988));
    CascadeBuf I__2079 (
            .O(N__12991),
            .I(N__12985));
    CascadeMux I__2078 (
            .O(N__12988),
            .I(N__12982));
    CascadeMux I__2077 (
            .O(N__12985),
            .I(N__12979));
    CascadeBuf I__2076 (
            .O(N__12982),
            .I(N__12976));
    CascadeBuf I__2075 (
            .O(N__12979),
            .I(N__12973));
    CascadeMux I__2074 (
            .O(N__12976),
            .I(N__12970));
    CascadeMux I__2073 (
            .O(N__12973),
            .I(N__12967));
    CascadeBuf I__2072 (
            .O(N__12970),
            .I(N__12964));
    CascadeBuf I__2071 (
            .O(N__12967),
            .I(N__12961));
    CascadeMux I__2070 (
            .O(N__12964),
            .I(N__12958));
    CascadeMux I__2069 (
            .O(N__12961),
            .I(N__12955));
    CascadeBuf I__2068 (
            .O(N__12958),
            .I(N__12952));
    CascadeBuf I__2067 (
            .O(N__12955),
            .I(N__12949));
    CascadeMux I__2066 (
            .O(N__12952),
            .I(N__12946));
    CascadeMux I__2065 (
            .O(N__12949),
            .I(N__12943));
    CascadeBuf I__2064 (
            .O(N__12946),
            .I(N__12940));
    CascadeBuf I__2063 (
            .O(N__12943),
            .I(N__12937));
    CascadeMux I__2062 (
            .O(N__12940),
            .I(N__12934));
    CascadeMux I__2061 (
            .O(N__12937),
            .I(N__12931));
    CascadeBuf I__2060 (
            .O(N__12934),
            .I(N__12928));
    CascadeBuf I__2059 (
            .O(N__12931),
            .I(N__12925));
    CascadeMux I__2058 (
            .O(N__12928),
            .I(N__12922));
    CascadeMux I__2057 (
            .O(N__12925),
            .I(N__12919));
    CascadeBuf I__2056 (
            .O(N__12922),
            .I(N__12916));
    CascadeBuf I__2055 (
            .O(N__12919),
            .I(N__12913));
    CascadeMux I__2054 (
            .O(N__12916),
            .I(N__12910));
    CascadeMux I__2053 (
            .O(N__12913),
            .I(N__12907));
    CascadeBuf I__2052 (
            .O(N__12910),
            .I(N__12904));
    CascadeBuf I__2051 (
            .O(N__12907),
            .I(N__12901));
    CascadeMux I__2050 (
            .O(N__12904),
            .I(N__12898));
    CascadeMux I__2049 (
            .O(N__12901),
            .I(N__12895));
    CascadeBuf I__2048 (
            .O(N__12898),
            .I(N__12892));
    CascadeBuf I__2047 (
            .O(N__12895),
            .I(N__12889));
    CascadeMux I__2046 (
            .O(N__12892),
            .I(N__12886));
    CascadeMux I__2045 (
            .O(N__12889),
            .I(N__12883));
    CascadeBuf I__2044 (
            .O(N__12886),
            .I(N__12880));
    CascadeBuf I__2043 (
            .O(N__12883),
            .I(N__12877));
    CascadeMux I__2042 (
            .O(N__12880),
            .I(N__12874));
    CascadeMux I__2041 (
            .O(N__12877),
            .I(N__12871));
    CascadeBuf I__2040 (
            .O(N__12874),
            .I(N__12868));
    CascadeBuf I__2039 (
            .O(N__12871),
            .I(N__12865));
    CascadeMux I__2038 (
            .O(N__12868),
            .I(N__12862));
    CascadeMux I__2037 (
            .O(N__12865),
            .I(N__12859));
    CascadeBuf I__2036 (
            .O(N__12862),
            .I(N__12856));
    InMux I__2035 (
            .O(N__12859),
            .I(N__12853));
    CascadeMux I__2034 (
            .O(N__12856),
            .I(N__12850));
    LocalMux I__2033 (
            .O(N__12853),
            .I(N__12847));
    InMux I__2032 (
            .O(N__12850),
            .I(N__12844));
    Span4Mux_s1_v I__2031 (
            .O(N__12847),
            .I(N__12841));
    LocalMux I__2030 (
            .O(N__12844),
            .I(N__12838));
    Span4Mux_h I__2029 (
            .O(N__12841),
            .I(N__12835));
    Span12Mux_s1_v I__2028 (
            .O(N__12838),
            .I(N__12832));
    Sp12to4 I__2027 (
            .O(N__12835),
            .I(N__12825));
    Span12Mux_h I__2026 (
            .O(N__12832),
            .I(N__12825));
    InMux I__2025 (
            .O(N__12831),
            .I(N__12822));
    InMux I__2024 (
            .O(N__12830),
            .I(N__12819));
    Span12Mux_v I__2023 (
            .O(N__12825),
            .I(N__12816));
    LocalMux I__2022 (
            .O(N__12822),
            .I(RX_ADDR_2));
    LocalMux I__2021 (
            .O(N__12819),
            .I(RX_ADDR_2));
    Odrv12 I__2020 (
            .O(N__12816),
            .I(RX_ADDR_2));
    SRMux I__2019 (
            .O(N__12809),
            .I(N__12805));
    SRMux I__2018 (
            .O(N__12808),
            .I(N__12802));
    LocalMux I__2017 (
            .O(N__12805),
            .I(N__12799));
    LocalMux I__2016 (
            .O(N__12802),
            .I(N__12796));
    Span4Mux_v I__2015 (
            .O(N__12799),
            .I(N__12790));
    Span4Mux_v I__2014 (
            .O(N__12796),
            .I(N__12790));
    SRMux I__2013 (
            .O(N__12795),
            .I(N__12787));
    Span4Mux_v I__2012 (
            .O(N__12790),
            .I(N__12781));
    LocalMux I__2011 (
            .O(N__12787),
            .I(N__12781));
    SRMux I__2010 (
            .O(N__12786),
            .I(N__12778));
    Span4Mux_v I__2009 (
            .O(N__12781),
            .I(N__12773));
    LocalMux I__2008 (
            .O(N__12778),
            .I(N__12773));
    Span4Mux_v I__2007 (
            .O(N__12773),
            .I(N__12768));
    SRMux I__2006 (
            .O(N__12772),
            .I(N__12765));
    SRMux I__2005 (
            .O(N__12771),
            .I(N__12762));
    Span4Mux_v I__2004 (
            .O(N__12768),
            .I(N__12755));
    LocalMux I__2003 (
            .O(N__12765),
            .I(N__12755));
    LocalMux I__2002 (
            .O(N__12762),
            .I(N__12752));
    SRMux I__2001 (
            .O(N__12761),
            .I(N__12749));
    SRMux I__2000 (
            .O(N__12760),
            .I(N__12746));
    Span4Mux_h I__1999 (
            .O(N__12755),
            .I(N__12743));
    Span4Mux_v I__1998 (
            .O(N__12752),
            .I(N__12736));
    LocalMux I__1997 (
            .O(N__12749),
            .I(N__12736));
    LocalMux I__1996 (
            .O(N__12746),
            .I(N__12736));
    Odrv4 I__1995 (
            .O(N__12743),
            .I(\receive_module.n3631 ));
    Odrv4 I__1994 (
            .O(N__12736),
            .I(\receive_module.n3631 ));
    InMux I__1993 (
            .O(N__12731),
            .I(bfn_13_12_0_));
    InMux I__1992 (
            .O(N__12728),
            .I(N__12725));
    LocalMux I__1991 (
            .O(N__12725),
            .I(\receive_module.rx_counter.n4_adj_605 ));
    CascadeMux I__1990 (
            .O(N__12722),
            .I(\receive_module.rx_counter.n3422_cascade_ ));
    InMux I__1989 (
            .O(N__12719),
            .I(N__12716));
    LocalMux I__1988 (
            .O(N__12716),
            .I(\receive_module.rx_counter.n55_adj_606 ));
    InMux I__1987 (
            .O(N__12713),
            .I(N__12710));
    LocalMux I__1986 (
            .O(N__12710),
            .I(\receive_module.rx_counter.n3394 ));
    InMux I__1985 (
            .O(N__12707),
            .I(N__12704));
    LocalMux I__1984 (
            .O(N__12704),
            .I(\receive_module.rx_counter.n5 ));
    InMux I__1983 (
            .O(N__12701),
            .I(N__12698));
    LocalMux I__1982 (
            .O(N__12698),
            .I(\receive_module.rx_counter.n3413 ));
    SRMux I__1981 (
            .O(N__12695),
            .I(N__12692));
    LocalMux I__1980 (
            .O(N__12692),
            .I(N__12687));
    SRMux I__1979 (
            .O(N__12691),
            .I(N__12684));
    SRMux I__1978 (
            .O(N__12690),
            .I(N__12681));
    Span4Mux_s2_v I__1977 (
            .O(N__12687),
            .I(N__12673));
    LocalMux I__1976 (
            .O(N__12684),
            .I(N__12673));
    LocalMux I__1975 (
            .O(N__12681),
            .I(N__12673));
    SRMux I__1974 (
            .O(N__12680),
            .I(N__12670));
    Span4Mux_v I__1973 (
            .O(N__12673),
            .I(N__12667));
    LocalMux I__1972 (
            .O(N__12670),
            .I(N__12664));
    Sp12to4 I__1971 (
            .O(N__12667),
            .I(N__12661));
    Span4Mux_v I__1970 (
            .O(N__12664),
            .I(N__12658));
    Span12Mux_v I__1969 (
            .O(N__12661),
            .I(N__12655));
    Span4Mux_v I__1968 (
            .O(N__12658),
            .I(N__12652));
    Span12Mux_h I__1967 (
            .O(N__12655),
            .I(N__12649));
    Span4Mux_h I__1966 (
            .O(N__12652),
            .I(N__12646));
    Odrv12 I__1965 (
            .O(N__12649),
            .I(\line_buffer.n596 ));
    Odrv4 I__1964 (
            .O(N__12646),
            .I(\line_buffer.n596 ));
    InMux I__1963 (
            .O(N__12641),
            .I(N__12638));
    LocalMux I__1962 (
            .O(N__12638),
            .I(\receive_module.rx_counter.n4_adj_604 ));
    InMux I__1961 (
            .O(N__12635),
            .I(bfn_13_9_0_));
    InMux I__1960 (
            .O(N__12632),
            .I(\receive_module.rx_counter.n3117 ));
    InMux I__1959 (
            .O(N__12629),
            .I(\receive_module.rx_counter.n3159 ));
    InMux I__1958 (
            .O(N__12626),
            .I(\receive_module.rx_counter.n3160 ));
    CEMux I__1957 (
            .O(N__12623),
            .I(N__12619));
    CEMux I__1956 (
            .O(N__12622),
            .I(N__12616));
    LocalMux I__1955 (
            .O(N__12619),
            .I(\receive_module.rx_counter.n3623 ));
    LocalMux I__1954 (
            .O(N__12616),
            .I(\receive_module.rx_counter.n3623 ));
    InMux I__1953 (
            .O(N__12611),
            .I(N__12607));
    InMux I__1952 (
            .O(N__12610),
            .I(N__12604));
    LocalMux I__1951 (
            .O(N__12607),
            .I(\receive_module.rx_counter.FRAME_COUNTER_4 ));
    LocalMux I__1950 (
            .O(N__12604),
            .I(\receive_module.rx_counter.FRAME_COUNTER_4 ));
    InMux I__1949 (
            .O(N__12599),
            .I(N__12595));
    InMux I__1948 (
            .O(N__12598),
            .I(N__12592));
    LocalMux I__1947 (
            .O(N__12595),
            .I(\receive_module.rx_counter.FRAME_COUNTER_2 ));
    LocalMux I__1946 (
            .O(N__12592),
            .I(\receive_module.rx_counter.FRAME_COUNTER_2 ));
    InMux I__1945 (
            .O(N__12587),
            .I(N__12583));
    InMux I__1944 (
            .O(N__12586),
            .I(N__12580));
    LocalMux I__1943 (
            .O(N__12583),
            .I(\receive_module.rx_counter.FRAME_COUNTER_5 ));
    LocalMux I__1942 (
            .O(N__12580),
            .I(\receive_module.rx_counter.FRAME_COUNTER_5 ));
    InMux I__1941 (
            .O(N__12575),
            .I(N__12571));
    InMux I__1940 (
            .O(N__12574),
            .I(N__12568));
    LocalMux I__1939 (
            .O(N__12571),
            .I(\receive_module.rx_counter.FRAME_COUNTER_1 ));
    LocalMux I__1938 (
            .O(N__12568),
            .I(\receive_module.rx_counter.FRAME_COUNTER_1 ));
    InMux I__1937 (
            .O(N__12563),
            .I(N__12559));
    InMux I__1936 (
            .O(N__12562),
            .I(N__12556));
    LocalMux I__1935 (
            .O(N__12559),
            .I(\receive_module.rx_counter.FRAME_COUNTER_0 ));
    LocalMux I__1934 (
            .O(N__12556),
            .I(\receive_module.rx_counter.FRAME_COUNTER_0 ));
    InMux I__1933 (
            .O(N__12551),
            .I(N__12547));
    InMux I__1932 (
            .O(N__12550),
            .I(N__12544));
    LocalMux I__1931 (
            .O(N__12547),
            .I(\receive_module.rx_counter.FRAME_COUNTER_3 ));
    LocalMux I__1930 (
            .O(N__12544),
            .I(\receive_module.rx_counter.FRAME_COUNTER_3 ));
    CascadeMux I__1929 (
            .O(N__12539),
            .I(\receive_module.rx_counter.n3473_cascade_ ));
    InMux I__1928 (
            .O(N__12536),
            .I(N__12533));
    LocalMux I__1927 (
            .O(N__12533),
            .I(\receive_module.rx_counter.n7 ));
    InMux I__1926 (
            .O(N__12530),
            .I(N__12527));
    LocalMux I__1925 (
            .O(N__12527),
            .I(N__12524));
    Odrv4 I__1924 (
            .O(N__12524),
            .I(\receive_module.rx_counter.n11 ));
    InMux I__1923 (
            .O(N__12521),
            .I(N__12517));
    InMux I__1922 (
            .O(N__12520),
            .I(N__12514));
    LocalMux I__1921 (
            .O(N__12517),
            .I(\receive_module.rx_counter.old_VS ));
    LocalMux I__1920 (
            .O(N__12514),
            .I(\receive_module.rx_counter.old_VS ));
    CascadeMux I__1919 (
            .O(N__12509),
            .I(\receive_module.rx_counter.n11_cascade_ ));
    SRMux I__1918 (
            .O(N__12506),
            .I(N__12503));
    LocalMux I__1917 (
            .O(N__12503),
            .I(N__12500));
    Span4Mux_h I__1916 (
            .O(N__12500),
            .I(N__12497));
    Odrv4 I__1915 (
            .O(N__12497),
            .I(\receive_module.rx_counter.n2529 ));
    InMux I__1914 (
            .O(N__12494),
            .I(N__12491));
    LocalMux I__1913 (
            .O(N__12491),
            .I(N__12488));
    Span12Mux_s10_v I__1912 (
            .O(N__12488),
            .I(N__12485));
    Odrv12 I__1911 (
            .O(N__12485),
            .I(\receive_module.n126 ));
    CascadeMux I__1910 (
            .O(N__12482),
            .I(N__12479));
    CascadeBuf I__1909 (
            .O(N__12479),
            .I(N__12476));
    CascadeMux I__1908 (
            .O(N__12476),
            .I(N__12473));
    CascadeBuf I__1907 (
            .O(N__12473),
            .I(N__12469));
    CascadeMux I__1906 (
            .O(N__12472),
            .I(N__12466));
    CascadeMux I__1905 (
            .O(N__12469),
            .I(N__12463));
    CascadeBuf I__1904 (
            .O(N__12466),
            .I(N__12460));
    CascadeBuf I__1903 (
            .O(N__12463),
            .I(N__12457));
    CascadeMux I__1902 (
            .O(N__12460),
            .I(N__12454));
    CascadeMux I__1901 (
            .O(N__12457),
            .I(N__12451));
    CascadeBuf I__1900 (
            .O(N__12454),
            .I(N__12448));
    CascadeBuf I__1899 (
            .O(N__12451),
            .I(N__12445));
    CascadeMux I__1898 (
            .O(N__12448),
            .I(N__12442));
    CascadeMux I__1897 (
            .O(N__12445),
            .I(N__12439));
    CascadeBuf I__1896 (
            .O(N__12442),
            .I(N__12436));
    CascadeBuf I__1895 (
            .O(N__12439),
            .I(N__12433));
    CascadeMux I__1894 (
            .O(N__12436),
            .I(N__12430));
    CascadeMux I__1893 (
            .O(N__12433),
            .I(N__12427));
    CascadeBuf I__1892 (
            .O(N__12430),
            .I(N__12424));
    CascadeBuf I__1891 (
            .O(N__12427),
            .I(N__12421));
    CascadeMux I__1890 (
            .O(N__12424),
            .I(N__12418));
    CascadeMux I__1889 (
            .O(N__12421),
            .I(N__12415));
    CascadeBuf I__1888 (
            .O(N__12418),
            .I(N__12412));
    CascadeBuf I__1887 (
            .O(N__12415),
            .I(N__12409));
    CascadeMux I__1886 (
            .O(N__12412),
            .I(N__12406));
    CascadeMux I__1885 (
            .O(N__12409),
            .I(N__12403));
    CascadeBuf I__1884 (
            .O(N__12406),
            .I(N__12400));
    CascadeBuf I__1883 (
            .O(N__12403),
            .I(N__12397));
    CascadeMux I__1882 (
            .O(N__12400),
            .I(N__12394));
    CascadeMux I__1881 (
            .O(N__12397),
            .I(N__12391));
    CascadeBuf I__1880 (
            .O(N__12394),
            .I(N__12388));
    CascadeBuf I__1879 (
            .O(N__12391),
            .I(N__12385));
    CascadeMux I__1878 (
            .O(N__12388),
            .I(N__12382));
    CascadeMux I__1877 (
            .O(N__12385),
            .I(N__12379));
    CascadeBuf I__1876 (
            .O(N__12382),
            .I(N__12376));
    CascadeBuf I__1875 (
            .O(N__12379),
            .I(N__12373));
    CascadeMux I__1874 (
            .O(N__12376),
            .I(N__12370));
    CascadeMux I__1873 (
            .O(N__12373),
            .I(N__12367));
    CascadeBuf I__1872 (
            .O(N__12370),
            .I(N__12364));
    CascadeBuf I__1871 (
            .O(N__12367),
            .I(N__12361));
    CascadeMux I__1870 (
            .O(N__12364),
            .I(N__12358));
    CascadeMux I__1869 (
            .O(N__12361),
            .I(N__12355));
    CascadeBuf I__1868 (
            .O(N__12358),
            .I(N__12352));
    CascadeBuf I__1867 (
            .O(N__12355),
            .I(N__12349));
    CascadeMux I__1866 (
            .O(N__12352),
            .I(N__12346));
    CascadeMux I__1865 (
            .O(N__12349),
            .I(N__12343));
    CascadeBuf I__1864 (
            .O(N__12346),
            .I(N__12340));
    CascadeBuf I__1863 (
            .O(N__12343),
            .I(N__12337));
    CascadeMux I__1862 (
            .O(N__12340),
            .I(N__12334));
    CascadeMux I__1861 (
            .O(N__12337),
            .I(N__12331));
    CascadeBuf I__1860 (
            .O(N__12334),
            .I(N__12328));
    CascadeBuf I__1859 (
            .O(N__12331),
            .I(N__12325));
    CascadeMux I__1858 (
            .O(N__12328),
            .I(N__12322));
    CascadeMux I__1857 (
            .O(N__12325),
            .I(N__12319));
    CascadeBuf I__1856 (
            .O(N__12322),
            .I(N__12316));
    CascadeBuf I__1855 (
            .O(N__12319),
            .I(N__12313));
    CascadeMux I__1854 (
            .O(N__12316),
            .I(N__12310));
    CascadeMux I__1853 (
            .O(N__12313),
            .I(N__12307));
    CascadeBuf I__1852 (
            .O(N__12310),
            .I(N__12304));
    InMux I__1851 (
            .O(N__12307),
            .I(N__12301));
    CascadeMux I__1850 (
            .O(N__12304),
            .I(N__12298));
    LocalMux I__1849 (
            .O(N__12301),
            .I(N__12295));
    CascadeBuf I__1848 (
            .O(N__12298),
            .I(N__12291));
    Span4Mux_s3_v I__1847 (
            .O(N__12295),
            .I(N__12288));
    InMux I__1846 (
            .O(N__12294),
            .I(N__12285));
    CascadeMux I__1845 (
            .O(N__12291),
            .I(N__12282));
    Span4Mux_h I__1844 (
            .O(N__12288),
            .I(N__12279));
    LocalMux I__1843 (
            .O(N__12285),
            .I(N__12276));
    InMux I__1842 (
            .O(N__12282),
            .I(N__12273));
    Span4Mux_h I__1841 (
            .O(N__12279),
            .I(N__12270));
    Span4Mux_v I__1840 (
            .O(N__12276),
            .I(N__12266));
    LocalMux I__1839 (
            .O(N__12273),
            .I(N__12263));
    Span4Mux_h I__1838 (
            .O(N__12270),
            .I(N__12260));
    InMux I__1837 (
            .O(N__12269),
            .I(N__12257));
    Span4Mux_v I__1836 (
            .O(N__12266),
            .I(N__12254));
    Span12Mux_s9_v I__1835 (
            .O(N__12263),
            .I(N__12251));
    Span4Mux_v I__1834 (
            .O(N__12260),
            .I(N__12248));
    LocalMux I__1833 (
            .O(N__12257),
            .I(RX_ADDR_10));
    Odrv4 I__1832 (
            .O(N__12254),
            .I(RX_ADDR_10));
    Odrv12 I__1831 (
            .O(N__12251),
            .I(RX_ADDR_10));
    Odrv4 I__1830 (
            .O(N__12248),
            .I(RX_ADDR_10));
    InMux I__1829 (
            .O(N__12239),
            .I(N__12236));
    LocalMux I__1828 (
            .O(N__12236),
            .I(N__12233));
    Span12Mux_s10_v I__1827 (
            .O(N__12233),
            .I(N__12230));
    Odrv12 I__1826 (
            .O(N__12230),
            .I(\receive_module.n133 ));
    CascadeMux I__1825 (
            .O(N__12227),
            .I(N__12224));
    CascadeBuf I__1824 (
            .O(N__12224),
            .I(N__12221));
    CascadeMux I__1823 (
            .O(N__12221),
            .I(N__12217));
    CascadeMux I__1822 (
            .O(N__12220),
            .I(N__12214));
    CascadeBuf I__1821 (
            .O(N__12217),
            .I(N__12211));
    CascadeBuf I__1820 (
            .O(N__12214),
            .I(N__12208));
    CascadeMux I__1819 (
            .O(N__12211),
            .I(N__12205));
    CascadeMux I__1818 (
            .O(N__12208),
            .I(N__12202));
    CascadeBuf I__1817 (
            .O(N__12205),
            .I(N__12199));
    CascadeBuf I__1816 (
            .O(N__12202),
            .I(N__12196));
    CascadeMux I__1815 (
            .O(N__12199),
            .I(N__12193));
    CascadeMux I__1814 (
            .O(N__12196),
            .I(N__12190));
    CascadeBuf I__1813 (
            .O(N__12193),
            .I(N__12187));
    CascadeBuf I__1812 (
            .O(N__12190),
            .I(N__12184));
    CascadeMux I__1811 (
            .O(N__12187),
            .I(N__12181));
    CascadeMux I__1810 (
            .O(N__12184),
            .I(N__12178));
    CascadeBuf I__1809 (
            .O(N__12181),
            .I(N__12175));
    CascadeBuf I__1808 (
            .O(N__12178),
            .I(N__12172));
    CascadeMux I__1807 (
            .O(N__12175),
            .I(N__12169));
    CascadeMux I__1806 (
            .O(N__12172),
            .I(N__12166));
    CascadeBuf I__1805 (
            .O(N__12169),
            .I(N__12163));
    CascadeBuf I__1804 (
            .O(N__12166),
            .I(N__12160));
    CascadeMux I__1803 (
            .O(N__12163),
            .I(N__12157));
    CascadeMux I__1802 (
            .O(N__12160),
            .I(N__12154));
    CascadeBuf I__1801 (
            .O(N__12157),
            .I(N__12151));
    CascadeBuf I__1800 (
            .O(N__12154),
            .I(N__12148));
    CascadeMux I__1799 (
            .O(N__12151),
            .I(N__12145));
    CascadeMux I__1798 (
            .O(N__12148),
            .I(N__12142));
    CascadeBuf I__1797 (
            .O(N__12145),
            .I(N__12139));
    CascadeBuf I__1796 (
            .O(N__12142),
            .I(N__12136));
    CascadeMux I__1795 (
            .O(N__12139),
            .I(N__12133));
    CascadeMux I__1794 (
            .O(N__12136),
            .I(N__12130));
    CascadeBuf I__1793 (
            .O(N__12133),
            .I(N__12127));
    CascadeBuf I__1792 (
            .O(N__12130),
            .I(N__12124));
    CascadeMux I__1791 (
            .O(N__12127),
            .I(N__12121));
    CascadeMux I__1790 (
            .O(N__12124),
            .I(N__12118));
    CascadeBuf I__1789 (
            .O(N__12121),
            .I(N__12115));
    CascadeBuf I__1788 (
            .O(N__12118),
            .I(N__12112));
    CascadeMux I__1787 (
            .O(N__12115),
            .I(N__12109));
    CascadeMux I__1786 (
            .O(N__12112),
            .I(N__12106));
    CascadeBuf I__1785 (
            .O(N__12109),
            .I(N__12103));
    CascadeBuf I__1784 (
            .O(N__12106),
            .I(N__12100));
    CascadeMux I__1783 (
            .O(N__12103),
            .I(N__12097));
    CascadeMux I__1782 (
            .O(N__12100),
            .I(N__12094));
    CascadeBuf I__1781 (
            .O(N__12097),
            .I(N__12091));
    CascadeBuf I__1780 (
            .O(N__12094),
            .I(N__12088));
    CascadeMux I__1779 (
            .O(N__12091),
            .I(N__12085));
    CascadeMux I__1778 (
            .O(N__12088),
            .I(N__12082));
    CascadeBuf I__1777 (
            .O(N__12085),
            .I(N__12079));
    CascadeBuf I__1776 (
            .O(N__12082),
            .I(N__12076));
    CascadeMux I__1775 (
            .O(N__12079),
            .I(N__12073));
    CascadeMux I__1774 (
            .O(N__12076),
            .I(N__12070));
    CascadeBuf I__1773 (
            .O(N__12073),
            .I(N__12067));
    CascadeBuf I__1772 (
            .O(N__12070),
            .I(N__12064));
    CascadeMux I__1771 (
            .O(N__12067),
            .I(N__12061));
    CascadeMux I__1770 (
            .O(N__12064),
            .I(N__12058));
    CascadeBuf I__1769 (
            .O(N__12061),
            .I(N__12055));
    CascadeBuf I__1768 (
            .O(N__12058),
            .I(N__12052));
    CascadeMux I__1767 (
            .O(N__12055),
            .I(N__12049));
    CascadeMux I__1766 (
            .O(N__12052),
            .I(N__12046));
    InMux I__1765 (
            .O(N__12049),
            .I(N__12042));
    CascadeBuf I__1764 (
            .O(N__12046),
            .I(N__12039));
    InMux I__1763 (
            .O(N__12045),
            .I(N__12036));
    LocalMux I__1762 (
            .O(N__12042),
            .I(N__12033));
    CascadeMux I__1761 (
            .O(N__12039),
            .I(N__12030));
    LocalMux I__1760 (
            .O(N__12036),
            .I(N__12027));
    Span4Mux_s3_v I__1759 (
            .O(N__12033),
            .I(N__12024));
    InMux I__1758 (
            .O(N__12030),
            .I(N__12021));
    Sp12to4 I__1757 (
            .O(N__12027),
            .I(N__12018));
    Span4Mux_h I__1756 (
            .O(N__12024),
            .I(N__12014));
    LocalMux I__1755 (
            .O(N__12021),
            .I(N__12011));
    Span12Mux_v I__1754 (
            .O(N__12018),
            .I(N__12008));
    InMux I__1753 (
            .O(N__12017),
            .I(N__12005));
    Sp12to4 I__1752 (
            .O(N__12014),
            .I(N__12002));
    Span4Mux_h I__1751 (
            .O(N__12011),
            .I(N__11999));
    Odrv12 I__1750 (
            .O(N__12008),
            .I(RX_ADDR_3));
    LocalMux I__1749 (
            .O(N__12005),
            .I(RX_ADDR_3));
    Odrv12 I__1748 (
            .O(N__12002),
            .I(RX_ADDR_3));
    Odrv4 I__1747 (
            .O(N__11999),
            .I(RX_ADDR_3));
    InMux I__1746 (
            .O(N__11990),
            .I(N__11987));
    LocalMux I__1745 (
            .O(N__11987),
            .I(N__11984));
    Span4Mux_v I__1744 (
            .O(N__11984),
            .I(N__11981));
    Span4Mux_v I__1743 (
            .O(N__11981),
            .I(N__11978));
    Span4Mux_v I__1742 (
            .O(N__11978),
            .I(N__11975));
    Span4Mux_v I__1741 (
            .O(N__11975),
            .I(N__11972));
    Odrv4 I__1740 (
            .O(N__11972),
            .I(\receive_module.n132 ));
    CascadeMux I__1739 (
            .O(N__11969),
            .I(N__11966));
    CascadeBuf I__1738 (
            .O(N__11966),
            .I(N__11963));
    CascadeMux I__1737 (
            .O(N__11963),
            .I(N__11959));
    CascadeMux I__1736 (
            .O(N__11962),
            .I(N__11956));
    CascadeBuf I__1735 (
            .O(N__11959),
            .I(N__11953));
    CascadeBuf I__1734 (
            .O(N__11956),
            .I(N__11950));
    CascadeMux I__1733 (
            .O(N__11953),
            .I(N__11947));
    CascadeMux I__1732 (
            .O(N__11950),
            .I(N__11944));
    CascadeBuf I__1731 (
            .O(N__11947),
            .I(N__11941));
    CascadeBuf I__1730 (
            .O(N__11944),
            .I(N__11938));
    CascadeMux I__1729 (
            .O(N__11941),
            .I(N__11935));
    CascadeMux I__1728 (
            .O(N__11938),
            .I(N__11932));
    CascadeBuf I__1727 (
            .O(N__11935),
            .I(N__11929));
    CascadeBuf I__1726 (
            .O(N__11932),
            .I(N__11926));
    CascadeMux I__1725 (
            .O(N__11929),
            .I(N__11923));
    CascadeMux I__1724 (
            .O(N__11926),
            .I(N__11920));
    CascadeBuf I__1723 (
            .O(N__11923),
            .I(N__11917));
    CascadeBuf I__1722 (
            .O(N__11920),
            .I(N__11914));
    CascadeMux I__1721 (
            .O(N__11917),
            .I(N__11911));
    CascadeMux I__1720 (
            .O(N__11914),
            .I(N__11908));
    CascadeBuf I__1719 (
            .O(N__11911),
            .I(N__11905));
    CascadeBuf I__1718 (
            .O(N__11908),
            .I(N__11902));
    CascadeMux I__1717 (
            .O(N__11905),
            .I(N__11899));
    CascadeMux I__1716 (
            .O(N__11902),
            .I(N__11896));
    CascadeBuf I__1715 (
            .O(N__11899),
            .I(N__11893));
    CascadeBuf I__1714 (
            .O(N__11896),
            .I(N__11890));
    CascadeMux I__1713 (
            .O(N__11893),
            .I(N__11887));
    CascadeMux I__1712 (
            .O(N__11890),
            .I(N__11884));
    CascadeBuf I__1711 (
            .O(N__11887),
            .I(N__11881));
    CascadeBuf I__1710 (
            .O(N__11884),
            .I(N__11878));
    CascadeMux I__1709 (
            .O(N__11881),
            .I(N__11875));
    CascadeMux I__1708 (
            .O(N__11878),
            .I(N__11872));
    CascadeBuf I__1707 (
            .O(N__11875),
            .I(N__11869));
    CascadeBuf I__1706 (
            .O(N__11872),
            .I(N__11866));
    CascadeMux I__1705 (
            .O(N__11869),
            .I(N__11863));
    CascadeMux I__1704 (
            .O(N__11866),
            .I(N__11860));
    CascadeBuf I__1703 (
            .O(N__11863),
            .I(N__11857));
    CascadeBuf I__1702 (
            .O(N__11860),
            .I(N__11854));
    CascadeMux I__1701 (
            .O(N__11857),
            .I(N__11851));
    CascadeMux I__1700 (
            .O(N__11854),
            .I(N__11848));
    CascadeBuf I__1699 (
            .O(N__11851),
            .I(N__11845));
    CascadeBuf I__1698 (
            .O(N__11848),
            .I(N__11842));
    CascadeMux I__1697 (
            .O(N__11845),
            .I(N__11839));
    CascadeMux I__1696 (
            .O(N__11842),
            .I(N__11836));
    CascadeBuf I__1695 (
            .O(N__11839),
            .I(N__11833));
    CascadeBuf I__1694 (
            .O(N__11836),
            .I(N__11830));
    CascadeMux I__1693 (
            .O(N__11833),
            .I(N__11827));
    CascadeMux I__1692 (
            .O(N__11830),
            .I(N__11824));
    CascadeBuf I__1691 (
            .O(N__11827),
            .I(N__11821));
    CascadeBuf I__1690 (
            .O(N__11824),
            .I(N__11818));
    CascadeMux I__1689 (
            .O(N__11821),
            .I(N__11815));
    CascadeMux I__1688 (
            .O(N__11818),
            .I(N__11812));
    CascadeBuf I__1687 (
            .O(N__11815),
            .I(N__11809));
    CascadeBuf I__1686 (
            .O(N__11812),
            .I(N__11806));
    CascadeMux I__1685 (
            .O(N__11809),
            .I(N__11803));
    CascadeMux I__1684 (
            .O(N__11806),
            .I(N__11800));
    CascadeBuf I__1683 (
            .O(N__11803),
            .I(N__11797));
    CascadeBuf I__1682 (
            .O(N__11800),
            .I(N__11794));
    CascadeMux I__1681 (
            .O(N__11797),
            .I(N__11791));
    CascadeMux I__1680 (
            .O(N__11794),
            .I(N__11788));
    InMux I__1679 (
            .O(N__11791),
            .I(N__11784));
    CascadeBuf I__1678 (
            .O(N__11788),
            .I(N__11781));
    InMux I__1677 (
            .O(N__11787),
            .I(N__11778));
    LocalMux I__1676 (
            .O(N__11784),
            .I(N__11775));
    CascadeMux I__1675 (
            .O(N__11781),
            .I(N__11772));
    LocalMux I__1674 (
            .O(N__11778),
            .I(N__11769));
    Span4Mux_h I__1673 (
            .O(N__11775),
            .I(N__11766));
    InMux I__1672 (
            .O(N__11772),
            .I(N__11763));
    Sp12to4 I__1671 (
            .O(N__11769),
            .I(N__11760));
    Sp12to4 I__1670 (
            .O(N__11766),
            .I(N__11756));
    LocalMux I__1669 (
            .O(N__11763),
            .I(N__11753));
    Span12Mux_v I__1668 (
            .O(N__11760),
            .I(N__11750));
    InMux I__1667 (
            .O(N__11759),
            .I(N__11747));
    Span12Mux_s2_v I__1666 (
            .O(N__11756),
            .I(N__11744));
    Span4Mux_s2_v I__1665 (
            .O(N__11753),
            .I(N__11741));
    Odrv12 I__1664 (
            .O(N__11750),
            .I(RX_ADDR_4));
    LocalMux I__1663 (
            .O(N__11747),
            .I(RX_ADDR_4));
    Odrv12 I__1662 (
            .O(N__11744),
            .I(RX_ADDR_4));
    Odrv4 I__1661 (
            .O(N__11741),
            .I(RX_ADDR_4));
    InMux I__1660 (
            .O(N__11732),
            .I(N__11729));
    LocalMux I__1659 (
            .O(N__11729),
            .I(N__11726));
    Odrv4 I__1658 (
            .O(N__11726),
            .I(\tvp_video_buffer.BUFFER_1_2 ));
    InMux I__1657 (
            .O(N__11723),
            .I(N__11718));
    InMux I__1656 (
            .O(N__11722),
            .I(N__11713));
    InMux I__1655 (
            .O(N__11721),
            .I(N__11709));
    LocalMux I__1654 (
            .O(N__11718),
            .I(N__11706));
    InMux I__1653 (
            .O(N__11717),
            .I(N__11703));
    InMux I__1652 (
            .O(N__11716),
            .I(N__11700));
    LocalMux I__1651 (
            .O(N__11713),
            .I(N__11695));
    InMux I__1650 (
            .O(N__11712),
            .I(N__11692));
    LocalMux I__1649 (
            .O(N__11709),
            .I(N__11689));
    Span12Mux_s4_v I__1648 (
            .O(N__11706),
            .I(N__11682));
    LocalMux I__1647 (
            .O(N__11703),
            .I(N__11682));
    LocalMux I__1646 (
            .O(N__11700),
            .I(N__11682));
    InMux I__1645 (
            .O(N__11699),
            .I(N__11679));
    InMux I__1644 (
            .O(N__11698),
            .I(N__11676));
    Span4Mux_v I__1643 (
            .O(N__11695),
            .I(N__11673));
    LocalMux I__1642 (
            .O(N__11692),
            .I(N__11670));
    Span12Mux_h I__1641 (
            .O(N__11689),
            .I(N__11667));
    Span12Mux_v I__1640 (
            .O(N__11682),
            .I(N__11660));
    LocalMux I__1639 (
            .O(N__11679),
            .I(N__11660));
    LocalMux I__1638 (
            .O(N__11676),
            .I(N__11660));
    Span4Mux_v I__1637 (
            .O(N__11673),
            .I(N__11655));
    Span4Mux_h I__1636 (
            .O(N__11670),
            .I(N__11655));
    Span12Mux_v I__1635 (
            .O(N__11667),
            .I(N__11652));
    Span12Mux_v I__1634 (
            .O(N__11660),
            .I(N__11649));
    Span4Mux_h I__1633 (
            .O(N__11655),
            .I(N__11646));
    Odrv12 I__1632 (
            .O(N__11652),
            .I(RX_DATA_0));
    Odrv12 I__1631 (
            .O(N__11649),
            .I(RX_DATA_0));
    Odrv4 I__1630 (
            .O(N__11646),
            .I(RX_DATA_0));
    InMux I__1629 (
            .O(N__11639),
            .I(bfn_13_6_0_));
    InMux I__1628 (
            .O(N__11636),
            .I(\receive_module.rx_counter.n3156 ));
    InMux I__1627 (
            .O(N__11633),
            .I(\receive_module.rx_counter.n3157 ));
    InMux I__1626 (
            .O(N__11630),
            .I(\receive_module.rx_counter.n3158 ));
    InMux I__1625 (
            .O(N__11627),
            .I(N__11624));
    LocalMux I__1624 (
            .O(N__11624),
            .I(N__11621));
    Span4Mux_h I__1623 (
            .O(N__11621),
            .I(N__11618));
    Odrv4 I__1622 (
            .O(N__11618),
            .I(\transmit_module.Y_DELTA_PATTERN_7 ));
    InMux I__1621 (
            .O(N__11615),
            .I(N__11612));
    LocalMux I__1620 (
            .O(N__11612),
            .I(\transmit_module.Y_DELTA_PATTERN_6 ));
    InMux I__1619 (
            .O(N__11609),
            .I(N__11606));
    LocalMux I__1618 (
            .O(N__11606),
            .I(N__11603));
    Span12Mux_v I__1617 (
            .O(N__11603),
            .I(N__11600));
    Odrv12 I__1616 (
            .O(N__11600),
            .I(\receive_module.n131 ));
    CascadeMux I__1615 (
            .O(N__11597),
            .I(N__11593));
    CascadeMux I__1614 (
            .O(N__11596),
            .I(N__11590));
    CascadeBuf I__1613 (
            .O(N__11593),
            .I(N__11587));
    CascadeBuf I__1612 (
            .O(N__11590),
            .I(N__11584));
    CascadeMux I__1611 (
            .O(N__11587),
            .I(N__11581));
    CascadeMux I__1610 (
            .O(N__11584),
            .I(N__11578));
    CascadeBuf I__1609 (
            .O(N__11581),
            .I(N__11575));
    CascadeBuf I__1608 (
            .O(N__11578),
            .I(N__11572));
    CascadeMux I__1607 (
            .O(N__11575),
            .I(N__11569));
    CascadeMux I__1606 (
            .O(N__11572),
            .I(N__11566));
    CascadeBuf I__1605 (
            .O(N__11569),
            .I(N__11563));
    CascadeBuf I__1604 (
            .O(N__11566),
            .I(N__11560));
    CascadeMux I__1603 (
            .O(N__11563),
            .I(N__11557));
    CascadeMux I__1602 (
            .O(N__11560),
            .I(N__11554));
    CascadeBuf I__1601 (
            .O(N__11557),
            .I(N__11551));
    CascadeBuf I__1600 (
            .O(N__11554),
            .I(N__11548));
    CascadeMux I__1599 (
            .O(N__11551),
            .I(N__11545));
    CascadeMux I__1598 (
            .O(N__11548),
            .I(N__11542));
    CascadeBuf I__1597 (
            .O(N__11545),
            .I(N__11539));
    CascadeBuf I__1596 (
            .O(N__11542),
            .I(N__11536));
    CascadeMux I__1595 (
            .O(N__11539),
            .I(N__11533));
    CascadeMux I__1594 (
            .O(N__11536),
            .I(N__11530));
    CascadeBuf I__1593 (
            .O(N__11533),
            .I(N__11527));
    CascadeBuf I__1592 (
            .O(N__11530),
            .I(N__11524));
    CascadeMux I__1591 (
            .O(N__11527),
            .I(N__11521));
    CascadeMux I__1590 (
            .O(N__11524),
            .I(N__11518));
    CascadeBuf I__1589 (
            .O(N__11521),
            .I(N__11515));
    CascadeBuf I__1588 (
            .O(N__11518),
            .I(N__11512));
    CascadeMux I__1587 (
            .O(N__11515),
            .I(N__11509));
    CascadeMux I__1586 (
            .O(N__11512),
            .I(N__11506));
    CascadeBuf I__1585 (
            .O(N__11509),
            .I(N__11503));
    CascadeBuf I__1584 (
            .O(N__11506),
            .I(N__11500));
    CascadeMux I__1583 (
            .O(N__11503),
            .I(N__11497));
    CascadeMux I__1582 (
            .O(N__11500),
            .I(N__11494));
    CascadeBuf I__1581 (
            .O(N__11497),
            .I(N__11491));
    CascadeBuf I__1580 (
            .O(N__11494),
            .I(N__11488));
    CascadeMux I__1579 (
            .O(N__11491),
            .I(N__11485));
    CascadeMux I__1578 (
            .O(N__11488),
            .I(N__11482));
    CascadeBuf I__1577 (
            .O(N__11485),
            .I(N__11479));
    CascadeBuf I__1576 (
            .O(N__11482),
            .I(N__11476));
    CascadeMux I__1575 (
            .O(N__11479),
            .I(N__11473));
    CascadeMux I__1574 (
            .O(N__11476),
            .I(N__11470));
    CascadeBuf I__1573 (
            .O(N__11473),
            .I(N__11467));
    CascadeBuf I__1572 (
            .O(N__11470),
            .I(N__11464));
    CascadeMux I__1571 (
            .O(N__11467),
            .I(N__11461));
    CascadeMux I__1570 (
            .O(N__11464),
            .I(N__11458));
    CascadeBuf I__1569 (
            .O(N__11461),
            .I(N__11455));
    CascadeBuf I__1568 (
            .O(N__11458),
            .I(N__11452));
    CascadeMux I__1567 (
            .O(N__11455),
            .I(N__11449));
    CascadeMux I__1566 (
            .O(N__11452),
            .I(N__11446));
    CascadeBuf I__1565 (
            .O(N__11449),
            .I(N__11443));
    CascadeBuf I__1564 (
            .O(N__11446),
            .I(N__11440));
    CascadeMux I__1563 (
            .O(N__11443),
            .I(N__11437));
    CascadeMux I__1562 (
            .O(N__11440),
            .I(N__11434));
    CascadeBuf I__1561 (
            .O(N__11437),
            .I(N__11431));
    CascadeBuf I__1560 (
            .O(N__11434),
            .I(N__11428));
    CascadeMux I__1559 (
            .O(N__11431),
            .I(N__11425));
    CascadeMux I__1558 (
            .O(N__11428),
            .I(N__11422));
    CascadeBuf I__1557 (
            .O(N__11425),
            .I(N__11419));
    CascadeBuf I__1556 (
            .O(N__11422),
            .I(N__11416));
    CascadeMux I__1555 (
            .O(N__11419),
            .I(N__11413));
    CascadeMux I__1554 (
            .O(N__11416),
            .I(N__11410));
    InMux I__1553 (
            .O(N__11413),
            .I(N__11407));
    InMux I__1552 (
            .O(N__11410),
            .I(N__11404));
    LocalMux I__1551 (
            .O(N__11407),
            .I(N__11400));
    LocalMux I__1550 (
            .O(N__11404),
            .I(N__11397));
    InMux I__1549 (
            .O(N__11403),
            .I(N__11394));
    Span4Mux_s1_v I__1548 (
            .O(N__11400),
            .I(N__11391));
    Span4Mux_s1_v I__1547 (
            .O(N__11397),
            .I(N__11388));
    LocalMux I__1546 (
            .O(N__11394),
            .I(N__11385));
    Span4Mux_h I__1545 (
            .O(N__11391),
            .I(N__11382));
    Span4Mux_v I__1544 (
            .O(N__11388),
            .I(N__11379));
    Span4Mux_h I__1543 (
            .O(N__11385),
            .I(N__11375));
    Sp12to4 I__1542 (
            .O(N__11382),
            .I(N__11372));
    Sp12to4 I__1541 (
            .O(N__11379),
            .I(N__11369));
    InMux I__1540 (
            .O(N__11378),
            .I(N__11366));
    Span4Mux_v I__1539 (
            .O(N__11375),
            .I(N__11363));
    Span12Mux_s5_v I__1538 (
            .O(N__11372),
            .I(N__11358));
    Span12Mux_h I__1537 (
            .O(N__11369),
            .I(N__11358));
    LocalMux I__1536 (
            .O(N__11366),
            .I(RX_ADDR_5));
    Odrv4 I__1535 (
            .O(N__11363),
            .I(RX_ADDR_5));
    Odrv12 I__1534 (
            .O(N__11358),
            .I(RX_ADDR_5));
    InMux I__1533 (
            .O(N__11351),
            .I(N__11348));
    LocalMux I__1532 (
            .O(N__11348),
            .I(N__11345));
    Span4Mux_v I__1531 (
            .O(N__11345),
            .I(N__11342));
    Span4Mux_v I__1530 (
            .O(N__11342),
            .I(N__11339));
    Odrv4 I__1529 (
            .O(N__11339),
            .I(\receive_module.n130 ));
    CascadeMux I__1528 (
            .O(N__11336),
            .I(N__11332));
    CascadeMux I__1527 (
            .O(N__11335),
            .I(N__11329));
    CascadeBuf I__1526 (
            .O(N__11332),
            .I(N__11326));
    CascadeBuf I__1525 (
            .O(N__11329),
            .I(N__11323));
    CascadeMux I__1524 (
            .O(N__11326),
            .I(N__11320));
    CascadeMux I__1523 (
            .O(N__11323),
            .I(N__11317));
    CascadeBuf I__1522 (
            .O(N__11320),
            .I(N__11314));
    CascadeBuf I__1521 (
            .O(N__11317),
            .I(N__11311));
    CascadeMux I__1520 (
            .O(N__11314),
            .I(N__11308));
    CascadeMux I__1519 (
            .O(N__11311),
            .I(N__11305));
    CascadeBuf I__1518 (
            .O(N__11308),
            .I(N__11302));
    CascadeBuf I__1517 (
            .O(N__11305),
            .I(N__11299));
    CascadeMux I__1516 (
            .O(N__11302),
            .I(N__11296));
    CascadeMux I__1515 (
            .O(N__11299),
            .I(N__11293));
    CascadeBuf I__1514 (
            .O(N__11296),
            .I(N__11290));
    CascadeBuf I__1513 (
            .O(N__11293),
            .I(N__11287));
    CascadeMux I__1512 (
            .O(N__11290),
            .I(N__11284));
    CascadeMux I__1511 (
            .O(N__11287),
            .I(N__11281));
    CascadeBuf I__1510 (
            .O(N__11284),
            .I(N__11278));
    CascadeBuf I__1509 (
            .O(N__11281),
            .I(N__11275));
    CascadeMux I__1508 (
            .O(N__11278),
            .I(N__11272));
    CascadeMux I__1507 (
            .O(N__11275),
            .I(N__11269));
    CascadeBuf I__1506 (
            .O(N__11272),
            .I(N__11266));
    CascadeBuf I__1505 (
            .O(N__11269),
            .I(N__11263));
    CascadeMux I__1504 (
            .O(N__11266),
            .I(N__11260));
    CascadeMux I__1503 (
            .O(N__11263),
            .I(N__11257));
    CascadeBuf I__1502 (
            .O(N__11260),
            .I(N__11254));
    CascadeBuf I__1501 (
            .O(N__11257),
            .I(N__11251));
    CascadeMux I__1500 (
            .O(N__11254),
            .I(N__11248));
    CascadeMux I__1499 (
            .O(N__11251),
            .I(N__11245));
    CascadeBuf I__1498 (
            .O(N__11248),
            .I(N__11242));
    CascadeBuf I__1497 (
            .O(N__11245),
            .I(N__11239));
    CascadeMux I__1496 (
            .O(N__11242),
            .I(N__11236));
    CascadeMux I__1495 (
            .O(N__11239),
            .I(N__11233));
    CascadeBuf I__1494 (
            .O(N__11236),
            .I(N__11230));
    CascadeBuf I__1493 (
            .O(N__11233),
            .I(N__11227));
    CascadeMux I__1492 (
            .O(N__11230),
            .I(N__11224));
    CascadeMux I__1491 (
            .O(N__11227),
            .I(N__11221));
    CascadeBuf I__1490 (
            .O(N__11224),
            .I(N__11218));
    CascadeBuf I__1489 (
            .O(N__11221),
            .I(N__11215));
    CascadeMux I__1488 (
            .O(N__11218),
            .I(N__11212));
    CascadeMux I__1487 (
            .O(N__11215),
            .I(N__11209));
    CascadeBuf I__1486 (
            .O(N__11212),
            .I(N__11206));
    CascadeBuf I__1485 (
            .O(N__11209),
            .I(N__11203));
    CascadeMux I__1484 (
            .O(N__11206),
            .I(N__11200));
    CascadeMux I__1483 (
            .O(N__11203),
            .I(N__11197));
    CascadeBuf I__1482 (
            .O(N__11200),
            .I(N__11194));
    CascadeBuf I__1481 (
            .O(N__11197),
            .I(N__11191));
    CascadeMux I__1480 (
            .O(N__11194),
            .I(N__11188));
    CascadeMux I__1479 (
            .O(N__11191),
            .I(N__11185));
    CascadeBuf I__1478 (
            .O(N__11188),
            .I(N__11182));
    CascadeBuf I__1477 (
            .O(N__11185),
            .I(N__11179));
    CascadeMux I__1476 (
            .O(N__11182),
            .I(N__11176));
    CascadeMux I__1475 (
            .O(N__11179),
            .I(N__11173));
    CascadeBuf I__1474 (
            .O(N__11176),
            .I(N__11170));
    CascadeBuf I__1473 (
            .O(N__11173),
            .I(N__11167));
    CascadeMux I__1472 (
            .O(N__11170),
            .I(N__11164));
    CascadeMux I__1471 (
            .O(N__11167),
            .I(N__11161));
    CascadeBuf I__1470 (
            .O(N__11164),
            .I(N__11158));
    CascadeBuf I__1469 (
            .O(N__11161),
            .I(N__11155));
    CascadeMux I__1468 (
            .O(N__11158),
            .I(N__11152));
    CascadeMux I__1467 (
            .O(N__11155),
            .I(N__11149));
    InMux I__1466 (
            .O(N__11152),
            .I(N__11146));
    InMux I__1465 (
            .O(N__11149),
            .I(N__11142));
    LocalMux I__1464 (
            .O(N__11146),
            .I(N__11139));
    InMux I__1463 (
            .O(N__11145),
            .I(N__11136));
    LocalMux I__1462 (
            .O(N__11142),
            .I(N__11133));
    Span4Mux_h I__1461 (
            .O(N__11139),
            .I(N__11130));
    LocalMux I__1460 (
            .O(N__11136),
            .I(N__11126));
    Span4Mux_h I__1459 (
            .O(N__11133),
            .I(N__11123));
    Span4Mux_h I__1458 (
            .O(N__11130),
            .I(N__11120));
    CascadeMux I__1457 (
            .O(N__11129),
            .I(N__11117));
    Span4Mux_h I__1456 (
            .O(N__11126),
            .I(N__11114));
    Sp12to4 I__1455 (
            .O(N__11123),
            .I(N__11111));
    Sp12to4 I__1454 (
            .O(N__11120),
            .I(N__11108));
    InMux I__1453 (
            .O(N__11117),
            .I(N__11105));
    Span4Mux_v I__1452 (
            .O(N__11114),
            .I(N__11102));
    Span12Mux_v I__1451 (
            .O(N__11111),
            .I(N__11097));
    Span12Mux_v I__1450 (
            .O(N__11108),
            .I(N__11097));
    LocalMux I__1449 (
            .O(N__11105),
            .I(RX_ADDR_6));
    Odrv4 I__1448 (
            .O(N__11102),
            .I(RX_ADDR_6));
    Odrv12 I__1447 (
            .O(N__11097),
            .I(RX_ADDR_6));
    InMux I__1446 (
            .O(N__11090),
            .I(N__11087));
    LocalMux I__1445 (
            .O(N__11087),
            .I(N__11084));
    Sp12to4 I__1444 (
            .O(N__11084),
            .I(N__11081));
    Odrv12 I__1443 (
            .O(N__11081),
            .I(\receive_module.n129 ));
    CascadeMux I__1442 (
            .O(N__11078),
            .I(N__11074));
    CascadeMux I__1441 (
            .O(N__11077),
            .I(N__11071));
    CascadeBuf I__1440 (
            .O(N__11074),
            .I(N__11068));
    CascadeBuf I__1439 (
            .O(N__11071),
            .I(N__11065));
    CascadeMux I__1438 (
            .O(N__11068),
            .I(N__11062));
    CascadeMux I__1437 (
            .O(N__11065),
            .I(N__11059));
    CascadeBuf I__1436 (
            .O(N__11062),
            .I(N__11056));
    CascadeBuf I__1435 (
            .O(N__11059),
            .I(N__11053));
    CascadeMux I__1434 (
            .O(N__11056),
            .I(N__11050));
    CascadeMux I__1433 (
            .O(N__11053),
            .I(N__11047));
    CascadeBuf I__1432 (
            .O(N__11050),
            .I(N__11044));
    CascadeBuf I__1431 (
            .O(N__11047),
            .I(N__11041));
    CascadeMux I__1430 (
            .O(N__11044),
            .I(N__11038));
    CascadeMux I__1429 (
            .O(N__11041),
            .I(N__11035));
    CascadeBuf I__1428 (
            .O(N__11038),
            .I(N__11032));
    CascadeBuf I__1427 (
            .O(N__11035),
            .I(N__11029));
    CascadeMux I__1426 (
            .O(N__11032),
            .I(N__11026));
    CascadeMux I__1425 (
            .O(N__11029),
            .I(N__11023));
    CascadeBuf I__1424 (
            .O(N__11026),
            .I(N__11020));
    CascadeBuf I__1423 (
            .O(N__11023),
            .I(N__11017));
    CascadeMux I__1422 (
            .O(N__11020),
            .I(N__11014));
    CascadeMux I__1421 (
            .O(N__11017),
            .I(N__11011));
    CascadeBuf I__1420 (
            .O(N__11014),
            .I(N__11008));
    CascadeBuf I__1419 (
            .O(N__11011),
            .I(N__11005));
    CascadeMux I__1418 (
            .O(N__11008),
            .I(N__11002));
    CascadeMux I__1417 (
            .O(N__11005),
            .I(N__10999));
    CascadeBuf I__1416 (
            .O(N__11002),
            .I(N__10996));
    CascadeBuf I__1415 (
            .O(N__10999),
            .I(N__10993));
    CascadeMux I__1414 (
            .O(N__10996),
            .I(N__10990));
    CascadeMux I__1413 (
            .O(N__10993),
            .I(N__10987));
    CascadeBuf I__1412 (
            .O(N__10990),
            .I(N__10984));
    CascadeBuf I__1411 (
            .O(N__10987),
            .I(N__10981));
    CascadeMux I__1410 (
            .O(N__10984),
            .I(N__10978));
    CascadeMux I__1409 (
            .O(N__10981),
            .I(N__10975));
    CascadeBuf I__1408 (
            .O(N__10978),
            .I(N__10972));
    CascadeBuf I__1407 (
            .O(N__10975),
            .I(N__10969));
    CascadeMux I__1406 (
            .O(N__10972),
            .I(N__10966));
    CascadeMux I__1405 (
            .O(N__10969),
            .I(N__10963));
    CascadeBuf I__1404 (
            .O(N__10966),
            .I(N__10960));
    CascadeBuf I__1403 (
            .O(N__10963),
            .I(N__10957));
    CascadeMux I__1402 (
            .O(N__10960),
            .I(N__10954));
    CascadeMux I__1401 (
            .O(N__10957),
            .I(N__10951));
    CascadeBuf I__1400 (
            .O(N__10954),
            .I(N__10948));
    CascadeBuf I__1399 (
            .O(N__10951),
            .I(N__10945));
    CascadeMux I__1398 (
            .O(N__10948),
            .I(N__10942));
    CascadeMux I__1397 (
            .O(N__10945),
            .I(N__10939));
    CascadeBuf I__1396 (
            .O(N__10942),
            .I(N__10936));
    CascadeBuf I__1395 (
            .O(N__10939),
            .I(N__10933));
    CascadeMux I__1394 (
            .O(N__10936),
            .I(N__10930));
    CascadeMux I__1393 (
            .O(N__10933),
            .I(N__10927));
    CascadeBuf I__1392 (
            .O(N__10930),
            .I(N__10924));
    CascadeBuf I__1391 (
            .O(N__10927),
            .I(N__10921));
    CascadeMux I__1390 (
            .O(N__10924),
            .I(N__10918));
    CascadeMux I__1389 (
            .O(N__10921),
            .I(N__10915));
    CascadeBuf I__1388 (
            .O(N__10918),
            .I(N__10912));
    CascadeBuf I__1387 (
            .O(N__10915),
            .I(N__10909));
    CascadeMux I__1386 (
            .O(N__10912),
            .I(N__10906));
    CascadeMux I__1385 (
            .O(N__10909),
            .I(N__10903));
    CascadeBuf I__1384 (
            .O(N__10906),
            .I(N__10900));
    CascadeBuf I__1383 (
            .O(N__10903),
            .I(N__10897));
    CascadeMux I__1382 (
            .O(N__10900),
            .I(N__10894));
    CascadeMux I__1381 (
            .O(N__10897),
            .I(N__10891));
    InMux I__1380 (
            .O(N__10894),
            .I(N__10888));
    InMux I__1379 (
            .O(N__10891),
            .I(N__10885));
    LocalMux I__1378 (
            .O(N__10888),
            .I(N__10882));
    LocalMux I__1377 (
            .O(N__10885),
            .I(N__10879));
    Span4Mux_s1_v I__1376 (
            .O(N__10882),
            .I(N__10876));
    Span4Mux_s2_v I__1375 (
            .O(N__10879),
            .I(N__10873));
    Sp12to4 I__1374 (
            .O(N__10876),
            .I(N__10869));
    Span4Mux_h I__1373 (
            .O(N__10873),
            .I(N__10866));
    InMux I__1372 (
            .O(N__10872),
            .I(N__10863));
    Span12Mux_h I__1371 (
            .O(N__10869),
            .I(N__10859));
    Span4Mux_v I__1370 (
            .O(N__10866),
            .I(N__10856));
    LocalMux I__1369 (
            .O(N__10863),
            .I(N__10853));
    InMux I__1368 (
            .O(N__10862),
            .I(N__10850));
    Span12Mux_v I__1367 (
            .O(N__10859),
            .I(N__10847));
    Span4Mux_v I__1366 (
            .O(N__10856),
            .I(N__10844));
    Odrv12 I__1365 (
            .O(N__10853),
            .I(RX_ADDR_7));
    LocalMux I__1364 (
            .O(N__10850),
            .I(RX_ADDR_7));
    Odrv12 I__1363 (
            .O(N__10847),
            .I(RX_ADDR_7));
    Odrv4 I__1362 (
            .O(N__10844),
            .I(RX_ADDR_7));
    InMux I__1361 (
            .O(N__10835),
            .I(N__10832));
    LocalMux I__1360 (
            .O(N__10832),
            .I(N__10829));
    Odrv12 I__1359 (
            .O(N__10829),
            .I(\receive_module.n128 ));
    CascadeMux I__1358 (
            .O(N__10826),
            .I(N__10822));
    CascadeMux I__1357 (
            .O(N__10825),
            .I(N__10819));
    CascadeBuf I__1356 (
            .O(N__10822),
            .I(N__10816));
    CascadeBuf I__1355 (
            .O(N__10819),
            .I(N__10813));
    CascadeMux I__1354 (
            .O(N__10816),
            .I(N__10810));
    CascadeMux I__1353 (
            .O(N__10813),
            .I(N__10807));
    CascadeBuf I__1352 (
            .O(N__10810),
            .I(N__10804));
    CascadeBuf I__1351 (
            .O(N__10807),
            .I(N__10801));
    CascadeMux I__1350 (
            .O(N__10804),
            .I(N__10798));
    CascadeMux I__1349 (
            .O(N__10801),
            .I(N__10795));
    CascadeBuf I__1348 (
            .O(N__10798),
            .I(N__10792));
    CascadeBuf I__1347 (
            .O(N__10795),
            .I(N__10789));
    CascadeMux I__1346 (
            .O(N__10792),
            .I(N__10786));
    CascadeMux I__1345 (
            .O(N__10789),
            .I(N__10783));
    CascadeBuf I__1344 (
            .O(N__10786),
            .I(N__10780));
    CascadeBuf I__1343 (
            .O(N__10783),
            .I(N__10777));
    CascadeMux I__1342 (
            .O(N__10780),
            .I(N__10774));
    CascadeMux I__1341 (
            .O(N__10777),
            .I(N__10771));
    CascadeBuf I__1340 (
            .O(N__10774),
            .I(N__10768));
    CascadeBuf I__1339 (
            .O(N__10771),
            .I(N__10765));
    CascadeMux I__1338 (
            .O(N__10768),
            .I(N__10762));
    CascadeMux I__1337 (
            .O(N__10765),
            .I(N__10759));
    CascadeBuf I__1336 (
            .O(N__10762),
            .I(N__10756));
    CascadeBuf I__1335 (
            .O(N__10759),
            .I(N__10753));
    CascadeMux I__1334 (
            .O(N__10756),
            .I(N__10750));
    CascadeMux I__1333 (
            .O(N__10753),
            .I(N__10747));
    CascadeBuf I__1332 (
            .O(N__10750),
            .I(N__10744));
    CascadeBuf I__1331 (
            .O(N__10747),
            .I(N__10741));
    CascadeMux I__1330 (
            .O(N__10744),
            .I(N__10738));
    CascadeMux I__1329 (
            .O(N__10741),
            .I(N__10735));
    CascadeBuf I__1328 (
            .O(N__10738),
            .I(N__10732));
    CascadeBuf I__1327 (
            .O(N__10735),
            .I(N__10729));
    CascadeMux I__1326 (
            .O(N__10732),
            .I(N__10726));
    CascadeMux I__1325 (
            .O(N__10729),
            .I(N__10723));
    CascadeBuf I__1324 (
            .O(N__10726),
            .I(N__10720));
    CascadeBuf I__1323 (
            .O(N__10723),
            .I(N__10717));
    CascadeMux I__1322 (
            .O(N__10720),
            .I(N__10714));
    CascadeMux I__1321 (
            .O(N__10717),
            .I(N__10711));
    CascadeBuf I__1320 (
            .O(N__10714),
            .I(N__10708));
    CascadeBuf I__1319 (
            .O(N__10711),
            .I(N__10705));
    CascadeMux I__1318 (
            .O(N__10708),
            .I(N__10702));
    CascadeMux I__1317 (
            .O(N__10705),
            .I(N__10699));
    CascadeBuf I__1316 (
            .O(N__10702),
            .I(N__10696));
    CascadeBuf I__1315 (
            .O(N__10699),
            .I(N__10693));
    CascadeMux I__1314 (
            .O(N__10696),
            .I(N__10690));
    CascadeMux I__1313 (
            .O(N__10693),
            .I(N__10687));
    CascadeBuf I__1312 (
            .O(N__10690),
            .I(N__10684));
    CascadeBuf I__1311 (
            .O(N__10687),
            .I(N__10681));
    CascadeMux I__1310 (
            .O(N__10684),
            .I(N__10678));
    CascadeMux I__1309 (
            .O(N__10681),
            .I(N__10675));
    CascadeBuf I__1308 (
            .O(N__10678),
            .I(N__10672));
    CascadeBuf I__1307 (
            .O(N__10675),
            .I(N__10669));
    CascadeMux I__1306 (
            .O(N__10672),
            .I(N__10666));
    CascadeMux I__1305 (
            .O(N__10669),
            .I(N__10663));
    CascadeBuf I__1304 (
            .O(N__10666),
            .I(N__10660));
    CascadeBuf I__1303 (
            .O(N__10663),
            .I(N__10657));
    CascadeMux I__1302 (
            .O(N__10660),
            .I(N__10654));
    CascadeMux I__1301 (
            .O(N__10657),
            .I(N__10651));
    CascadeBuf I__1300 (
            .O(N__10654),
            .I(N__10648));
    CascadeBuf I__1299 (
            .O(N__10651),
            .I(N__10645));
    CascadeMux I__1298 (
            .O(N__10648),
            .I(N__10642));
    CascadeMux I__1297 (
            .O(N__10645),
            .I(N__10639));
    InMux I__1296 (
            .O(N__10642),
            .I(N__10636));
    InMux I__1295 (
            .O(N__10639),
            .I(N__10633));
    LocalMux I__1294 (
            .O(N__10636),
            .I(N__10629));
    LocalMux I__1293 (
            .O(N__10633),
            .I(N__10626));
    InMux I__1292 (
            .O(N__10632),
            .I(N__10622));
    Span4Mux_s3_v I__1291 (
            .O(N__10629),
            .I(N__10619));
    Span4Mux_s2_v I__1290 (
            .O(N__10626),
            .I(N__10616));
    CascadeMux I__1289 (
            .O(N__10625),
            .I(N__10613));
    LocalMux I__1288 (
            .O(N__10622),
            .I(N__10610));
    Span4Mux_h I__1287 (
            .O(N__10619),
            .I(N__10607));
    Sp12to4 I__1286 (
            .O(N__10616),
            .I(N__10604));
    InMux I__1285 (
            .O(N__10613),
            .I(N__10601));
    Span4Mux_v I__1284 (
            .O(N__10610),
            .I(N__10598));
    Sp12to4 I__1283 (
            .O(N__10607),
            .I(N__10593));
    Span12Mux_h I__1282 (
            .O(N__10604),
            .I(N__10593));
    LocalMux I__1281 (
            .O(N__10601),
            .I(RX_ADDR_8));
    Odrv4 I__1280 (
            .O(N__10598),
            .I(RX_ADDR_8));
    Odrv12 I__1279 (
            .O(N__10593),
            .I(RX_ADDR_8));
    InMux I__1278 (
            .O(N__10586),
            .I(N__10583));
    LocalMux I__1277 (
            .O(N__10583),
            .I(N__10580));
    Odrv12 I__1276 (
            .O(N__10580),
            .I(\receive_module.n127 ));
    CascadeMux I__1275 (
            .O(N__10577),
            .I(N__10574));
    CascadeBuf I__1274 (
            .O(N__10574),
            .I(N__10570));
    CascadeMux I__1273 (
            .O(N__10573),
            .I(N__10567));
    CascadeMux I__1272 (
            .O(N__10570),
            .I(N__10564));
    CascadeBuf I__1271 (
            .O(N__10567),
            .I(N__10561));
    CascadeBuf I__1270 (
            .O(N__10564),
            .I(N__10558));
    CascadeMux I__1269 (
            .O(N__10561),
            .I(N__10555));
    CascadeMux I__1268 (
            .O(N__10558),
            .I(N__10552));
    CascadeBuf I__1267 (
            .O(N__10555),
            .I(N__10549));
    CascadeBuf I__1266 (
            .O(N__10552),
            .I(N__10546));
    CascadeMux I__1265 (
            .O(N__10549),
            .I(N__10543));
    CascadeMux I__1264 (
            .O(N__10546),
            .I(N__10540));
    CascadeBuf I__1263 (
            .O(N__10543),
            .I(N__10537));
    CascadeBuf I__1262 (
            .O(N__10540),
            .I(N__10534));
    CascadeMux I__1261 (
            .O(N__10537),
            .I(N__10531));
    CascadeMux I__1260 (
            .O(N__10534),
            .I(N__10528));
    CascadeBuf I__1259 (
            .O(N__10531),
            .I(N__10525));
    CascadeBuf I__1258 (
            .O(N__10528),
            .I(N__10522));
    CascadeMux I__1257 (
            .O(N__10525),
            .I(N__10519));
    CascadeMux I__1256 (
            .O(N__10522),
            .I(N__10516));
    CascadeBuf I__1255 (
            .O(N__10519),
            .I(N__10513));
    CascadeBuf I__1254 (
            .O(N__10516),
            .I(N__10510));
    CascadeMux I__1253 (
            .O(N__10513),
            .I(N__10507));
    CascadeMux I__1252 (
            .O(N__10510),
            .I(N__10504));
    CascadeBuf I__1251 (
            .O(N__10507),
            .I(N__10501));
    CascadeBuf I__1250 (
            .O(N__10504),
            .I(N__10498));
    CascadeMux I__1249 (
            .O(N__10501),
            .I(N__10495));
    CascadeMux I__1248 (
            .O(N__10498),
            .I(N__10492));
    CascadeBuf I__1247 (
            .O(N__10495),
            .I(N__10489));
    CascadeBuf I__1246 (
            .O(N__10492),
            .I(N__10486));
    CascadeMux I__1245 (
            .O(N__10489),
            .I(N__10483));
    CascadeMux I__1244 (
            .O(N__10486),
            .I(N__10480));
    CascadeBuf I__1243 (
            .O(N__10483),
            .I(N__10477));
    CascadeBuf I__1242 (
            .O(N__10480),
            .I(N__10474));
    CascadeMux I__1241 (
            .O(N__10477),
            .I(N__10471));
    CascadeMux I__1240 (
            .O(N__10474),
            .I(N__10468));
    CascadeBuf I__1239 (
            .O(N__10471),
            .I(N__10465));
    CascadeBuf I__1238 (
            .O(N__10468),
            .I(N__10462));
    CascadeMux I__1237 (
            .O(N__10465),
            .I(N__10459));
    CascadeMux I__1236 (
            .O(N__10462),
            .I(N__10456));
    CascadeBuf I__1235 (
            .O(N__10459),
            .I(N__10453));
    CascadeBuf I__1234 (
            .O(N__10456),
            .I(N__10450));
    CascadeMux I__1233 (
            .O(N__10453),
            .I(N__10447));
    CascadeMux I__1232 (
            .O(N__10450),
            .I(N__10444));
    CascadeBuf I__1231 (
            .O(N__10447),
            .I(N__10441));
    CascadeBuf I__1230 (
            .O(N__10444),
            .I(N__10438));
    CascadeMux I__1229 (
            .O(N__10441),
            .I(N__10435));
    CascadeMux I__1228 (
            .O(N__10438),
            .I(N__10432));
    CascadeBuf I__1227 (
            .O(N__10435),
            .I(N__10429));
    CascadeBuf I__1226 (
            .O(N__10432),
            .I(N__10426));
    CascadeMux I__1225 (
            .O(N__10429),
            .I(N__10423));
    CascadeMux I__1224 (
            .O(N__10426),
            .I(N__10420));
    CascadeBuf I__1223 (
            .O(N__10423),
            .I(N__10417));
    CascadeBuf I__1222 (
            .O(N__10420),
            .I(N__10414));
    CascadeMux I__1221 (
            .O(N__10417),
            .I(N__10411));
    CascadeMux I__1220 (
            .O(N__10414),
            .I(N__10408));
    CascadeBuf I__1219 (
            .O(N__10411),
            .I(N__10405));
    CascadeBuf I__1218 (
            .O(N__10408),
            .I(N__10402));
    CascadeMux I__1217 (
            .O(N__10405),
            .I(N__10399));
    CascadeMux I__1216 (
            .O(N__10402),
            .I(N__10396));
    CascadeBuf I__1215 (
            .O(N__10399),
            .I(N__10393));
    InMux I__1214 (
            .O(N__10396),
            .I(N__10390));
    CascadeMux I__1213 (
            .O(N__10393),
            .I(N__10387));
    LocalMux I__1212 (
            .O(N__10390),
            .I(N__10384));
    InMux I__1211 (
            .O(N__10387),
            .I(N__10381));
    Span4Mux_s2_v I__1210 (
            .O(N__10384),
            .I(N__10378));
    LocalMux I__1209 (
            .O(N__10381),
            .I(N__10375));
    Span4Mux_h I__1208 (
            .O(N__10378),
            .I(N__10372));
    Span4Mux_s2_v I__1207 (
            .O(N__10375),
            .I(N__10368));
    Span4Mux_h I__1206 (
            .O(N__10372),
            .I(N__10365));
    InMux I__1205 (
            .O(N__10371),
            .I(N__10362));
    Span4Mux_h I__1204 (
            .O(N__10368),
            .I(N__10357));
    Span4Mux_h I__1203 (
            .O(N__10365),
            .I(N__10357));
    LocalMux I__1202 (
            .O(N__10362),
            .I(N__10353));
    Span4Mux_v I__1201 (
            .O(N__10357),
            .I(N__10350));
    InMux I__1200 (
            .O(N__10356),
            .I(N__10347));
    Span4Mux_v I__1199 (
            .O(N__10353),
            .I(N__10344));
    Span4Mux_v I__1198 (
            .O(N__10350),
            .I(N__10341));
    LocalMux I__1197 (
            .O(N__10347),
            .I(RX_ADDR_9));
    Odrv4 I__1196 (
            .O(N__10344),
            .I(RX_ADDR_9));
    Odrv4 I__1195 (
            .O(N__10341),
            .I(RX_ADDR_9));
    InMux I__1194 (
            .O(N__10334),
            .I(N__10331));
    LocalMux I__1193 (
            .O(N__10331),
            .I(N__10328));
    Odrv12 I__1192 (
            .O(N__10328),
            .I(\receive_module.n136 ));
    CascadeMux I__1191 (
            .O(N__10325),
            .I(N__10321));
    CascadeMux I__1190 (
            .O(N__10324),
            .I(N__10318));
    CascadeBuf I__1189 (
            .O(N__10321),
            .I(N__10315));
    CascadeBuf I__1188 (
            .O(N__10318),
            .I(N__10312));
    CascadeMux I__1187 (
            .O(N__10315),
            .I(N__10309));
    CascadeMux I__1186 (
            .O(N__10312),
            .I(N__10306));
    CascadeBuf I__1185 (
            .O(N__10309),
            .I(N__10303));
    CascadeBuf I__1184 (
            .O(N__10306),
            .I(N__10300));
    CascadeMux I__1183 (
            .O(N__10303),
            .I(N__10297));
    CascadeMux I__1182 (
            .O(N__10300),
            .I(N__10294));
    CascadeBuf I__1181 (
            .O(N__10297),
            .I(N__10291));
    CascadeBuf I__1180 (
            .O(N__10294),
            .I(N__10288));
    CascadeMux I__1179 (
            .O(N__10291),
            .I(N__10285));
    CascadeMux I__1178 (
            .O(N__10288),
            .I(N__10282));
    CascadeBuf I__1177 (
            .O(N__10285),
            .I(N__10279));
    CascadeBuf I__1176 (
            .O(N__10282),
            .I(N__10276));
    CascadeMux I__1175 (
            .O(N__10279),
            .I(N__10273));
    CascadeMux I__1174 (
            .O(N__10276),
            .I(N__10270));
    CascadeBuf I__1173 (
            .O(N__10273),
            .I(N__10267));
    CascadeBuf I__1172 (
            .O(N__10270),
            .I(N__10264));
    CascadeMux I__1171 (
            .O(N__10267),
            .I(N__10261));
    CascadeMux I__1170 (
            .O(N__10264),
            .I(N__10258));
    CascadeBuf I__1169 (
            .O(N__10261),
            .I(N__10255));
    CascadeBuf I__1168 (
            .O(N__10258),
            .I(N__10252));
    CascadeMux I__1167 (
            .O(N__10255),
            .I(N__10249));
    CascadeMux I__1166 (
            .O(N__10252),
            .I(N__10246));
    CascadeBuf I__1165 (
            .O(N__10249),
            .I(N__10243));
    CascadeBuf I__1164 (
            .O(N__10246),
            .I(N__10240));
    CascadeMux I__1163 (
            .O(N__10243),
            .I(N__10237));
    CascadeMux I__1162 (
            .O(N__10240),
            .I(N__10234));
    CascadeBuf I__1161 (
            .O(N__10237),
            .I(N__10231));
    CascadeBuf I__1160 (
            .O(N__10234),
            .I(N__10228));
    CascadeMux I__1159 (
            .O(N__10231),
            .I(N__10225));
    CascadeMux I__1158 (
            .O(N__10228),
            .I(N__10222));
    CascadeBuf I__1157 (
            .O(N__10225),
            .I(N__10219));
    CascadeBuf I__1156 (
            .O(N__10222),
            .I(N__10216));
    CascadeMux I__1155 (
            .O(N__10219),
            .I(N__10213));
    CascadeMux I__1154 (
            .O(N__10216),
            .I(N__10210));
    CascadeBuf I__1153 (
            .O(N__10213),
            .I(N__10207));
    CascadeBuf I__1152 (
            .O(N__10210),
            .I(N__10204));
    CascadeMux I__1151 (
            .O(N__10207),
            .I(N__10201));
    CascadeMux I__1150 (
            .O(N__10204),
            .I(N__10198));
    CascadeBuf I__1149 (
            .O(N__10201),
            .I(N__10195));
    CascadeBuf I__1148 (
            .O(N__10198),
            .I(N__10192));
    CascadeMux I__1147 (
            .O(N__10195),
            .I(N__10189));
    CascadeMux I__1146 (
            .O(N__10192),
            .I(N__10186));
    CascadeBuf I__1145 (
            .O(N__10189),
            .I(N__10183));
    CascadeBuf I__1144 (
            .O(N__10186),
            .I(N__10180));
    CascadeMux I__1143 (
            .O(N__10183),
            .I(N__10177));
    CascadeMux I__1142 (
            .O(N__10180),
            .I(N__10174));
    CascadeBuf I__1141 (
            .O(N__10177),
            .I(N__10171));
    CascadeBuf I__1140 (
            .O(N__10174),
            .I(N__10168));
    CascadeMux I__1139 (
            .O(N__10171),
            .I(N__10165));
    CascadeMux I__1138 (
            .O(N__10168),
            .I(N__10162));
    CascadeBuf I__1137 (
            .O(N__10165),
            .I(N__10159));
    CascadeBuf I__1136 (
            .O(N__10162),
            .I(N__10156));
    CascadeMux I__1135 (
            .O(N__10159),
            .I(N__10153));
    CascadeMux I__1134 (
            .O(N__10156),
            .I(N__10150));
    CascadeBuf I__1133 (
            .O(N__10153),
            .I(N__10147));
    CascadeBuf I__1132 (
            .O(N__10150),
            .I(N__10144));
    CascadeMux I__1131 (
            .O(N__10147),
            .I(N__10141));
    CascadeMux I__1130 (
            .O(N__10144),
            .I(N__10138));
    InMux I__1129 (
            .O(N__10141),
            .I(N__10135));
    InMux I__1128 (
            .O(N__10138),
            .I(N__10132));
    LocalMux I__1127 (
            .O(N__10135),
            .I(N__10129));
    LocalMux I__1126 (
            .O(N__10132),
            .I(N__10125));
    Span4Mux_s1_v I__1125 (
            .O(N__10129),
            .I(N__10122));
    InMux I__1124 (
            .O(N__10128),
            .I(N__10119));
    Span4Mux_s2_v I__1123 (
            .O(N__10125),
            .I(N__10116));
    Span4Mux_h I__1122 (
            .O(N__10122),
            .I(N__10113));
    LocalMux I__1121 (
            .O(N__10119),
            .I(N__10110));
    Span4Mux_h I__1120 (
            .O(N__10116),
            .I(N__10107));
    Sp12to4 I__1119 (
            .O(N__10113),
            .I(N__10103));
    Span4Mux_v I__1118 (
            .O(N__10110),
            .I(N__10100));
    Span4Mux_v I__1117 (
            .O(N__10107),
            .I(N__10097));
    InMux I__1116 (
            .O(N__10106),
            .I(N__10094));
    Span12Mux_v I__1115 (
            .O(N__10103),
            .I(N__10091));
    Span4Mux_v I__1114 (
            .O(N__10100),
            .I(N__10086));
    Span4Mux_v I__1113 (
            .O(N__10097),
            .I(N__10086));
    LocalMux I__1112 (
            .O(N__10094),
            .I(RX_ADDR_0));
    Odrv12 I__1111 (
            .O(N__10091),
            .I(RX_ADDR_0));
    Odrv4 I__1110 (
            .O(N__10086),
            .I(RX_ADDR_0));
    CascadeMux I__1109 (
            .O(N__10079),
            .I(N__10076));
    InMux I__1108 (
            .O(N__10076),
            .I(N__10073));
    LocalMux I__1107 (
            .O(N__10073),
            .I(N__10070));
    Odrv12 I__1106 (
            .O(N__10070),
            .I(\receive_module.n135 ));
    CascadeMux I__1105 (
            .O(N__10067),
            .I(N__10063));
    CascadeMux I__1104 (
            .O(N__10066),
            .I(N__10060));
    CascadeBuf I__1103 (
            .O(N__10063),
            .I(N__10057));
    CascadeBuf I__1102 (
            .O(N__10060),
            .I(N__10054));
    CascadeMux I__1101 (
            .O(N__10057),
            .I(N__10051));
    CascadeMux I__1100 (
            .O(N__10054),
            .I(N__10048));
    CascadeBuf I__1099 (
            .O(N__10051),
            .I(N__10045));
    CascadeBuf I__1098 (
            .O(N__10048),
            .I(N__10042));
    CascadeMux I__1097 (
            .O(N__10045),
            .I(N__10039));
    CascadeMux I__1096 (
            .O(N__10042),
            .I(N__10036));
    CascadeBuf I__1095 (
            .O(N__10039),
            .I(N__10033));
    CascadeBuf I__1094 (
            .O(N__10036),
            .I(N__10030));
    CascadeMux I__1093 (
            .O(N__10033),
            .I(N__10027));
    CascadeMux I__1092 (
            .O(N__10030),
            .I(N__10024));
    CascadeBuf I__1091 (
            .O(N__10027),
            .I(N__10021));
    CascadeBuf I__1090 (
            .O(N__10024),
            .I(N__10018));
    CascadeMux I__1089 (
            .O(N__10021),
            .I(N__10015));
    CascadeMux I__1088 (
            .O(N__10018),
            .I(N__10012));
    CascadeBuf I__1087 (
            .O(N__10015),
            .I(N__10009));
    CascadeBuf I__1086 (
            .O(N__10012),
            .I(N__10006));
    CascadeMux I__1085 (
            .O(N__10009),
            .I(N__10003));
    CascadeMux I__1084 (
            .O(N__10006),
            .I(N__10000));
    CascadeBuf I__1083 (
            .O(N__10003),
            .I(N__9997));
    CascadeBuf I__1082 (
            .O(N__10000),
            .I(N__9994));
    CascadeMux I__1081 (
            .O(N__9997),
            .I(N__9991));
    CascadeMux I__1080 (
            .O(N__9994),
            .I(N__9988));
    CascadeBuf I__1079 (
            .O(N__9991),
            .I(N__9985));
    CascadeBuf I__1078 (
            .O(N__9988),
            .I(N__9982));
    CascadeMux I__1077 (
            .O(N__9985),
            .I(N__9979));
    CascadeMux I__1076 (
            .O(N__9982),
            .I(N__9976));
    CascadeBuf I__1075 (
            .O(N__9979),
            .I(N__9973));
    CascadeBuf I__1074 (
            .O(N__9976),
            .I(N__9970));
    CascadeMux I__1073 (
            .O(N__9973),
            .I(N__9967));
    CascadeMux I__1072 (
            .O(N__9970),
            .I(N__9964));
    CascadeBuf I__1071 (
            .O(N__9967),
            .I(N__9961));
    CascadeBuf I__1070 (
            .O(N__9964),
            .I(N__9958));
    CascadeMux I__1069 (
            .O(N__9961),
            .I(N__9955));
    CascadeMux I__1068 (
            .O(N__9958),
            .I(N__9952));
    CascadeBuf I__1067 (
            .O(N__9955),
            .I(N__9949));
    CascadeBuf I__1066 (
            .O(N__9952),
            .I(N__9946));
    CascadeMux I__1065 (
            .O(N__9949),
            .I(N__9943));
    CascadeMux I__1064 (
            .O(N__9946),
            .I(N__9940));
    CascadeBuf I__1063 (
            .O(N__9943),
            .I(N__9937));
    CascadeBuf I__1062 (
            .O(N__9940),
            .I(N__9934));
    CascadeMux I__1061 (
            .O(N__9937),
            .I(N__9931));
    CascadeMux I__1060 (
            .O(N__9934),
            .I(N__9928));
    CascadeBuf I__1059 (
            .O(N__9931),
            .I(N__9925));
    CascadeBuf I__1058 (
            .O(N__9928),
            .I(N__9922));
    CascadeMux I__1057 (
            .O(N__9925),
            .I(N__9919));
    CascadeMux I__1056 (
            .O(N__9922),
            .I(N__9916));
    CascadeBuf I__1055 (
            .O(N__9919),
            .I(N__9913));
    CascadeBuf I__1054 (
            .O(N__9916),
            .I(N__9910));
    CascadeMux I__1053 (
            .O(N__9913),
            .I(N__9907));
    CascadeMux I__1052 (
            .O(N__9910),
            .I(N__9904));
    CascadeBuf I__1051 (
            .O(N__9907),
            .I(N__9901));
    CascadeBuf I__1050 (
            .O(N__9904),
            .I(N__9898));
    CascadeMux I__1049 (
            .O(N__9901),
            .I(N__9895));
    CascadeMux I__1048 (
            .O(N__9898),
            .I(N__9892));
    CascadeBuf I__1047 (
            .O(N__9895),
            .I(N__9889));
    CascadeBuf I__1046 (
            .O(N__9892),
            .I(N__9886));
    CascadeMux I__1045 (
            .O(N__9889),
            .I(N__9883));
    CascadeMux I__1044 (
            .O(N__9886),
            .I(N__9880));
    InMux I__1043 (
            .O(N__9883),
            .I(N__9877));
    InMux I__1042 (
            .O(N__9880),
            .I(N__9874));
    LocalMux I__1041 (
            .O(N__9877),
            .I(N__9871));
    LocalMux I__1040 (
            .O(N__9874),
            .I(N__9867));
    Span4Mux_s2_v I__1039 (
            .O(N__9871),
            .I(N__9864));
    InMux I__1038 (
            .O(N__9870),
            .I(N__9861));
    Span12Mux_s1_v I__1037 (
            .O(N__9867),
            .I(N__9858));
    Span4Mux_h I__1036 (
            .O(N__9864),
            .I(N__9855));
    LocalMux I__1035 (
            .O(N__9861),
            .I(N__9852));
    Span12Mux_v I__1034 (
            .O(N__9858),
            .I(N__9848));
    Span4Mux_v I__1033 (
            .O(N__9855),
            .I(N__9845));
    Span12Mux_v I__1032 (
            .O(N__9852),
            .I(N__9842));
    InMux I__1031 (
            .O(N__9851),
            .I(N__9839));
    Span12Mux_h I__1030 (
            .O(N__9848),
            .I(N__9836));
    Span4Mux_v I__1029 (
            .O(N__9845),
            .I(N__9833));
    Odrv12 I__1028 (
            .O(N__9842),
            .I(RX_ADDR_1));
    LocalMux I__1027 (
            .O(N__9839),
            .I(RX_ADDR_1));
    Odrv12 I__1026 (
            .O(N__9836),
            .I(RX_ADDR_1));
    Odrv4 I__1025 (
            .O(N__9833),
            .I(RX_ADDR_1));
    InMux I__1024 (
            .O(N__9824),
            .I(N__9821));
    LocalMux I__1023 (
            .O(N__9821),
            .I(N__9818));
    Span12Mux_v I__1022 (
            .O(N__9818),
            .I(N__9815));
    Odrv12 I__1021 (
            .O(N__9815),
            .I(\line_buffer.n593 ));
    InMux I__1020 (
            .O(N__9812),
            .I(N__9809));
    LocalMux I__1019 (
            .O(N__9809),
            .I(N__9806));
    Span12Mux_v I__1018 (
            .O(N__9806),
            .I(N__9803));
    Odrv12 I__1017 (
            .O(N__9803),
            .I(\line_buffer.n585 ));
    InMux I__1016 (
            .O(N__9800),
            .I(\transmit_module.video_signal_controller.n3133 ));
    InMux I__1015 (
            .O(N__9797),
            .I(\transmit_module.video_signal_controller.n3134 ));
    InMux I__1014 (
            .O(N__9794),
            .I(\transmit_module.video_signal_controller.n3135 ));
    InMux I__1013 (
            .O(N__9791),
            .I(N__9788));
    LocalMux I__1012 (
            .O(N__9788),
            .I(\transmit_module.Y_DELTA_PATTERN_2 ));
    InMux I__1011 (
            .O(N__9785),
            .I(N__9782));
    LocalMux I__1010 (
            .O(N__9782),
            .I(\transmit_module.Y_DELTA_PATTERN_3 ));
    InMux I__1009 (
            .O(N__9779),
            .I(N__9776));
    LocalMux I__1008 (
            .O(N__9776),
            .I(\transmit_module.Y_DELTA_PATTERN_5 ));
    InMux I__1007 (
            .O(N__9773),
            .I(N__9770));
    LocalMux I__1006 (
            .O(N__9770),
            .I(\transmit_module.Y_DELTA_PATTERN_4 ));
    InMux I__1005 (
            .O(N__9767),
            .I(bfn_12_15_0_));
    InMux I__1004 (
            .O(N__9764),
            .I(\transmit_module.video_signal_controller.n3125 ));
    InMux I__1003 (
            .O(N__9761),
            .I(\transmit_module.video_signal_controller.n3126 ));
    InMux I__1002 (
            .O(N__9758),
            .I(\transmit_module.video_signal_controller.n3127 ));
    InMux I__1001 (
            .O(N__9755),
            .I(\transmit_module.video_signal_controller.n3128 ));
    InMux I__1000 (
            .O(N__9752),
            .I(\transmit_module.video_signal_controller.n3129 ));
    InMux I__999 (
            .O(N__9749),
            .I(\transmit_module.video_signal_controller.n3130 ));
    InMux I__998 (
            .O(N__9746),
            .I(\transmit_module.video_signal_controller.n3131 ));
    InMux I__997 (
            .O(N__9743),
            .I(bfn_12_16_0_));
    InMux I__996 (
            .O(N__9740),
            .I(\receive_module.n3102 ));
    InMux I__995 (
            .O(N__9737),
            .I(\receive_module.n3103 ));
    CEMux I__994 (
            .O(N__9734),
            .I(N__9731));
    LocalMux I__993 (
            .O(N__9731),
            .I(N__9728));
    Span4Mux_h I__992 (
            .O(N__9728),
            .I(N__9725));
    Odrv4 I__991 (
            .O(N__9725),
            .I(\receive_module.n3632 ));
    InMux I__990 (
            .O(N__9722),
            .I(N__9719));
    LocalMux I__989 (
            .O(N__9719),
            .I(\transmit_module.Y_DELTA_PATTERN_53 ));
    InMux I__988 (
            .O(N__9716),
            .I(N__9713));
    LocalMux I__987 (
            .O(N__9713),
            .I(\transmit_module.Y_DELTA_PATTERN_52 ));
    InMux I__986 (
            .O(N__9710),
            .I(N__9707));
    LocalMux I__985 (
            .O(N__9707),
            .I(\transmit_module.Y_DELTA_PATTERN_56 ));
    InMux I__984 (
            .O(N__9704),
            .I(N__9701));
    LocalMux I__983 (
            .O(N__9701),
            .I(\transmit_module.Y_DELTA_PATTERN_55 ));
    InMux I__982 (
            .O(N__9698),
            .I(N__9695));
    LocalMux I__981 (
            .O(N__9695),
            .I(\transmit_module.Y_DELTA_PATTERN_54 ));
    CascadeMux I__980 (
            .O(N__9692),
            .I(\transmit_module.video_signal_controller.n3629_cascade_ ));
    InMux I__979 (
            .O(N__9689),
            .I(N__9686));
    LocalMux I__978 (
            .O(N__9686),
            .I(\transmit_module.video_signal_controller.n2901 ));
    InMux I__977 (
            .O(N__9683),
            .I(\receive_module.n3093 ));
    InMux I__976 (
            .O(N__9680),
            .I(\receive_module.n3094 ));
    InMux I__975 (
            .O(N__9677),
            .I(\receive_module.n3095 ));
    InMux I__974 (
            .O(N__9674),
            .I(\receive_module.n3096 ));
    InMux I__973 (
            .O(N__9671),
            .I(\receive_module.n3097 ));
    InMux I__972 (
            .O(N__9668),
            .I(bfn_12_12_0_));
    InMux I__971 (
            .O(N__9665),
            .I(\receive_module.n3099 ));
    InMux I__970 (
            .O(N__9662),
            .I(\receive_module.n3100 ));
    InMux I__969 (
            .O(N__9659),
            .I(\receive_module.n3101 ));
    CascadeMux I__968 (
            .O(N__9656),
            .I(\receive_module.rx_counter.n4_cascade_ ));
    InMux I__967 (
            .O(N__9653),
            .I(N__9650));
    LocalMux I__966 (
            .O(N__9650),
            .I(\receive_module.rx_counter.n3400 ));
    SRMux I__965 (
            .O(N__9647),
            .I(N__9644));
    LocalMux I__964 (
            .O(N__9644),
            .I(N__9641));
    Span4Mux_v I__963 (
            .O(N__9641),
            .I(N__9637));
    SRMux I__962 (
            .O(N__9640),
            .I(N__9633));
    Span4Mux_v I__961 (
            .O(N__9637),
            .I(N__9630));
    SRMux I__960 (
            .O(N__9636),
            .I(N__9627));
    LocalMux I__959 (
            .O(N__9633),
            .I(N__9624));
    Span4Mux_v I__958 (
            .O(N__9630),
            .I(N__9619));
    LocalMux I__957 (
            .O(N__9627),
            .I(N__9619));
    Span4Mux_v I__956 (
            .O(N__9624),
            .I(N__9613));
    Span4Mux_v I__955 (
            .O(N__9619),
            .I(N__9613));
    SRMux I__954 (
            .O(N__9618),
            .I(N__9610));
    Sp12to4 I__953 (
            .O(N__9613),
            .I(N__9605));
    LocalMux I__952 (
            .O(N__9610),
            .I(N__9605));
    Odrv12 I__951 (
            .O(N__9605),
            .I(\line_buffer.n565 ));
    InMux I__950 (
            .O(N__9602),
            .I(N__9597));
    InMux I__949 (
            .O(N__9601),
            .I(N__9592));
    InMux I__948 (
            .O(N__9600),
            .I(N__9592));
    LocalMux I__947 (
            .O(N__9597),
            .I(\receive_module.rx_counter.X_5 ));
    LocalMux I__946 (
            .O(N__9592),
            .I(\receive_module.rx_counter.X_5 ));
    InMux I__945 (
            .O(N__9587),
            .I(N__9582));
    InMux I__944 (
            .O(N__9586),
            .I(N__9577));
    InMux I__943 (
            .O(N__9585),
            .I(N__9577));
    LocalMux I__942 (
            .O(N__9582),
            .I(\receive_module.rx_counter.X_4 ));
    LocalMux I__941 (
            .O(N__9577),
            .I(\receive_module.rx_counter.X_4 ));
    InMux I__940 (
            .O(N__9572),
            .I(N__9567));
    InMux I__939 (
            .O(N__9571),
            .I(N__9562));
    InMux I__938 (
            .O(N__9570),
            .I(N__9562));
    LocalMux I__937 (
            .O(N__9567),
            .I(\receive_module.rx_counter.X_3 ));
    LocalMux I__936 (
            .O(N__9562),
            .I(\receive_module.rx_counter.X_3 ));
    InMux I__935 (
            .O(N__9557),
            .I(N__9552));
    InMux I__934 (
            .O(N__9556),
            .I(N__9547));
    InMux I__933 (
            .O(N__9555),
            .I(N__9547));
    LocalMux I__932 (
            .O(N__9552),
            .I(\receive_module.rx_counter.X_6 ));
    LocalMux I__931 (
            .O(N__9547),
            .I(\receive_module.rx_counter.X_6 ));
    CascadeMux I__930 (
            .O(N__9542),
            .I(\receive_module.rx_counter.n6_cascade_ ));
    InMux I__929 (
            .O(N__9539),
            .I(N__9534));
    InMux I__928 (
            .O(N__9538),
            .I(N__9529));
    InMux I__927 (
            .O(N__9537),
            .I(N__9529));
    LocalMux I__926 (
            .O(N__9534),
            .I(\receive_module.rx_counter.X_7 ));
    LocalMux I__925 (
            .O(N__9529),
            .I(\receive_module.rx_counter.X_7 ));
    InMux I__924 (
            .O(N__9524),
            .I(N__9521));
    LocalMux I__923 (
            .O(N__9521),
            .I(\receive_module.rx_counter.n3385 ));
    InMux I__922 (
            .O(N__9518),
            .I(N__9515));
    LocalMux I__921 (
            .O(N__9515),
            .I(N__9512));
    Odrv4 I__920 (
            .O(N__9512),
            .I(\receive_module.rx_counter.old_HS ));
    InMux I__919 (
            .O(N__9509),
            .I(N__9505));
    InMux I__918 (
            .O(N__9508),
            .I(N__9501));
    LocalMux I__917 (
            .O(N__9505),
            .I(N__9498));
    InMux I__916 (
            .O(N__9504),
            .I(N__9495));
    LocalMux I__915 (
            .O(N__9501),
            .I(TVP_HSYNC_buff));
    Odrv4 I__914 (
            .O(N__9498),
            .I(TVP_HSYNC_buff));
    LocalMux I__913 (
            .O(N__9495),
            .I(TVP_HSYNC_buff));
    InMux I__912 (
            .O(N__9488),
            .I(bfn_12_11_0_));
    InMux I__911 (
            .O(N__9485),
            .I(\receive_module.n3091 ));
    InMux I__910 (
            .O(N__9482),
            .I(\receive_module.n3092 ));
    IoInMux I__909 (
            .O(N__9479),
            .I(N__9476));
    LocalMux I__908 (
            .O(N__9476),
            .I(N__9473));
    Span4Mux_s2_h I__907 (
            .O(N__9473),
            .I(N__9470));
    Span4Mux_h I__906 (
            .O(N__9470),
            .I(N__9466));
    InMux I__905 (
            .O(N__9469),
            .I(N__9463));
    Span4Mux_h I__904 (
            .O(N__9466),
            .I(N__9458));
    LocalMux I__903 (
            .O(N__9463),
            .I(N__9458));
    Span4Mux_h I__902 (
            .O(N__9458),
            .I(N__9455));
    Span4Mux_v I__901 (
            .O(N__9455),
            .I(N__9452));
    Odrv4 I__900 (
            .O(N__9452),
            .I(DEBUG_c_0_c));
    InMux I__899 (
            .O(N__9449),
            .I(N__9446));
    LocalMux I__898 (
            .O(N__9446),
            .I(\TVP_VSYNC_buff_I_0.BUFFER_0_0 ));
    InMux I__897 (
            .O(N__9443),
            .I(N__9439));
    InMux I__896 (
            .O(N__9442),
            .I(N__9436));
    LocalMux I__895 (
            .O(N__9439),
            .I(\receive_module.rx_counter.X_8 ));
    LocalMux I__894 (
            .O(N__9436),
            .I(\receive_module.rx_counter.X_8 ));
    CascadeMux I__893 (
            .O(N__9431),
            .I(N__9427));
    InMux I__892 (
            .O(N__9430),
            .I(N__9424));
    InMux I__891 (
            .O(N__9427),
            .I(N__9421));
    LocalMux I__890 (
            .O(N__9424),
            .I(\receive_module.rx_counter.X_9 ));
    LocalMux I__889 (
            .O(N__9421),
            .I(\receive_module.rx_counter.X_9 ));
    SRMux I__888 (
            .O(N__9416),
            .I(N__9412));
    SRMux I__887 (
            .O(N__9415),
            .I(N__9409));
    LocalMux I__886 (
            .O(N__9412),
            .I(N__9406));
    LocalMux I__885 (
            .O(N__9409),
            .I(N__9403));
    Sp12to4 I__884 (
            .O(N__9406),
            .I(N__9400));
    Span4Mux_h I__883 (
            .O(N__9403),
            .I(N__9397));
    Odrv12 I__882 (
            .O(N__9400),
            .I(\receive_module.rx_counter.n3630 ));
    Odrv4 I__881 (
            .O(N__9397),
            .I(\receive_module.rx_counter.n3630 ));
    InMux I__880 (
            .O(N__9392),
            .I(N__9389));
    LocalMux I__879 (
            .O(N__9389),
            .I(N__9386));
    Odrv4 I__878 (
            .O(N__9386),
            .I(\TVP_VSYNC_buff_I_0.BUFFER_1_0 ));
    SRMux I__877 (
            .O(N__9383),
            .I(N__9379));
    SRMux I__876 (
            .O(N__9382),
            .I(N__9376));
    LocalMux I__875 (
            .O(N__9379),
            .I(N__9370));
    LocalMux I__874 (
            .O(N__9376),
            .I(N__9370));
    SRMux I__873 (
            .O(N__9375),
            .I(N__9367));
    Span4Mux_v I__872 (
            .O(N__9370),
            .I(N__9362));
    LocalMux I__871 (
            .O(N__9367),
            .I(N__9362));
    Span4Mux_h I__870 (
            .O(N__9362),
            .I(N__9358));
    SRMux I__869 (
            .O(N__9361),
            .I(N__9355));
    Span4Mux_v I__868 (
            .O(N__9358),
            .I(N__9352));
    LocalMux I__867 (
            .O(N__9355),
            .I(N__9349));
    Span4Mux_v I__866 (
            .O(N__9352),
            .I(N__9346));
    Span4Mux_v I__865 (
            .O(N__9349),
            .I(N__9343));
    Span4Mux_v I__864 (
            .O(N__9346),
            .I(N__9340));
    Sp12to4 I__863 (
            .O(N__9343),
            .I(N__9337));
    Span4Mux_v I__862 (
            .O(N__9340),
            .I(N__9334));
    Span12Mux_h I__861 (
            .O(N__9337),
            .I(N__9331));
    Odrv4 I__860 (
            .O(N__9334),
            .I(\line_buffer.n467 ));
    Odrv12 I__859 (
            .O(N__9331),
            .I(\line_buffer.n467 ));
    InMux I__858 (
            .O(N__9326),
            .I(N__9323));
    LocalMux I__857 (
            .O(N__9323),
            .I(\transmit_module.Y_DELTA_PATTERN_43 ));
    InMux I__856 (
            .O(N__9320),
            .I(N__9317));
    LocalMux I__855 (
            .O(N__9317),
            .I(N__9314));
    Odrv12 I__854 (
            .O(N__9314),
            .I(\transmit_module.Y_DELTA_PATTERN_59 ));
    InMux I__853 (
            .O(N__9311),
            .I(N__9308));
    LocalMux I__852 (
            .O(N__9308),
            .I(\transmit_module.Y_DELTA_PATTERN_45 ));
    InMux I__851 (
            .O(N__9305),
            .I(N__9302));
    LocalMux I__850 (
            .O(N__9302),
            .I(\transmit_module.Y_DELTA_PATTERN_44 ));
    InMux I__849 (
            .O(N__9299),
            .I(N__9296));
    LocalMux I__848 (
            .O(N__9296),
            .I(N__9293));
    Odrv4 I__847 (
            .O(N__9293),
            .I(\transmit_module.Y_DELTA_PATTERN_47 ));
    InMux I__846 (
            .O(N__9290),
            .I(N__9287));
    LocalMux I__845 (
            .O(N__9287),
            .I(\transmit_module.Y_DELTA_PATTERN_46 ));
    InMux I__844 (
            .O(N__9284),
            .I(N__9281));
    LocalMux I__843 (
            .O(N__9281),
            .I(\transmit_module.Y_DELTA_PATTERN_61 ));
    InMux I__842 (
            .O(N__9278),
            .I(N__9275));
    LocalMux I__841 (
            .O(N__9275),
            .I(\transmit_module.Y_DELTA_PATTERN_60 ));
    InMux I__840 (
            .O(N__9272),
            .I(N__9269));
    LocalMux I__839 (
            .O(N__9269),
            .I(\transmit_module.Y_DELTA_PATTERN_77 ));
    InMux I__838 (
            .O(N__9266),
            .I(N__9263));
    LocalMux I__837 (
            .O(N__9263),
            .I(\transmit_module.Y_DELTA_PATTERN_76 ));
    CascadeMux I__836 (
            .O(N__9260),
            .I(N__9257));
    CascadeBuf I__835 (
            .O(N__9257),
            .I(N__9253));
    CascadeMux I__834 (
            .O(N__9256),
            .I(N__9250));
    CascadeMux I__833 (
            .O(N__9253),
            .I(N__9247));
    CascadeBuf I__832 (
            .O(N__9250),
            .I(N__9244));
    CascadeBuf I__831 (
            .O(N__9247),
            .I(N__9241));
    CascadeMux I__830 (
            .O(N__9244),
            .I(N__9238));
    CascadeMux I__829 (
            .O(N__9241),
            .I(N__9235));
    CascadeBuf I__828 (
            .O(N__9238),
            .I(N__9232));
    CascadeBuf I__827 (
            .O(N__9235),
            .I(N__9229));
    CascadeMux I__826 (
            .O(N__9232),
            .I(N__9226));
    CascadeMux I__825 (
            .O(N__9229),
            .I(N__9223));
    CascadeBuf I__824 (
            .O(N__9226),
            .I(N__9220));
    CascadeBuf I__823 (
            .O(N__9223),
            .I(N__9217));
    CascadeMux I__822 (
            .O(N__9220),
            .I(N__9214));
    CascadeMux I__821 (
            .O(N__9217),
            .I(N__9211));
    CascadeBuf I__820 (
            .O(N__9214),
            .I(N__9208));
    CascadeBuf I__819 (
            .O(N__9211),
            .I(N__9205));
    CascadeMux I__818 (
            .O(N__9208),
            .I(N__9202));
    CascadeMux I__817 (
            .O(N__9205),
            .I(N__9199));
    CascadeBuf I__816 (
            .O(N__9202),
            .I(N__9196));
    CascadeBuf I__815 (
            .O(N__9199),
            .I(N__9193));
    CascadeMux I__814 (
            .O(N__9196),
            .I(N__9190));
    CascadeMux I__813 (
            .O(N__9193),
            .I(N__9187));
    CascadeBuf I__812 (
            .O(N__9190),
            .I(N__9184));
    CascadeBuf I__811 (
            .O(N__9187),
            .I(N__9181));
    CascadeMux I__810 (
            .O(N__9184),
            .I(N__9178));
    CascadeMux I__809 (
            .O(N__9181),
            .I(N__9175));
    CascadeBuf I__808 (
            .O(N__9178),
            .I(N__9172));
    CascadeBuf I__807 (
            .O(N__9175),
            .I(N__9169));
    CascadeMux I__806 (
            .O(N__9172),
            .I(N__9166));
    CascadeMux I__805 (
            .O(N__9169),
            .I(N__9163));
    CascadeBuf I__804 (
            .O(N__9166),
            .I(N__9160));
    CascadeBuf I__803 (
            .O(N__9163),
            .I(N__9157));
    CascadeMux I__802 (
            .O(N__9160),
            .I(N__9154));
    CascadeMux I__801 (
            .O(N__9157),
            .I(N__9151));
    CascadeBuf I__800 (
            .O(N__9154),
            .I(N__9148));
    CascadeBuf I__799 (
            .O(N__9151),
            .I(N__9145));
    CascadeMux I__798 (
            .O(N__9148),
            .I(N__9142));
    CascadeMux I__797 (
            .O(N__9145),
            .I(N__9139));
    CascadeBuf I__796 (
            .O(N__9142),
            .I(N__9136));
    CascadeBuf I__795 (
            .O(N__9139),
            .I(N__9133));
    CascadeMux I__794 (
            .O(N__9136),
            .I(N__9130));
    CascadeMux I__793 (
            .O(N__9133),
            .I(N__9127));
    CascadeBuf I__792 (
            .O(N__9130),
            .I(N__9124));
    CascadeBuf I__791 (
            .O(N__9127),
            .I(N__9121));
    CascadeMux I__790 (
            .O(N__9124),
            .I(N__9118));
    CascadeMux I__789 (
            .O(N__9121),
            .I(N__9115));
    CascadeBuf I__788 (
            .O(N__9118),
            .I(N__9112));
    CascadeBuf I__787 (
            .O(N__9115),
            .I(N__9109));
    CascadeMux I__786 (
            .O(N__9112),
            .I(N__9106));
    CascadeMux I__785 (
            .O(N__9109),
            .I(N__9103));
    CascadeBuf I__784 (
            .O(N__9106),
            .I(N__9100));
    CascadeBuf I__783 (
            .O(N__9103),
            .I(N__9097));
    CascadeMux I__782 (
            .O(N__9100),
            .I(N__9094));
    CascadeMux I__781 (
            .O(N__9097),
            .I(N__9091));
    CascadeBuf I__780 (
            .O(N__9094),
            .I(N__9088));
    CascadeBuf I__779 (
            .O(N__9091),
            .I(N__9085));
    CascadeMux I__778 (
            .O(N__9088),
            .I(N__9082));
    CascadeMux I__777 (
            .O(N__9085),
            .I(N__9079));
    CascadeBuf I__776 (
            .O(N__9082),
            .I(N__9076));
    InMux I__775 (
            .O(N__9079),
            .I(N__9073));
    CascadeMux I__774 (
            .O(N__9076),
            .I(N__9070));
    LocalMux I__773 (
            .O(N__9073),
            .I(N__9067));
    InMux I__772 (
            .O(N__9070),
            .I(N__9064));
    Span12Mux_h I__771 (
            .O(N__9067),
            .I(N__9061));
    LocalMux I__770 (
            .O(N__9064),
            .I(N__9058));
    Odrv12 I__769 (
            .O(N__9061),
            .I(n24));
    Odrv4 I__768 (
            .O(N__9058),
            .I(n24));
    InMux I__767 (
            .O(N__9053),
            .I(N__9050));
    LocalMux I__766 (
            .O(N__9050),
            .I(N__9047));
    Span4Mux_h I__765 (
            .O(N__9047),
            .I(N__9044));
    Odrv4 I__764 (
            .O(N__9044),
            .I(TVP_VIDEO_c_4));
    InMux I__763 (
            .O(N__9041),
            .I(N__9038));
    LocalMux I__762 (
            .O(N__9038),
            .I(\transmit_module.Y_DELTA_PATTERN_99 ));
    InMux I__761 (
            .O(N__9035),
            .I(N__9032));
    LocalMux I__760 (
            .O(N__9032),
            .I(\transmit_module.Y_DELTA_PATTERN_10 ));
    InMux I__759 (
            .O(N__9029),
            .I(N__9026));
    LocalMux I__758 (
            .O(N__9026),
            .I(\transmit_module.Y_DELTA_PATTERN_9 ));
    InMux I__757 (
            .O(N__9023),
            .I(N__9020));
    LocalMux I__756 (
            .O(N__9020),
            .I(\transmit_module.Y_DELTA_PATTERN_12 ));
    InMux I__755 (
            .O(N__9017),
            .I(N__9014));
    LocalMux I__754 (
            .O(N__9014),
            .I(\transmit_module.Y_DELTA_PATTERN_11 ));
    InMux I__753 (
            .O(N__9011),
            .I(N__9008));
    LocalMux I__752 (
            .O(N__9008),
            .I(N__9005));
    Odrv4 I__751 (
            .O(N__9005),
            .I(\transmit_module.Y_DELTA_PATTERN_38 ));
    InMux I__750 (
            .O(N__9002),
            .I(N__8999));
    LocalMux I__749 (
            .O(N__8999),
            .I(\transmit_module.Y_DELTA_PATTERN_40 ));
    InMux I__748 (
            .O(N__8996),
            .I(N__8993));
    LocalMux I__747 (
            .O(N__8993),
            .I(\transmit_module.Y_DELTA_PATTERN_39 ));
    InMux I__746 (
            .O(N__8990),
            .I(N__8987));
    LocalMux I__745 (
            .O(N__8987),
            .I(\transmit_module.Y_DELTA_PATTERN_41 ));
    InMux I__744 (
            .O(N__8984),
            .I(N__8981));
    LocalMux I__743 (
            .O(N__8981),
            .I(\transmit_module.Y_DELTA_PATTERN_42 ));
    InMux I__742 (
            .O(N__8978),
            .I(N__8975));
    LocalMux I__741 (
            .O(N__8975),
            .I(\transmit_module.Y_DELTA_PATTERN_24 ));
    InMux I__740 (
            .O(N__8972),
            .I(N__8969));
    LocalMux I__739 (
            .O(N__8969),
            .I(\transmit_module.Y_DELTA_PATTERN_23 ));
    InMux I__738 (
            .O(N__8966),
            .I(N__8963));
    LocalMux I__737 (
            .O(N__8963),
            .I(\transmit_module.Y_DELTA_PATTERN_28 ));
    InMux I__736 (
            .O(N__8960),
            .I(N__8957));
    LocalMux I__735 (
            .O(N__8957),
            .I(\transmit_module.Y_DELTA_PATTERN_27 ));
    InMux I__734 (
            .O(N__8954),
            .I(N__8951));
    LocalMux I__733 (
            .O(N__8951),
            .I(\transmit_module.Y_DELTA_PATTERN_13 ));
    InMux I__732 (
            .O(N__8948),
            .I(N__8945));
    LocalMux I__731 (
            .O(N__8945),
            .I(\transmit_module.Y_DELTA_PATTERN_15 ));
    InMux I__730 (
            .O(N__8942),
            .I(N__8939));
    LocalMux I__729 (
            .O(N__8939),
            .I(\transmit_module.Y_DELTA_PATTERN_14 ));
    InMux I__728 (
            .O(N__8936),
            .I(N__8933));
    LocalMux I__727 (
            .O(N__8933),
            .I(\transmit_module.Y_DELTA_PATTERN_26 ));
    InMux I__726 (
            .O(N__8930),
            .I(N__8927));
    LocalMux I__725 (
            .O(N__8927),
            .I(\transmit_module.Y_DELTA_PATTERN_25 ));
    InMux I__724 (
            .O(N__8924),
            .I(N__8921));
    LocalMux I__723 (
            .O(N__8921),
            .I(\transmit_module.Y_DELTA_PATTERN_8 ));
    InMux I__722 (
            .O(N__8918),
            .I(N__8915));
    LocalMux I__721 (
            .O(N__8915),
            .I(\transmit_module.Y_DELTA_PATTERN_50 ));
    InMux I__720 (
            .O(N__8912),
            .I(N__8909));
    LocalMux I__719 (
            .O(N__8909),
            .I(\transmit_module.Y_DELTA_PATTERN_51 ));
    InMux I__718 (
            .O(N__8906),
            .I(N__8903));
    LocalMux I__717 (
            .O(N__8903),
            .I(\transmit_module.Y_DELTA_PATTERN_58 ));
    InMux I__716 (
            .O(N__8900),
            .I(N__8897));
    LocalMux I__715 (
            .O(N__8897),
            .I(\transmit_module.Y_DELTA_PATTERN_57 ));
    InMux I__714 (
            .O(N__8894),
            .I(N__8891));
    LocalMux I__713 (
            .O(N__8891),
            .I(\transmit_module.Y_DELTA_PATTERN_22 ));
    InMux I__712 (
            .O(N__8888),
            .I(N__8885));
    LocalMux I__711 (
            .O(N__8885),
            .I(\transmit_module.Y_DELTA_PATTERN_21 ));
    InMux I__710 (
            .O(N__8882),
            .I(N__8879));
    LocalMux I__709 (
            .O(N__8879),
            .I(\receive_module.rx_counter.n9_adj_612 ));
    InMux I__708 (
            .O(N__8876),
            .I(\receive_module.rx_counter.n3147 ));
    InMux I__707 (
            .O(N__8873),
            .I(N__8870));
    LocalMux I__706 (
            .O(N__8870),
            .I(\receive_module.rx_counter.n8_adj_611 ));
    InMux I__705 (
            .O(N__8867),
            .I(\receive_module.rx_counter.n3148 ));
    InMux I__704 (
            .O(N__8864),
            .I(\receive_module.rx_counter.n3149 ));
    InMux I__703 (
            .O(N__8861),
            .I(\receive_module.rx_counter.n3150 ));
    InMux I__702 (
            .O(N__8858),
            .I(\receive_module.rx_counter.n3151 ));
    InMux I__701 (
            .O(N__8855),
            .I(\receive_module.rx_counter.n3152 ));
    InMux I__700 (
            .O(N__8852),
            .I(\receive_module.rx_counter.n3153 ));
    InMux I__699 (
            .O(N__8849),
            .I(bfn_11_10_0_));
    InMux I__698 (
            .O(N__8846),
            .I(\receive_module.rx_counter.n3155 ));
    InMux I__697 (
            .O(N__8843),
            .I(N__8840));
    LocalMux I__696 (
            .O(N__8840),
            .I(\transmit_module.Y_DELTA_PATTERN_75 ));
    InMux I__695 (
            .O(N__8837),
            .I(N__8834));
    LocalMux I__694 (
            .O(N__8834),
            .I(\transmit_module.Y_DELTA_PATTERN_62 ));
    InMux I__693 (
            .O(N__8831),
            .I(N__8828));
    LocalMux I__692 (
            .O(N__8828),
            .I(N__8825));
    Odrv4 I__691 (
            .O(N__8825),
            .I(\transmit_module.Y_DELTA_PATTERN_78 ));
    InMux I__690 (
            .O(N__8822),
            .I(N__8819));
    LocalMux I__689 (
            .O(N__8819),
            .I(\tvp_video_buffer.BUFFER_0_2 ));
    IoInMux I__688 (
            .O(N__8816),
            .I(N__8813));
    LocalMux I__687 (
            .O(N__8813),
            .I(N__8810));
    Span12Mux_s6_v I__686 (
            .O(N__8810),
            .I(N__8806));
    InMux I__685 (
            .O(N__8809),
            .I(N__8803));
    Odrv12 I__684 (
            .O(N__8806),
            .I(LED_c));
    LocalMux I__683 (
            .O(N__8803),
            .I(LED_c));
    IoInMux I__682 (
            .O(N__8798),
            .I(N__8795));
    LocalMux I__681 (
            .O(N__8795),
            .I(N__8792));
    IoSpan4Mux I__680 (
            .O(N__8792),
            .I(N__8789));
    Span4Mux_s3_h I__679 (
            .O(N__8789),
            .I(N__8785));
    InMux I__678 (
            .O(N__8788),
            .I(N__8782));
    Span4Mux_h I__677 (
            .O(N__8785),
            .I(N__8779));
    LocalMux I__676 (
            .O(N__8782),
            .I(N__8776));
    Span4Mux_h I__675 (
            .O(N__8779),
            .I(N__8771));
    Span4Mux_v I__674 (
            .O(N__8776),
            .I(N__8771));
    Span4Mux_h I__673 (
            .O(N__8771),
            .I(N__8768));
    Span4Mux_h I__672 (
            .O(N__8768),
            .I(N__8765));
    Odrv4 I__671 (
            .O(N__8765),
            .I(DEBUG_c_1_c));
    InMux I__670 (
            .O(N__8762),
            .I(N__8759));
    LocalMux I__669 (
            .O(N__8759),
            .I(\tvp_hs_buffer.BUFFER_0_0 ));
    InMux I__668 (
            .O(N__8756),
            .I(N__8753));
    LocalMux I__667 (
            .O(N__8753),
            .I(\tvp_hs_buffer.BUFFER_1_0 ));
    InMux I__666 (
            .O(N__8750),
            .I(N__8747));
    LocalMux I__665 (
            .O(N__8747),
            .I(\receive_module.rx_counter.n10 ));
    InMux I__664 (
            .O(N__8744),
            .I(bfn_11_9_0_));
    InMux I__663 (
            .O(N__8741),
            .I(N__8738));
    LocalMux I__662 (
            .O(N__8738),
            .I(N__8735));
    Odrv4 I__661 (
            .O(N__8735),
            .I(\transmit_module.Y_DELTA_PATTERN_33 ));
    InMux I__660 (
            .O(N__8732),
            .I(N__8729));
    LocalMux I__659 (
            .O(N__8729),
            .I(\transmit_module.Y_DELTA_PATTERN_29 ));
    InMux I__658 (
            .O(N__8726),
            .I(N__8723));
    LocalMux I__657 (
            .O(N__8723),
            .I(\transmit_module.Y_DELTA_PATTERN_32 ));
    InMux I__656 (
            .O(N__8720),
            .I(N__8717));
    LocalMux I__655 (
            .O(N__8717),
            .I(\transmit_module.Y_DELTA_PATTERN_31 ));
    InMux I__654 (
            .O(N__8714),
            .I(N__8711));
    LocalMux I__653 (
            .O(N__8711),
            .I(\transmit_module.Y_DELTA_PATTERN_30 ));
    InMux I__652 (
            .O(N__8708),
            .I(N__8705));
    LocalMux I__651 (
            .O(N__8705),
            .I(\transmit_module.Y_DELTA_PATTERN_74 ));
    InMux I__650 (
            .O(N__8702),
            .I(N__8699));
    LocalMux I__649 (
            .O(N__8699),
            .I(N__8696));
    Odrv4 I__648 (
            .O(N__8696),
            .I(\transmit_module.Y_DELTA_PATTERN_73 ));
    InMux I__647 (
            .O(N__8693),
            .I(N__8690));
    LocalMux I__646 (
            .O(N__8690),
            .I(\transmit_module.Y_DELTA_PATTERN_65 ));
    InMux I__645 (
            .O(N__8687),
            .I(N__8684));
    LocalMux I__644 (
            .O(N__8684),
            .I(\transmit_module.Y_DELTA_PATTERN_64 ));
    InMux I__643 (
            .O(N__8681),
            .I(N__8678));
    LocalMux I__642 (
            .O(N__8678),
            .I(\transmit_module.Y_DELTA_PATTERN_63 ));
    InMux I__641 (
            .O(N__8675),
            .I(N__8672));
    LocalMux I__640 (
            .O(N__8672),
            .I(\transmit_module.Y_DELTA_PATTERN_91 ));
    InMux I__639 (
            .O(N__8669),
            .I(N__8666));
    LocalMux I__638 (
            .O(N__8666),
            .I(\transmit_module.Y_DELTA_PATTERN_93 ));
    InMux I__637 (
            .O(N__8663),
            .I(N__8660));
    LocalMux I__636 (
            .O(N__8660),
            .I(\transmit_module.Y_DELTA_PATTERN_92 ));
    InMux I__635 (
            .O(N__8657),
            .I(N__8654));
    LocalMux I__634 (
            .O(N__8654),
            .I(\transmit_module.Y_DELTA_PATTERN_94 ));
    InMux I__633 (
            .O(N__8651),
            .I(N__8648));
    LocalMux I__632 (
            .O(N__8648),
            .I(\transmit_module.Y_DELTA_PATTERN_97 ));
    InMux I__631 (
            .O(N__8645),
            .I(N__8642));
    LocalMux I__630 (
            .O(N__8642),
            .I(\transmit_module.Y_DELTA_PATTERN_98 ));
    InMux I__629 (
            .O(N__8639),
            .I(N__8636));
    LocalMux I__628 (
            .O(N__8636),
            .I(\transmit_module.Y_DELTA_PATTERN_96 ));
    InMux I__627 (
            .O(N__8633),
            .I(N__8630));
    LocalMux I__626 (
            .O(N__8630),
            .I(\transmit_module.Y_DELTA_PATTERN_95 ));
    InMux I__625 (
            .O(N__8627),
            .I(N__8624));
    LocalMux I__624 (
            .O(N__8624),
            .I(N__8621));
    IoSpan4Mux I__623 (
            .O(N__8621),
            .I(N__8618));
    Odrv4 I__622 (
            .O(N__8618),
            .I(TVP_VIDEO_c_2));
    SRMux I__621 (
            .O(N__8615),
            .I(N__8610));
    SRMux I__620 (
            .O(N__8614),
            .I(N__8607));
    SRMux I__619 (
            .O(N__8613),
            .I(N__8604));
    LocalMux I__618 (
            .O(N__8610),
            .I(N__8600));
    LocalMux I__617 (
            .O(N__8607),
            .I(N__8595));
    LocalMux I__616 (
            .O(N__8604),
            .I(N__8595));
    SRMux I__615 (
            .O(N__8603),
            .I(N__8592));
    Span4Mux_h I__614 (
            .O(N__8600),
            .I(N__8589));
    Span4Mux_v I__613 (
            .O(N__8595),
            .I(N__8584));
    LocalMux I__612 (
            .O(N__8592),
            .I(N__8584));
    Sp12to4 I__611 (
            .O(N__8589),
            .I(N__8581));
    Span4Mux_v I__610 (
            .O(N__8584),
            .I(N__8578));
    Span12Mux_v I__609 (
            .O(N__8581),
            .I(N__8575));
    Span4Mux_h I__608 (
            .O(N__8578),
            .I(N__8572));
    Odrv12 I__607 (
            .O(N__8575),
            .I(\line_buffer.n533 ));
    Odrv4 I__606 (
            .O(N__8572),
            .I(\line_buffer.n533 ));
    InMux I__605 (
            .O(N__8567),
            .I(N__8564));
    LocalMux I__604 (
            .O(N__8564),
            .I(N__8561));
    Span4Mux_h I__603 (
            .O(N__8561),
            .I(N__8558));
    Odrv4 I__602 (
            .O(N__8558),
            .I(\tvp_video_buffer.BUFFER_0_3 ));
    InMux I__601 (
            .O(N__8555),
            .I(N__8552));
    LocalMux I__600 (
            .O(N__8552),
            .I(N__8549));
    Span4Mux_v I__599 (
            .O(N__8549),
            .I(N__8546));
    Odrv4 I__598 (
            .O(N__8546),
            .I(\transmit_module.Y_DELTA_PATTERN_82 ));
    InMux I__597 (
            .O(N__8543),
            .I(N__8540));
    LocalMux I__596 (
            .O(N__8540),
            .I(N__8537));
    Span4Mux_v I__595 (
            .O(N__8537),
            .I(N__8534));
    Odrv4 I__594 (
            .O(N__8534),
            .I(\transmit_module.Y_DELTA_PATTERN_49 ));
    InMux I__593 (
            .O(N__8531),
            .I(N__8528));
    LocalMux I__592 (
            .O(N__8528),
            .I(\transmit_module.Y_DELTA_PATTERN_84 ));
    InMux I__591 (
            .O(N__8525),
            .I(N__8522));
    LocalMux I__590 (
            .O(N__8522),
            .I(\transmit_module.Y_DELTA_PATTERN_83 ));
    InMux I__589 (
            .O(N__8519),
            .I(N__8516));
    LocalMux I__588 (
            .O(N__8516),
            .I(\transmit_module.Y_DELTA_PATTERN_85 ));
    InMux I__587 (
            .O(N__8513),
            .I(N__8510));
    LocalMux I__586 (
            .O(N__8510),
            .I(\transmit_module.Y_DELTA_PATTERN_87 ));
    InMux I__585 (
            .O(N__8507),
            .I(N__8504));
    LocalMux I__584 (
            .O(N__8504),
            .I(\transmit_module.Y_DELTA_PATTERN_86 ));
    InMux I__583 (
            .O(N__8501),
            .I(N__8498));
    LocalMux I__582 (
            .O(N__8498),
            .I(\transmit_module.Y_DELTA_PATTERN_81 ));
    InMux I__581 (
            .O(N__8495),
            .I(N__8492));
    LocalMux I__580 (
            .O(N__8492),
            .I(\transmit_module.Y_DELTA_PATTERN_80 ));
    InMux I__579 (
            .O(N__8489),
            .I(N__8486));
    LocalMux I__578 (
            .O(N__8486),
            .I(\transmit_module.Y_DELTA_PATTERN_37 ));
    InMux I__577 (
            .O(N__8483),
            .I(N__8480));
    LocalMux I__576 (
            .O(N__8480),
            .I(\transmit_module.Y_DELTA_PATTERN_79 ));
    InMux I__575 (
            .O(N__8477),
            .I(N__8474));
    LocalMux I__574 (
            .O(N__8474),
            .I(\transmit_module.Y_DELTA_PATTERN_66 ));
    InMux I__573 (
            .O(N__8471),
            .I(N__8468));
    LocalMux I__572 (
            .O(N__8468),
            .I(N__8465));
    Span4Mux_v I__571 (
            .O(N__8465),
            .I(N__8462));
    Odrv4 I__570 (
            .O(N__8462),
            .I(\transmit_module.Y_DELTA_PATTERN_69 ));
    InMux I__569 (
            .O(N__8459),
            .I(N__8456));
    LocalMux I__568 (
            .O(N__8456),
            .I(\transmit_module.Y_DELTA_PATTERN_68 ));
    InMux I__567 (
            .O(N__8453),
            .I(N__8450));
    LocalMux I__566 (
            .O(N__8450),
            .I(\transmit_module.Y_DELTA_PATTERN_67 ));
    InMux I__565 (
            .O(N__8447),
            .I(N__8444));
    LocalMux I__564 (
            .O(N__8444),
            .I(\transmit_module.Y_DELTA_PATTERN_48 ));
    InMux I__563 (
            .O(N__8441),
            .I(N__8438));
    LocalMux I__562 (
            .O(N__8438),
            .I(\transmit_module.Y_DELTA_PATTERN_34 ));
    InMux I__561 (
            .O(N__8435),
            .I(N__8432));
    LocalMux I__560 (
            .O(N__8432),
            .I(N__8429));
    Odrv4 I__559 (
            .O(N__8429),
            .I(\transmit_module.Y_DELTA_PATTERN_72 ));
    InMux I__558 (
            .O(N__8426),
            .I(N__8423));
    LocalMux I__557 (
            .O(N__8423),
            .I(\transmit_module.Y_DELTA_PATTERN_90 ));
    InMux I__556 (
            .O(N__8420),
            .I(N__8417));
    LocalMux I__555 (
            .O(N__8417),
            .I(\transmit_module.Y_DELTA_PATTERN_89 ));
    InMux I__554 (
            .O(N__8414),
            .I(N__8411));
    LocalMux I__553 (
            .O(N__8411),
            .I(\transmit_module.Y_DELTA_PATTERN_88 ));
    InMux I__552 (
            .O(N__8408),
            .I(N__8405));
    LocalMux I__551 (
            .O(N__8405),
            .I(N__8402));
    Odrv4 I__550 (
            .O(N__8402),
            .I(\transmit_module.Y_DELTA_PATTERN_36 ));
    IoInMux I__549 (
            .O(N__8399),
            .I(N__8396));
    LocalMux I__548 (
            .O(N__8396),
            .I(N__8392));
    IoInMux I__547 (
            .O(N__8395),
            .I(N__8389));
    IoSpan4Mux I__546 (
            .O(N__8392),
            .I(N__8386));
    LocalMux I__545 (
            .O(N__8389),
            .I(N__8383));
    Span4Mux_s3_v I__544 (
            .O(N__8386),
            .I(N__8380));
    Span4Mux_s2_h I__543 (
            .O(N__8383),
            .I(N__8377));
    Span4Mux_v I__542 (
            .O(N__8380),
            .I(N__8374));
    Sp12to4 I__541 (
            .O(N__8377),
            .I(N__8371));
    Sp12to4 I__540 (
            .O(N__8374),
            .I(N__8366));
    Span12Mux_v I__539 (
            .O(N__8371),
            .I(N__8366));
    Odrv12 I__538 (
            .O(N__8366),
            .I(GB_BUFFER_DEBUG_c_2_c_THRU_CO));
    InMux I__537 (
            .O(N__8363),
            .I(N__8360));
    LocalMux I__536 (
            .O(N__8360),
            .I(\transmit_module.Y_DELTA_PATTERN_70 ));
    InMux I__535 (
            .O(N__8357),
            .I(N__8354));
    LocalMux I__534 (
            .O(N__8354),
            .I(N__8351));
    Odrv12 I__533 (
            .O(N__8351),
            .I(TVP_VIDEO_c_3));
    InMux I__532 (
            .O(N__8348),
            .I(N__8345));
    LocalMux I__531 (
            .O(N__8345),
            .I(\transmit_module.Y_DELTA_PATTERN_71 ));
    InMux I__530 (
            .O(N__8342),
            .I(N__8339));
    LocalMux I__529 (
            .O(N__8339),
            .I(\transmit_module.Y_DELTA_PATTERN_35 ));
    INV \INVTVP_VSYNC_buff_I_0.WIRE_OUT_0__9C  (
            .O(\INVTVP_VSYNC_buff_I_0.WIRE_OUT_0__9C_net ),
            .I(N__24595));
    INV \INVTVP_VSYNC_buff_I_0.BUFFER_0__i2C  (
            .O(\INVTVP_VSYNC_buff_I_0.BUFFER_0__i2C_net ),
            .I(N__24586));
    INV \INVTVP_VSYNC_buff_I_0.BUFFER_0__i1C  (
            .O(\INVTVP_VSYNC_buff_I_0.BUFFER_0__i1C_net ),
            .I(N__24582));
    defparam IN_MUX_bfv_13_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_12_0_));
    defparam IN_MUX_bfv_13_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_13_0_ (
            .carryinitin(\transmit_module.video_signal_controller.n3143 ),
            .carryinitout(bfn_13_13_0_));
    defparam IN_MUX_bfv_12_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_15_0_));
    defparam IN_MUX_bfv_12_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_16_0_ (
            .carryinitin(\transmit_module.video_signal_controller.n3132 ),
            .carryinitout(bfn_12_16_0_));
    defparam IN_MUX_bfv_15_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_13_0_));
    defparam IN_MUX_bfv_15_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_14_0_ (
            .carryinitin(\transmit_module.n3111 ),
            .carryinitout(bfn_15_14_0_));
    defparam IN_MUX_bfv_13_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_9_0_));
    defparam IN_MUX_bfv_13_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_10_0_ (
            .carryinitin(\receive_module.rx_counter.n3124 ),
            .carryinitout(bfn_13_10_0_));
    defparam IN_MUX_bfv_11_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_9_0_));
    defparam IN_MUX_bfv_11_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_10_0_ (
            .carryinitin(\receive_module.rx_counter.n3154 ),
            .carryinitout(bfn_11_10_0_));
    defparam IN_MUX_bfv_13_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_6_0_));
    defparam IN_MUX_bfv_12_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_11_0_));
    defparam IN_MUX_bfv_12_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_12_0_ (
            .carryinitin(\receive_module.n3098 ),
            .carryinitout(bfn_12_12_0_));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam GB_BUFFER_DEBUG_c_2_c_THRU_LUT4_0_LC_3_25_4.C_ON=1'b0;
    defparam GB_BUFFER_DEBUG_c_2_c_THRU_LUT4_0_LC_3_25_4.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_DEBUG_c_2_c_THRU_LUT4_0_LC_3_25_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 GB_BUFFER_DEBUG_c_2_c_THRU_LUT4_0_LC_3_25_4 (
            .in0(N__24641),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(GB_BUFFER_DEBUG_c_2_c_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.Y_DELTA_PATTERN_i70_LC_6_15_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i70_LC_6_15_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i70_LC_6_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i70_LC_6_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8348),
            .lcout(\transmit_module.Y_DELTA_PATTERN_70 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23482),
            .ce(N__15257),
            .sr(N__20409));
    defparam \transmit_module.Y_DELTA_PATTERN_i69_LC_6_16_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i69_LC_6_16_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i69_LC_6_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i69_LC_6_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8363),
            .lcout(\transmit_module.Y_DELTA_PATTERN_69 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23500),
            .ce(N__15251),
            .sr(N__20285));
    defparam \tvp_video_buffer.BUFFER_0__i2_LC_7_9_0 .C_ON=1'b0;
    defparam \tvp_video_buffer.BUFFER_0__i2_LC_7_9_0 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.BUFFER_0__i2_LC_7_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.BUFFER_0__i2_LC_7_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8357),
            .lcout(\tvp_video_buffer.BUFFER_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24609),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.Y_DELTA_PATTERN_i71_LC_7_15_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i71_LC_7_15_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i71_LC_7_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i71_LC_7_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8435),
            .lcout(\transmit_module.Y_DELTA_PATTERN_71 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23457),
            .ce(N__15255),
            .sr(N__20354));
    defparam \transmit_module.Y_DELTA_PATTERN_i35_LC_7_16_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i35_LC_7_16_2 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i35_LC_7_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i35_LC_7_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8408),
            .lcout(\transmit_module.Y_DELTA_PATTERN_35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23317),
            .ce(N__15250),
            .sr(N__20298));
    defparam \transmit_module.Y_DELTA_PATTERN_i34_LC_7_16_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i34_LC_7_16_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i34_LC_7_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i34_LC_7_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8342),
            .lcout(\transmit_module.Y_DELTA_PATTERN_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23317),
            .ce(N__15250),
            .sr(N__20298));
    defparam \transmit_module.Y_DELTA_PATTERN_i33_LC_7_17_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i33_LC_7_17_2 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i33_LC_7_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i33_LC_7_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8441),
            .lcout(\transmit_module.Y_DELTA_PATTERN_33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23319),
            .ce(N__15248),
            .sr(N__20414));
    defparam \transmit_module.Y_DELTA_PATTERN_i72_LC_7_18_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i72_LC_7_18_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i72_LC_7_18_4 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i72_LC_7_18_4  (
            .in0(_gnd_net_),
            .in1(N__8702),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.Y_DELTA_PATTERN_72 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23316),
            .ce(N__15221),
            .sr(N__20385));
    defparam \transmit_module.Y_DELTA_PATTERN_i87_LC_9_13_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i87_LC_9_13_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i87_LC_9_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i87_LC_9_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8414),
            .lcout(\transmit_module.Y_DELTA_PATTERN_87 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23506),
            .ce(N__18406),
            .sr(N__20416));
    defparam \transmit_module.Y_DELTA_PATTERN_i89_LC_9_14_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i89_LC_9_14_2 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i89_LC_9_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i89_LC_9_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8426),
            .lcout(\transmit_module.Y_DELTA_PATTERN_89 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23498),
            .ce(N__18392),
            .sr(N__20327));
    defparam \transmit_module.Y_DELTA_PATTERN_i90_LC_9_14_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i90_LC_9_14_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i90_LC_9_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i90_LC_9_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8675),
            .lcout(\transmit_module.Y_DELTA_PATTERN_90 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23498),
            .ce(N__18392),
            .sr(N__20327));
    defparam \transmit_module.Y_DELTA_PATTERN_i88_LC_9_14_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i88_LC_9_14_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i88_LC_9_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i88_LC_9_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8420),
            .lcout(\transmit_module.Y_DELTA_PATTERN_88 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23498),
            .ce(N__18392),
            .sr(N__20327));
    defparam \transmit_module.Y_DELTA_PATTERN_i96_LC_9_15_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i96_LC_9_15_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i96_LC_9_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i96_LC_9_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8651),
            .lcout(\transmit_module.Y_DELTA_PATTERN_96 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23422),
            .ce(N__21047),
            .sr(N__20413));
    defparam \transmit_module.Y_DELTA_PATTERN_i36_LC_9_16_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i36_LC_9_16_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i36_LC_9_16_0 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i36_LC_9_16_0  (
            .in0(_gnd_net_),
            .in1(N__8489),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.Y_DELTA_PATTERN_36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23505),
            .ce(N__15256),
            .sr(N__20338));
    defparam \transmit_module.Y_DELTA_PATTERN_i79_LC_9_16_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i79_LC_9_16_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i79_LC_9_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i79_LC_9_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8495),
            .lcout(\transmit_module.Y_DELTA_PATTERN_79 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23505),
            .ce(N__15256),
            .sr(N__20338));
    defparam \transmit_module.Y_DELTA_PATTERN_i81_LC_9_16_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i81_LC_9_16_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i81_LC_9_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i81_LC_9_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8555),
            .lcout(\transmit_module.Y_DELTA_PATTERN_81 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23505),
            .ce(N__15256),
            .sr(N__20338));
    defparam \transmit_module.Y_DELTA_PATTERN_i80_LC_9_16_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i80_LC_9_16_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i80_LC_9_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i80_LC_9_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8501),
            .lcout(\transmit_module.Y_DELTA_PATTERN_80 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23505),
            .ce(N__15256),
            .sr(N__20338));
    defparam \transmit_module.Y_DELTA_PATTERN_i37_LC_9_17_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i37_LC_9_17_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i37_LC_9_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i37_LC_9_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9011),
            .lcout(\transmit_module.Y_DELTA_PATTERN_37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23435),
            .ce(N__15244),
            .sr(N__20393));
    defparam \transmit_module.Y_DELTA_PATTERN_i78_LC_9_17_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i78_LC_9_17_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i78_LC_9_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i78_LC_9_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8483),
            .lcout(\transmit_module.Y_DELTA_PATTERN_78 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23435),
            .ce(N__15244),
            .sr(N__20393));
    defparam \transmit_module.Y_DELTA_PATTERN_i66_LC_9_18_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i66_LC_9_18_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i66_LC_9_18_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i66_LC_9_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8453),
            .lcout(\transmit_module.Y_DELTA_PATTERN_66 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23372),
            .ce(N__15220),
            .sr(N__20384));
    defparam \transmit_module.Y_DELTA_PATTERN_i48_LC_9_18_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i48_LC_9_18_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i48_LC_9_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i48_LC_9_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8543),
            .lcout(\transmit_module.Y_DELTA_PATTERN_48 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23372),
            .ce(N__15220),
            .sr(N__20384));
    defparam \transmit_module.Y_DELTA_PATTERN_i65_LC_9_18_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i65_LC_9_18_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i65_LC_9_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i65_LC_9_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8477),
            .lcout(\transmit_module.Y_DELTA_PATTERN_65 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23372),
            .ce(N__15220),
            .sr(N__20384));
    defparam \transmit_module.Y_DELTA_PATTERN_i68_LC_9_18_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i68_LC_9_18_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i68_LC_9_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i68_LC_9_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8471),
            .lcout(\transmit_module.Y_DELTA_PATTERN_68 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23372),
            .ce(N__15220),
            .sr(N__20384));
    defparam \transmit_module.Y_DELTA_PATTERN_i67_LC_9_18_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i67_LC_9_18_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i67_LC_9_18_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i67_LC_9_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8459),
            .lcout(\transmit_module.Y_DELTA_PATTERN_67 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23372),
            .ce(N__15220),
            .sr(N__20384));
    defparam \transmit_module.Y_DELTA_PATTERN_i47_LC_9_18_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i47_LC_9_18_7 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i47_LC_9_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i47_LC_9_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8447),
            .lcout(\transmit_module.Y_DELTA_PATTERN_47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23372),
            .ce(N__15220),
            .sr(N__20384));
    defparam \tvp_video_buffer.BUFFER_0__i1_LC_10_4_0 .C_ON=1'b0;
    defparam \tvp_video_buffer.BUFFER_0__i1_LC_10_4_0 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.BUFFER_0__i1_LC_10_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.BUFFER_0__i1_LC_10_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8627),
            .lcout(\tvp_video_buffer.BUFFER_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24581),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_LC_10_9_5 .C_ON=1'b0;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_LC_10_9_5 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_LC_10_9_5 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \line_buffer.i1_2_lut_3_lut_4_lut_LC_10_9_5  (
            .in0(N__14812),
            .in1(N__14668),
            .in2(N__14575),
            .in3(N__14474),
            .lcout(\line_buffer.n533 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.BUFFER_0__i10_LC_10_10_4 .C_ON=1'b0;
    defparam \tvp_video_buffer.BUFFER_0__i10_LC_10_10_4 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.BUFFER_0__i10_LC_10_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.BUFFER_0__i10_LC_10_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8567),
            .lcout(\tvp_video_buffer.BUFFER_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24604),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.Y_DELTA_PATTERN_i82_LC_10_12_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i82_LC_10_12_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i82_LC_10_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i82_LC_10_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8525),
            .lcout(\transmit_module.Y_DELTA_PATTERN_82 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23516),
            .ce(N__15254),
            .sr(N__20336));
    defparam \transmit_module.Y_DELTA_PATTERN_i49_LC_10_12_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i49_LC_10_12_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i49_LC_10_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i49_LC_10_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8918),
            .lcout(\transmit_module.Y_DELTA_PATTERN_49 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23516),
            .ce(N__15254),
            .sr(N__20336));
    defparam \transmit_module.Y_DELTA_PATTERN_i84_LC_10_13_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i84_LC_10_13_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i84_LC_10_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i84_LC_10_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8519),
            .lcout(\transmit_module.Y_DELTA_PATTERN_84 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23455),
            .ce(N__18407),
            .sr(N__20295));
    defparam \transmit_module.Y_DELTA_PATTERN_i83_LC_10_13_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i83_LC_10_13_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i83_LC_10_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i83_LC_10_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8531),
            .lcout(\transmit_module.Y_DELTA_PATTERN_83 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23455),
            .ce(N__18407),
            .sr(N__20295));
    defparam \transmit_module.Y_DELTA_PATTERN_i85_LC_10_13_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i85_LC_10_13_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i85_LC_10_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i85_LC_10_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8507),
            .lcout(\transmit_module.Y_DELTA_PATTERN_85 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23455),
            .ce(N__18407),
            .sr(N__20295));
    defparam \transmit_module.Y_DELTA_PATTERN_i86_LC_10_13_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i86_LC_10_13_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i86_LC_10_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i86_LC_10_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8513),
            .lcout(\transmit_module.Y_DELTA_PATTERN_86 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23455),
            .ce(N__18407),
            .sr(N__20295));
    defparam \transmit_module.Y_DELTA_PATTERN_i93_LC_10_14_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i93_LC_10_14_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i93_LC_10_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i93_LC_10_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8657),
            .lcout(\transmit_module.Y_DELTA_PATTERN_93 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23458),
            .ce(N__18402),
            .sr(N__20284));
    defparam \transmit_module.Y_DELTA_PATTERN_i91_LC_10_14_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i91_LC_10_14_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i91_LC_10_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i91_LC_10_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8663),
            .lcout(\transmit_module.Y_DELTA_PATTERN_91 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23458),
            .ce(N__18402),
            .sr(N__20284));
    defparam \transmit_module.Y_DELTA_PATTERN_i92_LC_10_14_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i92_LC_10_14_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i92_LC_10_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i92_LC_10_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8669),
            .lcout(\transmit_module.Y_DELTA_PATTERN_92 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23458),
            .ce(N__18402),
            .sr(N__20284));
    defparam \transmit_module.Y_DELTA_PATTERN_i94_LC_10_15_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i94_LC_10_15_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i94_LC_10_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i94_LC_10_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8633),
            .lcout(\transmit_module.Y_DELTA_PATTERN_94 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23303),
            .ce(N__18391),
            .sr(N__20293));
    defparam \transmit_module.Y_DELTA_PATTERN_i97_LC_10_15_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i97_LC_10_15_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i97_LC_10_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i97_LC_10_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8645),
            .lcout(\transmit_module.Y_DELTA_PATTERN_97 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23303),
            .ce(N__18391),
            .sr(N__20293));
    defparam \transmit_module.Y_DELTA_PATTERN_i98_LC_10_15_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i98_LC_10_15_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i98_LC_10_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i98_LC_10_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9041),
            .lcout(\transmit_module.Y_DELTA_PATTERN_98 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23303),
            .ce(N__18391),
            .sr(N__20293));
    defparam \transmit_module.Y_DELTA_PATTERN_i95_LC_10_15_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i95_LC_10_15_7 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i95_LC_10_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i95_LC_10_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8639),
            .lcout(\transmit_module.Y_DELTA_PATTERN_95 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23303),
            .ce(N__18391),
            .sr(N__20293));
    defparam \transmit_module.Y_DELTA_PATTERN_i28_LC_10_16_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i28_LC_10_16_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i28_LC_10_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i28_LC_10_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8732),
            .lcout(\transmit_module.Y_DELTA_PATTERN_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23468),
            .ce(N__21032),
            .sr(N__20337));
    defparam \transmit_module.Y_DELTA_PATTERN_i7_LC_10_16_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i7_LC_10_16_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i7_LC_10_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i7_LC_10_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8924),
            .lcout(\transmit_module.Y_DELTA_PATTERN_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23468),
            .ce(N__21032),
            .sr(N__20337));
    defparam \transmit_module.Y_DELTA_PATTERN_i32_LC_10_17_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i32_LC_10_17_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i32_LC_10_17_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i32_LC_10_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8741),
            .lcout(\transmit_module.Y_DELTA_PATTERN_32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23436),
            .ce(N__21022),
            .sr(N__20397));
    defparam \transmit_module.Y_DELTA_PATTERN_i29_LC_10_17_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i29_LC_10_17_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i29_LC_10_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i29_LC_10_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8714),
            .lcout(\transmit_module.Y_DELTA_PATTERN_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23436),
            .ce(N__21022),
            .sr(N__20397));
    defparam \transmit_module.Y_DELTA_PATTERN_i31_LC_10_17_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i31_LC_10_17_2 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i31_LC_10_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i31_LC_10_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8726),
            .lcout(\transmit_module.Y_DELTA_PATTERN_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23436),
            .ce(N__21022),
            .sr(N__20397));
    defparam \transmit_module.Y_DELTA_PATTERN_i30_LC_10_17_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i30_LC_10_17_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i30_LC_10_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i30_LC_10_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8720),
            .lcout(\transmit_module.Y_DELTA_PATTERN_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23436),
            .ce(N__21022),
            .sr(N__20397));
    defparam \transmit_module.Y_DELTA_PATTERN_i74_LC_10_18_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i74_LC_10_18_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i74_LC_10_18_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i74_LC_10_18_1  (
            .in0(N__8843),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.Y_DELTA_PATTERN_74 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23376),
            .ce(N__15164),
            .sr(N__20267));
    defparam \transmit_module.Y_DELTA_PATTERN_i73_LC_10_18_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i73_LC_10_18_2 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i73_LC_10_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i73_LC_10_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8708),
            .lcout(\transmit_module.Y_DELTA_PATTERN_73 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23376),
            .ce(N__15164),
            .sr(N__20267));
    defparam \transmit_module.Y_DELTA_PATTERN_i64_LC_10_18_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i64_LC_10_18_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i64_LC_10_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i64_LC_10_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8693),
            .lcout(\transmit_module.Y_DELTA_PATTERN_64 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23376),
            .ce(N__15164),
            .sr(N__20267));
    defparam \transmit_module.Y_DELTA_PATTERN_i62_LC_10_19_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i62_LC_10_19_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i62_LC_10_19_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i62_LC_10_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8681),
            .lcout(\transmit_module.Y_DELTA_PATTERN_62 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23161),
            .ce(N__15240),
            .sr(N__20297));
    defparam \transmit_module.Y_DELTA_PATTERN_i63_LC_10_19_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i63_LC_10_19_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i63_LC_10_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i63_LC_10_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8687),
            .lcout(\transmit_module.Y_DELTA_PATTERN_63 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23161),
            .ce(N__15240),
            .sr(N__20297));
    defparam \transmit_module.Y_DELTA_PATTERN_i75_LC_10_19_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i75_LC_10_19_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i75_LC_10_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i75_LC_10_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9266),
            .lcout(\transmit_module.Y_DELTA_PATTERN_75 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23161),
            .ce(N__15240),
            .sr(N__20297));
    defparam \transmit_module.Y_DELTA_PATTERN_i61_LC_10_19_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i61_LC_10_19_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i61_LC_10_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i61_LC_10_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8837),
            .lcout(\transmit_module.Y_DELTA_PATTERN_61 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23161),
            .ce(N__15240),
            .sr(N__20297));
    defparam \transmit_module.Y_DELTA_PATTERN_i77_LC_10_19_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i77_LC_10_19_7 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i77_LC_10_19_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i77_LC_10_19_7  (
            .in0(N__8831),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.Y_DELTA_PATTERN_77 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23161),
            .ce(N__15240),
            .sr(N__20297));
    defparam \tvp_video_buffer.BUFFER_0__i9_LC_11_4_5 .C_ON=1'b0;
    defparam \tvp_video_buffer.BUFFER_0__i9_LC_11_4_5 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.BUFFER_0__i9_LC_11_4_5 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \tvp_video_buffer.BUFFER_0__i9_LC_11_4_5  (
            .in0(_gnd_net_),
            .in1(N__8822),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\tvp_video_buffer.BUFFER_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24575),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.PULSE_1HZ_49_LC_11_7_5 .C_ON=1'b0;
    defparam \receive_module.rx_counter.PULSE_1HZ_49_LC_11_7_5 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.PULSE_1HZ_49_LC_11_7_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \receive_module.rx_counter.PULSE_1HZ_49_LC_11_7_5  (
            .in0(_gnd_net_),
            .in1(N__8809),
            .in2(_gnd_net_),
            .in3(N__12530),
            .lcout(LED_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24590),
            .ce(N__12622),
            .sr(_gnd_net_));
    defparam \tvp_hs_buffer.BUFFER_0__i2_LC_11_8_0 .C_ON=1'b0;
    defparam \tvp_hs_buffer.BUFFER_0__i2_LC_11_8_0 .SEQ_MODE=4'b1000;
    defparam \tvp_hs_buffer.BUFFER_0__i2_LC_11_8_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_hs_buffer.BUFFER_0__i2_LC_11_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8762),
            .lcout(\tvp_hs_buffer.BUFFER_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24594),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_hs_buffer.BUFFER_0__i1_LC_11_8_2 .C_ON=1'b0;
    defparam \tvp_hs_buffer.BUFFER_0__i1_LC_11_8_2 .SEQ_MODE=4'b1000;
    defparam \tvp_hs_buffer.BUFFER_0__i1_LC_11_8_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_hs_buffer.BUFFER_0__i1_LC_11_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8788),
            .lcout(\tvp_hs_buffer.BUFFER_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24594),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_hs_buffer.WIRE_OUT_0__9_LC_11_8_3 .C_ON=1'b0;
    defparam \tvp_hs_buffer.WIRE_OUT_0__9_LC_11_8_3 .SEQ_MODE=4'b1000;
    defparam \tvp_hs_buffer.WIRE_OUT_0__9_LC_11_8_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_hs_buffer.WIRE_OUT_0__9_LC_11_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8756),
            .lcout(TVP_HSYNC_buff),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24594),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.X_243__i0_LC_11_9_0 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_243__i0_LC_11_9_0 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_243__i0_LC_11_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_243__i0_LC_11_9_0  (
            .in0(_gnd_net_),
            .in1(N__8750),
            .in2(_gnd_net_),
            .in3(N__8744),
            .lcout(\receive_module.rx_counter.n10 ),
            .ltout(),
            .carryin(bfn_11_9_0_),
            .carryout(\receive_module.rx_counter.n3147 ),
            .clk(N__24599),
            .ce(),
            .sr(N__9415));
    defparam \receive_module.rx_counter.X_243__i1_LC_11_9_1 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_243__i1_LC_11_9_1 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_243__i1_LC_11_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_243__i1_LC_11_9_1  (
            .in0(_gnd_net_),
            .in1(N__8882),
            .in2(_gnd_net_),
            .in3(N__8876),
            .lcout(\receive_module.rx_counter.n9_adj_612 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3147 ),
            .carryout(\receive_module.rx_counter.n3148 ),
            .clk(N__24599),
            .ce(),
            .sr(N__9415));
    defparam \receive_module.rx_counter.X_243__i2_LC_11_9_2 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_243__i2_LC_11_9_2 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_243__i2_LC_11_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_243__i2_LC_11_9_2  (
            .in0(_gnd_net_),
            .in1(N__8873),
            .in2(_gnd_net_),
            .in3(N__8867),
            .lcout(\receive_module.rx_counter.n8_adj_611 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3148 ),
            .carryout(\receive_module.rx_counter.n3149 ),
            .clk(N__24599),
            .ce(),
            .sr(N__9415));
    defparam \receive_module.rx_counter.X_243__i3_LC_11_9_3 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_243__i3_LC_11_9_3 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_243__i3_LC_11_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_243__i3_LC_11_9_3  (
            .in0(_gnd_net_),
            .in1(N__9572),
            .in2(_gnd_net_),
            .in3(N__8864),
            .lcout(\receive_module.rx_counter.X_3 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3149 ),
            .carryout(\receive_module.rx_counter.n3150 ),
            .clk(N__24599),
            .ce(),
            .sr(N__9415));
    defparam \receive_module.rx_counter.X_243__i4_LC_11_9_4 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_243__i4_LC_11_9_4 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_243__i4_LC_11_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_243__i4_LC_11_9_4  (
            .in0(_gnd_net_),
            .in1(N__9587),
            .in2(_gnd_net_),
            .in3(N__8861),
            .lcout(\receive_module.rx_counter.X_4 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3150 ),
            .carryout(\receive_module.rx_counter.n3151 ),
            .clk(N__24599),
            .ce(),
            .sr(N__9415));
    defparam \receive_module.rx_counter.X_243__i5_LC_11_9_5 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_243__i5_LC_11_9_5 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_243__i5_LC_11_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_243__i5_LC_11_9_5  (
            .in0(_gnd_net_),
            .in1(N__9602),
            .in2(_gnd_net_),
            .in3(N__8858),
            .lcout(\receive_module.rx_counter.X_5 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3151 ),
            .carryout(\receive_module.rx_counter.n3152 ),
            .clk(N__24599),
            .ce(),
            .sr(N__9415));
    defparam \receive_module.rx_counter.X_243__i6_LC_11_9_6 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_243__i6_LC_11_9_6 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_243__i6_LC_11_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_243__i6_LC_11_9_6  (
            .in0(_gnd_net_),
            .in1(N__9557),
            .in2(_gnd_net_),
            .in3(N__8855),
            .lcout(\receive_module.rx_counter.X_6 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3152 ),
            .carryout(\receive_module.rx_counter.n3153 ),
            .clk(N__24599),
            .ce(),
            .sr(N__9415));
    defparam \receive_module.rx_counter.X_243__i7_LC_11_9_7 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_243__i7_LC_11_9_7 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_243__i7_LC_11_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_243__i7_LC_11_9_7  (
            .in0(_gnd_net_),
            .in1(N__9539),
            .in2(_gnd_net_),
            .in3(N__8852),
            .lcout(\receive_module.rx_counter.X_7 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3153 ),
            .carryout(\receive_module.rx_counter.n3154 ),
            .clk(N__24599),
            .ce(),
            .sr(N__9415));
    defparam \receive_module.rx_counter.X_243__i8_LC_11_10_0 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_243__i8_LC_11_10_0 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_243__i8_LC_11_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_243__i8_LC_11_10_0  (
            .in0(_gnd_net_),
            .in1(N__9443),
            .in2(_gnd_net_),
            .in3(N__8849),
            .lcout(\receive_module.rx_counter.X_8 ),
            .ltout(),
            .carryin(bfn_11_10_0_),
            .carryout(\receive_module.rx_counter.n3155 ),
            .clk(N__24602),
            .ce(),
            .sr(N__9416));
    defparam \receive_module.rx_counter.X_243__i9_LC_11_10_1 .C_ON=1'b0;
    defparam \receive_module.rx_counter.X_243__i9_LC_11_10_1 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_243__i9_LC_11_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_243__i9_LC_11_10_1  (
            .in0(_gnd_net_),
            .in1(N__9430),
            .in2(_gnd_net_),
            .in3(N__8846),
            .lcout(\receive_module.rx_counter.X_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24602),
            .ce(),
            .sr(N__9416));
    defparam \receive_module.i246_2_lut_rep_26_LC_11_11_0 .C_ON=1'b0;
    defparam \receive_module.i246_2_lut_rep_26_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \receive_module.i246_2_lut_rep_26_LC_11_11_0 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \receive_module.i246_2_lut_rep_26_LC_11_11_0  (
            .in0(_gnd_net_),
            .in1(N__14675),
            .in2(_gnd_net_),
            .in3(N__13089),
            .lcout(\receive_module.n3632 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.Y_DELTA_PATTERN_i57_LC_11_12_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i57_LC_11_12_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i57_LC_11_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i57_LC_11_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8906),
            .lcout(\transmit_module.Y_DELTA_PATTERN_57 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23459),
            .ce(N__15253),
            .sr(N__20335));
    defparam \transmit_module.Y_DELTA_PATTERN_i50_LC_11_12_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i50_LC_11_12_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i50_LC_11_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i50_LC_11_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8912),
            .lcout(\transmit_module.Y_DELTA_PATTERN_50 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23459),
            .ce(N__15253),
            .sr(N__20335));
    defparam \transmit_module.Y_DELTA_PATTERN_i51_LC_11_12_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i51_LC_11_12_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i51_LC_11_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i51_LC_11_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9716),
            .lcout(\transmit_module.Y_DELTA_PATTERN_51 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23459),
            .ce(N__15253),
            .sr(N__20335));
    defparam \transmit_module.Y_DELTA_PATTERN_i58_LC_11_12_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i58_LC_11_12_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i58_LC_11_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i58_LC_11_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9320),
            .lcout(\transmit_module.Y_DELTA_PATTERN_58 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23459),
            .ce(N__15253),
            .sr(N__20335));
    defparam \transmit_module.Y_DELTA_PATTERN_i56_LC_11_13_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i56_LC_11_13_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i56_LC_11_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i56_LC_11_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8900),
            .lcout(\transmit_module.Y_DELTA_PATTERN_56 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23305),
            .ce(N__15252),
            .sr(N__20294));
    defparam \transmit_module.Y_DELTA_PATTERN_i22_LC_11_14_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i22_LC_11_14_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i22_LC_11_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i22_LC_11_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8972),
            .lcout(\transmit_module.Y_DELTA_PATTERN_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23472),
            .ce(N__21033),
            .sr(N__20251));
    defparam \transmit_module.Y_DELTA_PATTERN_i21_LC_11_14_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i21_LC_11_14_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i21_LC_11_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i21_LC_11_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8894),
            .lcout(\transmit_module.Y_DELTA_PATTERN_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23472),
            .ce(N__21033),
            .sr(N__20251));
    defparam \transmit_module.Y_DELTA_PATTERN_i20_LC_11_14_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i20_LC_11_14_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i20_LC_11_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i20_LC_11_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8888),
            .lcout(\transmit_module.Y_DELTA_PATTERN_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23472),
            .ce(N__21033),
            .sr(N__20251));
    defparam \transmit_module.Y_DELTA_PATTERN_i24_LC_11_14_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i24_LC_11_14_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i24_LC_11_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i24_LC_11_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8930),
            .lcout(\transmit_module.Y_DELTA_PATTERN_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23472),
            .ce(N__21033),
            .sr(N__20251));
    defparam \transmit_module.Y_DELTA_PATTERN_i23_LC_11_14_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i23_LC_11_14_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i23_LC_11_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i23_LC_11_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8978),
            .lcout(\transmit_module.Y_DELTA_PATTERN_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23472),
            .ce(N__21033),
            .sr(N__20251));
    defparam \transmit_module.Y_DELTA_PATTERN_i27_LC_11_15_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i27_LC_11_15_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i27_LC_11_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i27_LC_11_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8966),
            .lcout(\transmit_module.Y_DELTA_PATTERN_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23484),
            .ce(N__21046),
            .sr(N__20292));
    defparam \transmit_module.Y_DELTA_PATTERN_i26_LC_11_15_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i26_LC_11_15_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i26_LC_11_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i26_LC_11_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8960),
            .lcout(\transmit_module.Y_DELTA_PATTERN_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23484),
            .ce(N__21046),
            .sr(N__20292));
    defparam \transmit_module.Y_DELTA_PATTERN_i15_LC_11_15_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i15_LC_11_15_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i15_LC_11_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i15_LC_11_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18311),
            .lcout(\transmit_module.Y_DELTA_PATTERN_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23484),
            .ce(N__21046),
            .sr(N__20292));
    defparam \transmit_module.Y_DELTA_PATTERN_i12_LC_11_15_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i12_LC_11_15_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i12_LC_11_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i12_LC_11_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8954),
            .lcout(\transmit_module.Y_DELTA_PATTERN_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23484),
            .ce(N__21046),
            .sr(N__20292));
    defparam \transmit_module.Y_DELTA_PATTERN_i13_LC_11_15_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i13_LC_11_15_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i13_LC_11_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i13_LC_11_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8942),
            .lcout(\transmit_module.Y_DELTA_PATTERN_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23484),
            .ce(N__21046),
            .sr(N__20292));
    defparam \transmit_module.Y_DELTA_PATTERN_i14_LC_11_15_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i14_LC_11_15_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i14_LC_11_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i14_LC_11_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8948),
            .lcout(\transmit_module.Y_DELTA_PATTERN_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23484),
            .ce(N__21046),
            .sr(N__20292));
    defparam \transmit_module.Y_DELTA_PATTERN_i25_LC_11_15_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i25_LC_11_15_7 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i25_LC_11_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i25_LC_11_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8936),
            .lcout(\transmit_module.Y_DELTA_PATTERN_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23484),
            .ce(N__21046),
            .sr(N__20292));
    defparam \transmit_module.Y_DELTA_PATTERN_i8_LC_11_16_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i8_LC_11_16_2 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i8_LC_11_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i8_LC_11_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9029),
            .lcout(\transmit_module.Y_DELTA_PATTERN_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23377),
            .ce(N__21009),
            .sr(N__20164));
    defparam \transmit_module.Y_DELTA_PATTERN_i99_LC_11_16_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i99_LC_11_16_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i99_LC_11_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i99_LC_11_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20657),
            .lcout(\transmit_module.Y_DELTA_PATTERN_99 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23377),
            .ce(N__21009),
            .sr(N__20164));
    defparam \transmit_module.Y_DELTA_PATTERN_i10_LC_11_16_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i10_LC_11_16_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i10_LC_11_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i10_LC_11_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9017),
            .lcout(\transmit_module.Y_DELTA_PATTERN_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23377),
            .ce(N__21009),
            .sr(N__20164));
    defparam \transmit_module.Y_DELTA_PATTERN_i9_LC_11_16_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i9_LC_11_16_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i9_LC_11_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i9_LC_11_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9035),
            .lcout(\transmit_module.Y_DELTA_PATTERN_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23377),
            .ce(N__21009),
            .sr(N__20164));
    defparam \transmit_module.Y_DELTA_PATTERN_i11_LC_11_16_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i11_LC_11_16_7 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i11_LC_11_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i11_LC_11_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9023),
            .lcout(\transmit_module.Y_DELTA_PATTERN_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23377),
            .ce(N__21009),
            .sr(N__20164));
    defparam \transmit_module.Y_DELTA_PATTERN_i40_LC_11_17_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i40_LC_11_17_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i40_LC_11_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i40_LC_11_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8990),
            .lcout(\transmit_module.Y_DELTA_PATTERN_40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23434),
            .ce(N__15212),
            .sr(N__20392));
    defparam \transmit_module.Y_DELTA_PATTERN_i38_LC_11_17_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i38_LC_11_17_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i38_LC_11_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i38_LC_11_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8996),
            .lcout(\transmit_module.Y_DELTA_PATTERN_38 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23434),
            .ce(N__15212),
            .sr(N__20392));
    defparam \transmit_module.Y_DELTA_PATTERN_i39_LC_11_17_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i39_LC_11_17_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i39_LC_11_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i39_LC_11_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9002),
            .lcout(\transmit_module.Y_DELTA_PATTERN_39 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23434),
            .ce(N__15212),
            .sr(N__20392));
    defparam \transmit_module.Y_DELTA_PATTERN_i41_LC_11_17_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i41_LC_11_17_7 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i41_LC_11_17_7 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i41_LC_11_17_7  (
            .in0(_gnd_net_),
            .in1(N__8984),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.Y_DELTA_PATTERN_41 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23434),
            .ce(N__15212),
            .sr(N__20392));
    defparam \transmit_module.Y_DELTA_PATTERN_i42_LC_11_18_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i42_LC_11_18_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i42_LC_11_18_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i42_LC_11_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9326),
            .lcout(\transmit_module.Y_DELTA_PATTERN_42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23371),
            .ce(N__15199),
            .sr(N__20339));
    defparam \transmit_module.Y_DELTA_PATTERN_i45_LC_11_18_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i45_LC_11_18_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i45_LC_11_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i45_LC_11_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9290),
            .lcout(\transmit_module.Y_DELTA_PATTERN_45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23371),
            .ce(N__15199),
            .sr(N__20339));
    defparam \transmit_module.Y_DELTA_PATTERN_i43_LC_11_18_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i43_LC_11_18_2 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i43_LC_11_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i43_LC_11_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9305),
            .lcout(\transmit_module.Y_DELTA_PATTERN_43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23371),
            .ce(N__15199),
            .sr(N__20339));
    defparam \transmit_module.Y_DELTA_PATTERN_i59_LC_11_18_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i59_LC_11_18_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i59_LC_11_18_5 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i59_LC_11_18_5  (
            .in0(_gnd_net_),
            .in1(N__9278),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.Y_DELTA_PATTERN_59 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23371),
            .ce(N__15199),
            .sr(N__20339));
    defparam \transmit_module.Y_DELTA_PATTERN_i44_LC_11_18_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i44_LC_11_18_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i44_LC_11_18_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i44_LC_11_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9311),
            .lcout(\transmit_module.Y_DELTA_PATTERN_44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23371),
            .ce(N__15199),
            .sr(N__20339));
    defparam \transmit_module.Y_DELTA_PATTERN_i46_LC_11_18_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i46_LC_11_18_7 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i46_LC_11_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i46_LC_11_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9299),
            .lcout(\transmit_module.Y_DELTA_PATTERN_46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23371),
            .ce(N__15199),
            .sr(N__20339));
    defparam \transmit_module.Y_DELTA_PATTERN_i60_LC_11_19_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i60_LC_11_19_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i60_LC_11_19_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i60_LC_11_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9284),
            .lcout(\transmit_module.Y_DELTA_PATTERN_60 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23154),
            .ce(N__15219),
            .sr(N__20296));
    defparam \transmit_module.Y_DELTA_PATTERN_i76_LC_11_19_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i76_LC_11_19_2 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i76_LC_11_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i76_LC_11_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9272),
            .lcout(\transmit_module.Y_DELTA_PATTERN_76 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23154),
            .ce(N__15219),
            .sr(N__20296));
    defparam \transmit_module.i1613_4_lut_LC_11_31_3 .C_ON=1'b0;
    defparam \transmit_module.i1613_4_lut_LC_11_31_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1613_4_lut_LC_11_31_3 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \transmit_module.i1613_4_lut_LC_11_31_3  (
            .in0(N__20877),
            .in1(N__20557),
            .in2(N__20408),
            .in3(N__18245),
            .lcout(n24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.BUFFER_0__i3_LC_12_3_1 .C_ON=1'b0;
    defparam \tvp_video_buffer.BUFFER_0__i3_LC_12_3_1 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.BUFFER_0__i3_LC_12_3_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.BUFFER_0__i3_LC_12_3_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9053),
            .lcout(\tvp_video_buffer.BUFFER_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24568),
            .ce(),
            .sr(_gnd_net_));
    defparam \TVP_VSYNC_buff_I_0.BUFFER_0__i1_LC_12_6_6 .C_ON=1'b0;
    defparam \TVP_VSYNC_buff_I_0.BUFFER_0__i1_LC_12_6_6 .SEQ_MODE=4'b1000;
    defparam \TVP_VSYNC_buff_I_0.BUFFER_0__i1_LC_12_6_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \TVP_VSYNC_buff_I_0.BUFFER_0__i1_LC_12_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9469),
            .lcout(\TVP_VSYNC_buff_I_0.BUFFER_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVTVP_VSYNC_buff_I_0.BUFFER_0__i1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i130_2_lut_rep_17_LC_12_7_3 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i130_2_lut_rep_17_LC_12_7_3 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i130_2_lut_rep_17_LC_12_7_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \receive_module.rx_counter.i130_2_lut_rep_17_LC_12_7_3  (
            .in0(N__13088),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12521),
            .lcout(\receive_module.rx_counter.n3623 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \TVP_VSYNC_buff_I_0.BUFFER_0__i2_LC_12_7_4 .C_ON=1'b0;
    defparam \TVP_VSYNC_buff_I_0.BUFFER_0__i2_LC_12_7_4 .SEQ_MODE=4'b1000;
    defparam \TVP_VSYNC_buff_I_0.BUFFER_0__i2_LC_12_7_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \TVP_VSYNC_buff_I_0.BUFFER_0__i2_LC_12_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9449),
            .lcout(\TVP_VSYNC_buff_I_0.BUFFER_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVTVP_VSYNC_buff_I_0.BUFFER_0__i2C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.old_HS_51_LC_12_8_1 .C_ON=1'b0;
    defparam \receive_module.rx_counter.old_HS_51_LC_12_8_1 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.old_HS_51_LC_12_8_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \receive_module.rx_counter.old_HS_51_LC_12_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9508),
            .lcout(\receive_module.rx_counter.old_HS ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24591),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i59_4_lut_LC_12_9_2 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i59_4_lut_LC_12_9_2 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i59_4_lut_LC_12_9_2 .LUT_INIT=16'b1110000011100101;
    LogicCell40 \receive_module.rx_counter.i59_4_lut_LC_12_9_2  (
            .in0(N__9442),
            .in1(N__9653),
            .in2(N__9431),
            .in3(N__9524),
            .lcout(\receive_module.rx_counter.n55_adj_606 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i5_1_lut_rep_24_LC_12_9_3 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i5_1_lut_rep_24_LC_12_9_3 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i5_1_lut_rep_24_LC_12_9_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \receive_module.rx_counter.i5_1_lut_rep_24_LC_12_9_3  (
            .in0(N__9504),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\receive_module.rx_counter.n3630 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \TVP_VSYNC_buff_I_0.WIRE_OUT_0__9_LC_12_9_6 .C_ON=1'b0;
    defparam \TVP_VSYNC_buff_I_0.WIRE_OUT_0__9_LC_12_9_6 .SEQ_MODE=4'b1000;
    defparam \TVP_VSYNC_buff_I_0.WIRE_OUT_0__9_LC_12_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \TVP_VSYNC_buff_I_0.WIRE_OUT_0__9_LC_12_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9392),
            .lcout(TVP_VSYNC_buff),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVTVP_VSYNC_buff_I_0.WIRE_OUT_0__9C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_14_LC_12_9_7 .C_ON=1'b0;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_14_LC_12_9_7 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_14_LC_12_9_7 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \line_buffer.i1_2_lut_3_lut_4_lut_adj_14_LC_12_9_7  (
            .in0(N__14794),
            .in1(N__14643),
            .in2(N__14560),
            .in3(N__14455),
            .lcout(\line_buffer.n467 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i1_2_lut_adj_18_LC_12_10_0 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i1_2_lut_adj_18_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i1_2_lut_adj_18_LC_12_10_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \receive_module.rx_counter.i1_2_lut_adj_18_LC_12_10_0  (
            .in0(_gnd_net_),
            .in1(N__9570),
            .in2(_gnd_net_),
            .in3(N__9585),
            .lcout(),
            .ltout(\receive_module.rx_counter.n4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i2_4_lut_adj_19_LC_12_10_1 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i2_4_lut_adj_19_LC_12_10_1 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i2_4_lut_adj_19_LC_12_10_1 .LUT_INIT=16'b1100100000000000;
    LogicCell40 \receive_module.rx_counter.i2_4_lut_adj_19_LC_12_10_1  (
            .in0(N__9601),
            .in1(N__9555),
            .in2(N__9656),
            .in3(N__9537),
            .lcout(\receive_module.rx_counter.n3400 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_15_LC_12_10_2 .C_ON=1'b0;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_15_LC_12_10_2 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_15_LC_12_10_2 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \line_buffer.i1_2_lut_3_lut_4_lut_adj_15_LC_12_10_2  (
            .in0(N__14649),
            .in1(N__14795),
            .in2(N__14561),
            .in3(N__14467),
            .lcout(\line_buffer.n565 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i2_2_lut_adj_20_LC_12_10_4 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i2_2_lut_adj_20_LC_12_10_4 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i2_2_lut_adj_20_LC_12_10_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \receive_module.rx_counter.i2_2_lut_adj_20_LC_12_10_4  (
            .in0(_gnd_net_),
            .in1(N__9600),
            .in2(_gnd_net_),
            .in3(N__9586),
            .lcout(),
            .ltout(\receive_module.rx_counter.n6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i2042_4_lut_LC_12_10_5 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i2042_4_lut_LC_12_10_5 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i2042_4_lut_LC_12_10_5 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \receive_module.rx_counter.i2042_4_lut_LC_12_10_5  (
            .in0(N__9571),
            .in1(N__9556),
            .in2(N__9542),
            .in3(N__9538),
            .lcout(\receive_module.rx_counter.n3385 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.O_VS_I_0_1_lut_rep_25_LC_12_10_6 .C_ON=1'b0;
    defparam \receive_module.rx_counter.O_VS_I_0_1_lut_rep_25_LC_12_10_6 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.O_VS_I_0_1_lut_rep_25_LC_12_10_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \receive_module.rx_counter.O_VS_I_0_1_lut_rep_25_LC_12_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13067),
            .lcout(\receive_module.n3631 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i249_3_lut_3_lut_3_lut_LC_12_10_7 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i249_3_lut_3_lut_3_lut_LC_12_10_7 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i249_3_lut_3_lut_3_lut_LC_12_10_7 .LUT_INIT=16'b0101010111011101;
    LogicCell40 \receive_module.rx_counter.i249_3_lut_3_lut_3_lut_LC_12_10_7  (
            .in0(N__13068),
            .in1(N__9518),
            .in2(_gnd_net_),
            .in3(N__9509),
            .lcout(\receive_module.rx_counter.n2063 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_2_lut_LC_12_11_0 .C_ON=1'b1;
    defparam \receive_module.add_12_2_lut_LC_12_11_0 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_2_lut_LC_12_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_2_lut_LC_12_11_0  (
            .in0(_gnd_net_),
            .in1(N__10128),
            .in2(_gnd_net_),
            .in3(N__9488),
            .lcout(\receive_module.n136 ),
            .ltout(),
            .carryin(bfn_12_11_0_),
            .carryout(\receive_module.n3091 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_3_lut_LC_12_11_1 .C_ON=1'b1;
    defparam \receive_module.add_12_3_lut_LC_12_11_1 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_3_lut_LC_12_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_3_lut_LC_12_11_1  (
            .in0(_gnd_net_),
            .in1(N__9870),
            .in2(_gnd_net_),
            .in3(N__9485),
            .lcout(\receive_module.n135 ),
            .ltout(),
            .carryin(\receive_module.n3091 ),
            .carryout(\receive_module.n3092 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_4_lut_LC_12_11_2 .C_ON=1'b1;
    defparam \receive_module.add_12_4_lut_LC_12_11_2 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_4_lut_LC_12_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_4_lut_LC_12_11_2  (
            .in0(_gnd_net_),
            .in1(N__12831),
            .in2(_gnd_net_),
            .in3(N__9482),
            .lcout(\receive_module.n134 ),
            .ltout(),
            .carryin(\receive_module.n3092 ),
            .carryout(\receive_module.n3093 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_5_lut_LC_12_11_3 .C_ON=1'b1;
    defparam \receive_module.add_12_5_lut_LC_12_11_3 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_5_lut_LC_12_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_5_lut_LC_12_11_3  (
            .in0(_gnd_net_),
            .in1(N__12045),
            .in2(_gnd_net_),
            .in3(N__9683),
            .lcout(\receive_module.n133 ),
            .ltout(),
            .carryin(\receive_module.n3093 ),
            .carryout(\receive_module.n3094 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_6_lut_LC_12_11_4 .C_ON=1'b1;
    defparam \receive_module.add_12_6_lut_LC_12_11_4 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_6_lut_LC_12_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_6_lut_LC_12_11_4  (
            .in0(_gnd_net_),
            .in1(N__11787),
            .in2(_gnd_net_),
            .in3(N__9680),
            .lcout(\receive_module.n132 ),
            .ltout(),
            .carryin(\receive_module.n3094 ),
            .carryout(\receive_module.n3095 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_7_lut_LC_12_11_5 .C_ON=1'b1;
    defparam \receive_module.add_12_7_lut_LC_12_11_5 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_7_lut_LC_12_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_7_lut_LC_12_11_5  (
            .in0(_gnd_net_),
            .in1(N__11403),
            .in2(_gnd_net_),
            .in3(N__9677),
            .lcout(\receive_module.n131 ),
            .ltout(),
            .carryin(\receive_module.n3095 ),
            .carryout(\receive_module.n3096 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_8_lut_LC_12_11_6 .C_ON=1'b1;
    defparam \receive_module.add_12_8_lut_LC_12_11_6 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_8_lut_LC_12_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_8_lut_LC_12_11_6  (
            .in0(_gnd_net_),
            .in1(N__11145),
            .in2(_gnd_net_),
            .in3(N__9674),
            .lcout(\receive_module.n130 ),
            .ltout(),
            .carryin(\receive_module.n3096 ),
            .carryout(\receive_module.n3097 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_9_lut_LC_12_11_7 .C_ON=1'b1;
    defparam \receive_module.add_12_9_lut_LC_12_11_7 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_9_lut_LC_12_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_9_lut_LC_12_11_7  (
            .in0(_gnd_net_),
            .in1(N__10872),
            .in2(_gnd_net_),
            .in3(N__9671),
            .lcout(\receive_module.n129 ),
            .ltout(),
            .carryin(\receive_module.n3097 ),
            .carryout(\receive_module.n3098 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_10_lut_LC_12_12_0 .C_ON=1'b1;
    defparam \receive_module.add_12_10_lut_LC_12_12_0 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_10_lut_LC_12_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_10_lut_LC_12_12_0  (
            .in0(_gnd_net_),
            .in1(N__10632),
            .in2(_gnd_net_),
            .in3(N__9668),
            .lcout(\receive_module.n128 ),
            .ltout(),
            .carryin(bfn_12_12_0_),
            .carryout(\receive_module.n3099 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_11_lut_LC_12_12_1 .C_ON=1'b1;
    defparam \receive_module.add_12_11_lut_LC_12_12_1 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_11_lut_LC_12_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_11_lut_LC_12_12_1  (
            .in0(_gnd_net_),
            .in1(N__10371),
            .in2(_gnd_net_),
            .in3(N__9665),
            .lcout(\receive_module.n127 ),
            .ltout(),
            .carryin(\receive_module.n3099 ),
            .carryout(\receive_module.n3100 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_12_lut_LC_12_12_2 .C_ON=1'b1;
    defparam \receive_module.add_12_12_lut_LC_12_12_2 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_12_lut_LC_12_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_12_lut_LC_12_12_2  (
            .in0(_gnd_net_),
            .in1(N__12294),
            .in2(_gnd_net_),
            .in3(N__9662),
            .lcout(\receive_module.n126 ),
            .ltout(),
            .carryin(\receive_module.n3100 ),
            .carryout(\receive_module.n3101 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.BRAM_ADDR__i11_LC_12_12_3 .C_ON=1'b1;
    defparam \receive_module.BRAM_ADDR__i11_LC_12_12_3 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i11_LC_12_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.BRAM_ADDR__i11_LC_12_12_3  (
            .in0(_gnd_net_),
            .in1(N__14430),
            .in2(_gnd_net_),
            .in3(N__9659),
            .lcout(RX_ADDR_11),
            .ltout(),
            .carryin(\receive_module.n3101 ),
            .carryout(\receive_module.n3102 ),
            .clk(N__24605),
            .ce(N__9734),
            .sr(N__12761));
    defparam \receive_module.BRAM_ADDR__i12_LC_12_12_4 .C_ON=1'b1;
    defparam \receive_module.BRAM_ADDR__i12_LC_12_12_4 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i12_LC_12_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.BRAM_ADDR__i12_LC_12_12_4  (
            .in0(_gnd_net_),
            .in1(N__14778),
            .in2(_gnd_net_),
            .in3(N__9740),
            .lcout(RX_ADDR_12),
            .ltout(),
            .carryin(\receive_module.n3102 ),
            .carryout(\receive_module.n3103 ),
            .clk(N__24605),
            .ce(N__9734),
            .sr(N__12761));
    defparam \receive_module.BRAM_ADDR__i13_LC_12_12_5 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i13_LC_12_12_5 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i13_LC_12_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.BRAM_ADDR__i13_LC_12_12_5  (
            .in0(_gnd_net_),
            .in1(N__14532),
            .in2(_gnd_net_),
            .in3(N__9737),
            .lcout(RX_ADDR_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24605),
            .ce(N__9734),
            .sr(N__12761));
    defparam \transmit_module.Y_DELTA_PATTERN_i53_LC_12_13_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i53_LC_12_13_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i53_LC_12_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i53_LC_12_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9698),
            .lcout(\transmit_module.Y_DELTA_PATTERN_53 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23486),
            .ce(N__15249),
            .sr(N__20415));
    defparam \transmit_module.Y_DELTA_PATTERN_i52_LC_12_13_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i52_LC_12_13_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i52_LC_12_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i52_LC_12_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9722),
            .lcout(\transmit_module.Y_DELTA_PATTERN_52 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23486),
            .ce(N__15249),
            .sr(N__20415));
    defparam \transmit_module.Y_DELTA_PATTERN_i55_LC_12_13_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i55_LC_12_13_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i55_LC_12_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i55_LC_12_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9710),
            .lcout(\transmit_module.Y_DELTA_PATTERN_55 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23486),
            .ce(N__15249),
            .sr(N__20415));
    defparam \transmit_module.Y_DELTA_PATTERN_i54_LC_12_13_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i54_LC_12_13_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i54_LC_12_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i54_LC_12_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9704),
            .lcout(\transmit_module.Y_DELTA_PATTERN_54 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23486),
            .ce(N__15249),
            .sr(N__20415));
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_23_LC_12_14_4 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_23_LC_12_14_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_23_LC_12_14_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \transmit_module.video_signal_controller.i1_2_lut_rep_23_LC_12_14_4  (
            .in0(_gnd_net_),
            .in1(N__15299),
            .in2(_gnd_net_),
            .in3(N__13632),
            .lcout(),
            .ltout(\transmit_module.video_signal_controller.n3629_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_4_lut_adj_24_LC_12_14_5 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_4_lut_adj_24_LC_12_14_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_4_lut_adj_24_LC_12_14_5 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \transmit_module.video_signal_controller.i1_4_lut_adj_24_LC_12_14_5  (
            .in0(N__9689),
            .in1(N__13656),
            .in2(N__9692),
            .in3(N__13340),
            .lcout(\transmit_module.video_signal_controller.n4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1653_2_lut_LC_12_14_7 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1653_2_lut_LC_12_14_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1653_2_lut_LC_12_14_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \transmit_module.video_signal_controller.i1653_2_lut_LC_12_14_7  (
            .in0(_gnd_net_),
            .in1(N__13291),
            .in2(_gnd_net_),
            .in3(N__13312),
            .lcout(\transmit_module.video_signal_controller.n2901 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.VGA_X_i0_LC_12_15_0 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i0_LC_12_15_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i0_LC_12_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i0_LC_12_15_0  (
            .in0(_gnd_net_),
            .in1(N__13292),
            .in2(_gnd_net_),
            .in3(N__9767),
            .lcout(\transmit_module.video_signal_controller.VGA_X_0 ),
            .ltout(),
            .carryin(bfn_12_15_0_),
            .carryout(\transmit_module.video_signal_controller.n3125 ),
            .clk(N__23132),
            .ce(),
            .sr(N__14248));
    defparam \transmit_module.video_signal_controller.VGA_X_i1_LC_12_15_1 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i1_LC_12_15_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i1_LC_12_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i1_LC_12_15_1  (
            .in0(_gnd_net_),
            .in1(N__13313),
            .in2(_gnd_net_),
            .in3(N__9764),
            .lcout(\transmit_module.video_signal_controller.VGA_X_1 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3125 ),
            .carryout(\transmit_module.video_signal_controller.n3126 ),
            .clk(N__23132),
            .ce(),
            .sr(N__14248));
    defparam \transmit_module.video_signal_controller.VGA_X_i2_LC_12_15_2 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i2_LC_12_15_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i2_LC_12_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i2_LC_12_15_2  (
            .in0(_gnd_net_),
            .in1(N__13341),
            .in2(_gnd_net_),
            .in3(N__9761),
            .lcout(\transmit_module.video_signal_controller.VGA_X_2 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3126 ),
            .carryout(\transmit_module.video_signal_controller.n3127 ),
            .clk(N__23132),
            .ce(),
            .sr(N__14248));
    defparam \transmit_module.video_signal_controller.VGA_X_i3_LC_12_15_3 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i3_LC_12_15_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i3_LC_12_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i3_LC_12_15_3  (
            .in0(_gnd_net_),
            .in1(N__13657),
            .in2(_gnd_net_),
            .in3(N__9758),
            .lcout(\transmit_module.video_signal_controller.VGA_X_3 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3127 ),
            .carryout(\transmit_module.video_signal_controller.n3128 ),
            .clk(N__23132),
            .ce(),
            .sr(N__14248));
    defparam \transmit_module.video_signal_controller.VGA_X_i4_LC_12_15_4 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i4_LC_12_15_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i4_LC_12_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i4_LC_12_15_4  (
            .in0(_gnd_net_),
            .in1(N__13514),
            .in2(_gnd_net_),
            .in3(N__9755),
            .lcout(\transmit_module.video_signal_controller.VGA_X_4 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3128 ),
            .carryout(\transmit_module.video_signal_controller.n3129 ),
            .clk(N__23132),
            .ce(),
            .sr(N__14248));
    defparam \transmit_module.video_signal_controller.VGA_X_i5_LC_12_15_5 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i5_LC_12_15_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i5_LC_12_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i5_LC_12_15_5  (
            .in0(_gnd_net_),
            .in1(N__13634),
            .in2(_gnd_net_),
            .in3(N__9752),
            .lcout(\transmit_module.video_signal_controller.VGA_X_5 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3129 ),
            .carryout(\transmit_module.video_signal_controller.n3130 ),
            .clk(N__23132),
            .ce(),
            .sr(N__14248));
    defparam \transmit_module.video_signal_controller.VGA_X_i6_LC_12_15_6 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i6_LC_12_15_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i6_LC_12_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i6_LC_12_15_6  (
            .in0(_gnd_net_),
            .in1(N__15300),
            .in2(_gnd_net_),
            .in3(N__9749),
            .lcout(\transmit_module.video_signal_controller.VGA_X_6 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3130 ),
            .carryout(\transmit_module.video_signal_controller.n3131 ),
            .clk(N__23132),
            .ce(),
            .sr(N__14248));
    defparam \transmit_module.video_signal_controller.VGA_X_i7_LC_12_15_7 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i7_LC_12_15_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i7_LC_12_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i7_LC_12_15_7  (
            .in0(_gnd_net_),
            .in1(N__13539),
            .in2(_gnd_net_),
            .in3(N__9746),
            .lcout(\transmit_module.video_signal_controller.VGA_X_7 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3131 ),
            .carryout(\transmit_module.video_signal_controller.n3132 ),
            .clk(N__23132),
            .ce(),
            .sr(N__14248));
    defparam \transmit_module.video_signal_controller.VGA_X_i8_LC_12_16_0 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i8_LC_12_16_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i8_LC_12_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i8_LC_12_16_0  (
            .in0(_gnd_net_),
            .in1(N__15350),
            .in2(_gnd_net_),
            .in3(N__9743),
            .lcout(\transmit_module.video_signal_controller.VGA_X_8 ),
            .ltout(),
            .carryin(bfn_12_16_0_),
            .carryout(\transmit_module.video_signal_controller.n3133 ),
            .clk(N__23404),
            .ce(),
            .sr(N__14252));
    defparam \transmit_module.video_signal_controller.VGA_X_i9_LC_12_16_1 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i9_LC_12_16_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i9_LC_12_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i9_LC_12_16_1  (
            .in0(_gnd_net_),
            .in1(N__13602),
            .in2(_gnd_net_),
            .in3(N__9800),
            .lcout(\transmit_module.video_signal_controller.VGA_X_9 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3133 ),
            .carryout(\transmit_module.video_signal_controller.n3134 ),
            .clk(N__23404),
            .ce(),
            .sr(N__14252));
    defparam \transmit_module.video_signal_controller.VGA_X_i10_LC_12_16_2 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i10_LC_12_16_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i10_LC_12_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i10_LC_12_16_2  (
            .in0(_gnd_net_),
            .in1(N__13573),
            .in2(_gnd_net_),
            .in3(N__9797),
            .lcout(\transmit_module.video_signal_controller.VGA_X_10 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3134 ),
            .carryout(\transmit_module.video_signal_controller.n3135 ),
            .clk(N__23404),
            .ce(),
            .sr(N__14252));
    defparam \transmit_module.video_signal_controller.VGA_X_i11_LC_12_16_3 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.VGA_X_i11_LC_12_16_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i11_LC_12_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i11_LC_12_16_3  (
            .in0(_gnd_net_),
            .in1(N__16716),
            .in2(_gnd_net_),
            .in3(N__9794),
            .lcout(\transmit_module.video_signal_controller.VGA_X_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23404),
            .ce(),
            .sr(N__14252));
    defparam \transmit_module.i123_2_lut_4_lut_rep_29_LC_12_17_7 .C_ON=1'b0;
    defparam \transmit_module.i123_2_lut_4_lut_rep_29_LC_12_17_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i123_2_lut_4_lut_rep_29_LC_12_17_7 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \transmit_module.i123_2_lut_4_lut_rep_29_LC_12_17_7  (
            .in0(N__16403),
            .in1(N__16427),
            .in2(N__20326),
            .in3(N__16369),
            .lcout(\transmit_module.n3635 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.Y_DELTA_PATTERN_i1_LC_12_18_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i1_LC_12_18_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i1_LC_12_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i1_LC_12_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9791),
            .lcout(\transmit_module.Y_DELTA_PATTERN_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23229),
            .ce(N__20990),
            .sr(N__20260));
    defparam \transmit_module.Y_DELTA_PATTERN_i2_LC_12_18_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i2_LC_12_18_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i2_LC_12_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i2_LC_12_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9785),
            .lcout(\transmit_module.Y_DELTA_PATTERN_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23229),
            .ce(N__20990),
            .sr(N__20260));
    defparam \transmit_module.Y_DELTA_PATTERN_i3_LC_12_18_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i3_LC_12_18_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i3_LC_12_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i3_LC_12_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9773),
            .lcout(\transmit_module.Y_DELTA_PATTERN_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23229),
            .ce(N__20990),
            .sr(N__20260));
    defparam \transmit_module.Y_DELTA_PATTERN_i5_LC_12_18_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i5_LC_12_18_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i5_LC_12_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i5_LC_12_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11615),
            .lcout(\transmit_module.Y_DELTA_PATTERN_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23229),
            .ce(N__20990),
            .sr(N__20260));
    defparam \transmit_module.Y_DELTA_PATTERN_i4_LC_12_18_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i4_LC_12_18_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i4_LC_12_18_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i4_LC_12_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9779),
            .lcout(\transmit_module.Y_DELTA_PATTERN_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23229),
            .ce(N__20990),
            .sr(N__20260));
    defparam \transmit_module.Y_DELTA_PATTERN_i6_LC_12_18_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i6_LC_12_18_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i6_LC_12_18_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i6_LC_12_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11627),
            .lcout(\transmit_module.Y_DELTA_PATTERN_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23229),
            .ce(N__20990),
            .sr(N__20260));
    defparam \receive_module.BRAM_ADDR__i5_LC_12_19_0 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i5_LC_12_19_0 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i5_LC_12_19_0 .LUT_INIT=16'b1010110010101010;
    LogicCell40 \receive_module.BRAM_ADDR__i5_LC_12_19_0  (
            .in0(N__11609),
            .in1(N__11378),
            .in2(N__14732),
            .in3(N__13118),
            .lcout(RX_ADDR_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24614),
            .ce(),
            .sr(N__12786));
    defparam \receive_module.BRAM_ADDR__i6_LC_12_19_1 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i6_LC_12_19_1 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i6_LC_12_19_1 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \receive_module.BRAM_ADDR__i6_LC_12_19_1  (
            .in0(N__13119),
            .in1(N__14718),
            .in2(N__11129),
            .in3(N__11351),
            .lcout(RX_ADDR_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24614),
            .ce(),
            .sr(N__12786));
    defparam \receive_module.BRAM_ADDR__i7_LC_12_19_2 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i7_LC_12_19_2 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i7_LC_12_19_2 .LUT_INIT=16'b1100101011001100;
    LogicCell40 \receive_module.BRAM_ADDR__i7_LC_12_19_2  (
            .in0(N__10862),
            .in1(N__11090),
            .in2(N__14733),
            .in3(N__13120),
            .lcout(RX_ADDR_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24614),
            .ce(),
            .sr(N__12786));
    defparam \receive_module.BRAM_ADDR__i8_LC_12_19_3 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i8_LC_12_19_3 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i8_LC_12_19_3 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \receive_module.BRAM_ADDR__i8_LC_12_19_3  (
            .in0(N__13121),
            .in1(N__14722),
            .in2(N__10625),
            .in3(N__10835),
            .lcout(RX_ADDR_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24614),
            .ce(),
            .sr(N__12786));
    defparam \receive_module.BRAM_ADDR__i9_LC_12_19_4 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i9_LC_12_19_4 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i9_LC_12_19_4 .LUT_INIT=16'b1100101011001100;
    LogicCell40 \receive_module.BRAM_ADDR__i9_LC_12_19_4  (
            .in0(N__10356),
            .in1(N__10586),
            .in2(N__14734),
            .in3(N__13122),
            .lcout(RX_ADDR_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24614),
            .ce(),
            .sr(N__12786));
    defparam \receive_module.BRAM_ADDR__i0_LC_12_19_6 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i0_LC_12_19_6 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i0_LC_12_19_6 .LUT_INIT=16'b1010110010101010;
    LogicCell40 \receive_module.BRAM_ADDR__i0_LC_12_19_6  (
            .in0(N__10334),
            .in1(N__10106),
            .in2(N__14731),
            .in3(N__13116),
            .lcout(RX_ADDR_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24614),
            .ce(),
            .sr(N__12786));
    defparam \receive_module.BRAM_ADDR__i1_LC_12_19_7 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i1_LC_12_19_7 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i1_LC_12_19_7 .LUT_INIT=16'b1111001011010000;
    LogicCell40 \receive_module.BRAM_ADDR__i1_LC_12_19_7  (
            .in0(N__13117),
            .in1(N__14714),
            .in2(N__10079),
            .in3(N__9851),
            .lcout(RX_ADDR_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24614),
            .ce(),
            .sr(N__12786));
    defparam \line_buffer.i2158_3_lut_LC_12_21_3 .C_ON=1'b0;
    defparam \line_buffer.i2158_3_lut_LC_12_21_3 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2158_3_lut_LC_12_21_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \line_buffer.i2158_3_lut_LC_12_21_3  (
            .in0(N__24358),
            .in1(N__9824),
            .in2(_gnd_net_),
            .in3(N__9812),
            .lcout(\line_buffer.n3501 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.BRAM_ADDR__i10_LC_12_23_0 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i10_LC_12_23_0 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i10_LC_12_23_0 .LUT_INIT=16'b1100101011001100;
    LogicCell40 \receive_module.BRAM_ADDR__i10_LC_12_23_0  (
            .in0(N__12269),
            .in1(N__12494),
            .in2(N__14738),
            .in3(N__13129),
            .lcout(RX_ADDR_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24619),
            .ce(),
            .sr(N__12795));
    defparam \receive_module.BRAM_ADDR__i3_LC_12_29_6 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i3_LC_12_29_6 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i3_LC_12_29_6 .LUT_INIT=16'b1010110010101010;
    LogicCell40 \receive_module.BRAM_ADDR__i3_LC_12_29_6  (
            .in0(N__12239),
            .in1(N__12017),
            .in2(N__14729),
            .in3(N__13141),
            .lcout(RX_ADDR_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24626),
            .ce(),
            .sr(N__12808));
    defparam \receive_module.BRAM_ADDR__i4_LC_12_30_6 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i4_LC_12_30_6 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i4_LC_12_30_6 .LUT_INIT=16'b1010110010101010;
    LogicCell40 \receive_module.BRAM_ADDR__i4_LC_12_30_6  (
            .in0(N__11990),
            .in1(N__11759),
            .in2(N__14730),
            .in3(N__13142),
            .lcout(RX_ADDR_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24628),
            .ce(),
            .sr(N__12809));
    defparam \tvp_video_buffer.WIRE_OUT_i0_LC_13_4_4 .C_ON=1'b0;
    defparam \tvp_video_buffer.WIRE_OUT_i0_LC_13_4_4 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.WIRE_OUT_i0_LC_13_4_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.WIRE_OUT_i0_LC_13_4_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11732),
            .lcout(RX_DATA_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24569),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.FRAME_COUNTER_244__i0_LC_13_6_0 .C_ON=1'b1;
    defparam \receive_module.rx_counter.FRAME_COUNTER_244__i0_LC_13_6_0 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.FRAME_COUNTER_244__i0_LC_13_6_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.FRAME_COUNTER_244__i0_LC_13_6_0  (
            .in0(_gnd_net_),
            .in1(N__12563),
            .in2(_gnd_net_),
            .in3(N__11639),
            .lcout(\receive_module.rx_counter.FRAME_COUNTER_0 ),
            .ltout(),
            .carryin(bfn_13_6_0_),
            .carryout(\receive_module.rx_counter.n3156 ),
            .clk(N__24576),
            .ce(N__12623),
            .sr(N__12506));
    defparam \receive_module.rx_counter.FRAME_COUNTER_244__i1_LC_13_6_1 .C_ON=1'b1;
    defparam \receive_module.rx_counter.FRAME_COUNTER_244__i1_LC_13_6_1 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.FRAME_COUNTER_244__i1_LC_13_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.FRAME_COUNTER_244__i1_LC_13_6_1  (
            .in0(_gnd_net_),
            .in1(N__12575),
            .in2(_gnd_net_),
            .in3(N__11636),
            .lcout(\receive_module.rx_counter.FRAME_COUNTER_1 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3156 ),
            .carryout(\receive_module.rx_counter.n3157 ),
            .clk(N__24576),
            .ce(N__12623),
            .sr(N__12506));
    defparam \receive_module.rx_counter.FRAME_COUNTER_244__i2_LC_13_6_2 .C_ON=1'b1;
    defparam \receive_module.rx_counter.FRAME_COUNTER_244__i2_LC_13_6_2 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.FRAME_COUNTER_244__i2_LC_13_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.FRAME_COUNTER_244__i2_LC_13_6_2  (
            .in0(_gnd_net_),
            .in1(N__12599),
            .in2(_gnd_net_),
            .in3(N__11633),
            .lcout(\receive_module.rx_counter.FRAME_COUNTER_2 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3157 ),
            .carryout(\receive_module.rx_counter.n3158 ),
            .clk(N__24576),
            .ce(N__12623),
            .sr(N__12506));
    defparam \receive_module.rx_counter.FRAME_COUNTER_244__i3_LC_13_6_3 .C_ON=1'b1;
    defparam \receive_module.rx_counter.FRAME_COUNTER_244__i3_LC_13_6_3 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.FRAME_COUNTER_244__i3_LC_13_6_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.FRAME_COUNTER_244__i3_LC_13_6_3  (
            .in0(_gnd_net_),
            .in1(N__12551),
            .in2(_gnd_net_),
            .in3(N__11630),
            .lcout(\receive_module.rx_counter.FRAME_COUNTER_3 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3158 ),
            .carryout(\receive_module.rx_counter.n3159 ),
            .clk(N__24576),
            .ce(N__12623),
            .sr(N__12506));
    defparam \receive_module.rx_counter.FRAME_COUNTER_244__i4_LC_13_6_4 .C_ON=1'b1;
    defparam \receive_module.rx_counter.FRAME_COUNTER_244__i4_LC_13_6_4 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.FRAME_COUNTER_244__i4_LC_13_6_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.FRAME_COUNTER_244__i4_LC_13_6_4  (
            .in0(_gnd_net_),
            .in1(N__12611),
            .in2(_gnd_net_),
            .in3(N__12629),
            .lcout(\receive_module.rx_counter.FRAME_COUNTER_4 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3159 ),
            .carryout(\receive_module.rx_counter.n3160 ),
            .clk(N__24576),
            .ce(N__12623),
            .sr(N__12506));
    defparam \receive_module.rx_counter.FRAME_COUNTER_244__i5_LC_13_6_5 .C_ON=1'b0;
    defparam \receive_module.rx_counter.FRAME_COUNTER_244__i5_LC_13_6_5 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.FRAME_COUNTER_244__i5_LC_13_6_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.FRAME_COUNTER_244__i5_LC_13_6_5  (
            .in0(_gnd_net_),
            .in1(N__12587),
            .in2(_gnd_net_),
            .in3(N__12626),
            .lcout(\receive_module.rx_counter.FRAME_COUNTER_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24576),
            .ce(N__12623),
            .sr(N__12506));
    defparam \receive_module.rx_counter.i1_4_lut_LC_13_7_0 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i1_4_lut_LC_13_7_0 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i1_4_lut_LC_13_7_0 .LUT_INIT=16'b1010100010001000;
    LogicCell40 \receive_module.rx_counter.i1_4_lut_LC_13_7_0  (
            .in0(N__13868),
            .in1(N__13708),
            .in2(N__13898),
            .in3(N__12701),
            .lcout(\receive_module.rx_counter.n4_adj_605 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i1_2_lut_adj_22_LC_13_7_1 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i1_2_lut_adj_22_LC_13_7_1 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i1_2_lut_adj_22_LC_13_7_1 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \receive_module.rx_counter.i1_2_lut_adj_22_LC_13_7_1  (
            .in0(_gnd_net_),
            .in1(N__12610),
            .in2(_gnd_net_),
            .in3(N__12598),
            .lcout(\receive_module.rx_counter.n7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.old_VS_52_LC_13_7_2 .C_ON=1'b0;
    defparam \receive_module.rx_counter.old_VS_52_LC_13_7_2 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.old_VS_52_LC_13_7_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \receive_module.rx_counter.old_VS_52_LC_13_7_2  (
            .in0(N__13087),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\receive_module.rx_counter.old_VS ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24583),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i2130_2_lut_LC_13_7_5 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i2130_2_lut_LC_13_7_5 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i2130_2_lut_LC_13_7_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \receive_module.rx_counter.i2130_2_lut_LC_13_7_5  (
            .in0(_gnd_net_),
            .in1(N__12586),
            .in2(_gnd_net_),
            .in3(N__12574),
            .lcout(),
            .ltout(\receive_module.rx_counter.n3473_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i5_4_lut_LC_13_7_6 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i5_4_lut_LC_13_7_6 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i5_4_lut_LC_13_7_6 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \receive_module.rx_counter.i5_4_lut_LC_13_7_6  (
            .in0(N__12562),
            .in1(N__12550),
            .in2(N__12539),
            .in3(N__12536),
            .lcout(\receive_module.rx_counter.n11 ),
            .ltout(\receive_module.rx_counter.n11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i1281_2_lut_3_lut_LC_13_7_7 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i1281_2_lut_3_lut_LC_13_7_7 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i1281_2_lut_3_lut_LC_13_7_7 .LUT_INIT=16'b0000000000001100;
    LogicCell40 \receive_module.rx_counter.i1281_2_lut_3_lut_LC_13_7_7  (
            .in0(_gnd_net_),
            .in1(N__12520),
            .in2(N__12509),
            .in3(N__13086),
            .lcout(\receive_module.rx_counter.n2529 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i3_4_lut_LC_13_8_0 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i3_4_lut_LC_13_8_0 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i3_4_lut_LC_13_8_0 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \receive_module.rx_counter.i3_4_lut_LC_13_8_0  (
            .in0(N__12641),
            .in1(N__12713),
            .in2(N__13769),
            .in3(N__12707),
            .lcout(),
            .ltout(\receive_module.rx_counter.n3422_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.O_VISIBLE_53_LC_13_8_1 .C_ON=1'b0;
    defparam \receive_module.rx_counter.O_VISIBLE_53_LC_13_8_1 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.O_VISIBLE_53_LC_13_8_1 .LUT_INIT=16'b0000000001110000;
    LogicCell40 \receive_module.rx_counter.O_VISIBLE_53_LC_13_8_1  (
            .in0(N__12728),
            .in1(N__13768),
            .in2(N__12722),
            .in3(N__12719),
            .lcout(RX_WE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24587),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i2_3_lut_LC_13_8_2 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i2_3_lut_LC_13_8_2 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i2_3_lut_LC_13_8_2 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \receive_module.rx_counter.i2_3_lut_LC_13_8_2  (
            .in0(N__13736),
            .in1(N__13838),
            .in2(_gnd_net_),
            .in3(N__13788),
            .lcout(\receive_module.rx_counter.n3394 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i1_2_lut_3_lut_LC_13_8_3 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i1_2_lut_3_lut_LC_13_8_3 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i1_2_lut_3_lut_LC_13_8_3 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \receive_module.rx_counter.i1_2_lut_3_lut_LC_13_8_3  (
            .in0(N__13210),
            .in1(N__13862),
            .in2(_gnd_net_),
            .in3(N__13192),
            .lcout(\receive_module.rx_counter.n5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i2_4_lut_LC_13_8_4 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i2_4_lut_LC_13_8_4 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i2_4_lut_LC_13_8_4 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \receive_module.rx_counter.i2_4_lut_LC_13_8_4  (
            .in0(N__13735),
            .in1(N__13811),
            .in2(N__13841),
            .in3(N__13787),
            .lcout(\receive_module.rx_counter.n3413 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_13_LC_13_8_5 .C_ON=1'b0;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_13_LC_13_8_5 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_13_LC_13_8_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \line_buffer.i1_2_lut_3_lut_4_lut_adj_13_LC_13_8_5  (
            .in0(N__14620),
            .in1(N__14810),
            .in2(N__14573),
            .in3(N__14471),
            .lcout(\line_buffer.n596 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i595_2_lut_rep_27_LC_13_8_6 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i595_2_lut_rep_27_LC_13_8_6 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i595_2_lut_rep_27_LC_13_8_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \receive_module.rx_counter.i595_2_lut_rep_27_LC_13_8_6  (
            .in0(_gnd_net_),
            .in1(N__13191),
            .in2(_gnd_net_),
            .in3(N__13209),
            .lcout(\receive_module.rx_counter.n3633 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i1_2_lut_adj_21_LC_13_8_7 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i1_2_lut_adj_21_LC_13_8_7 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i1_2_lut_adj_21_LC_13_8_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \receive_module.rx_counter.i1_2_lut_adj_21_LC_13_8_7  (
            .in0(N__13812),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13889),
            .lcout(\receive_module.rx_counter.n4_adj_604 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.Y__i0_LC_13_9_0 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i0_LC_13_9_0 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i0_LC_13_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i0_LC_13_9_0  (
            .in0(_gnd_net_),
            .in1(N__13733),
            .in2(_gnd_net_),
            .in3(N__12635),
            .lcout(\receive_module.rx_counter.Y_0 ),
            .ltout(),
            .carryin(bfn_13_9_0_),
            .carryout(\receive_module.rx_counter.n3117 ),
            .clk(N__24592),
            .ce(N__13166),
            .sr(N__12771));
    defparam \receive_module.rx_counter.Y__i1_LC_13_9_1 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i1_LC_13_9_1 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i1_LC_13_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i1_LC_13_9_1  (
            .in0(_gnd_net_),
            .in1(N__13839),
            .in2(_gnd_net_),
            .in3(N__12632),
            .lcout(\receive_module.rx_counter.Y_1 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3117 ),
            .carryout(\receive_module.rx_counter.n3118 ),
            .clk(N__24592),
            .ce(N__13166),
            .sr(N__12771));
    defparam \receive_module.rx_counter.Y__i2_LC_13_9_2 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i2_LC_13_9_2 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i2_LC_13_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i2_LC_13_9_2  (
            .in0(_gnd_net_),
            .in1(N__13789),
            .in2(_gnd_net_),
            .in3(N__13220),
            .lcout(\receive_module.rx_counter.Y_2 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3118 ),
            .carryout(\receive_module.rx_counter.n3119 ),
            .clk(N__24592),
            .ce(N__13166),
            .sr(N__12771));
    defparam \receive_module.rx_counter.Y__i3_LC_13_9_3 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i3_LC_13_9_3 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i3_LC_13_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i3_LC_13_9_3  (
            .in0(_gnd_net_),
            .in1(N__13813),
            .in2(_gnd_net_),
            .in3(N__13217),
            .lcout(\receive_module.rx_counter.Y_3 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3119 ),
            .carryout(\receive_module.rx_counter.n3120 ),
            .clk(N__24592),
            .ce(N__13166),
            .sr(N__12771));
    defparam \receive_module.rx_counter.Y__i4_LC_13_9_4 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i4_LC_13_9_4 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i4_LC_13_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i4_LC_13_9_4  (
            .in0(_gnd_net_),
            .in1(N__13890),
            .in2(_gnd_net_),
            .in3(N__13214),
            .lcout(\receive_module.rx_counter.Y_4 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3120 ),
            .carryout(\receive_module.rx_counter.n3121 ),
            .clk(N__24592),
            .ce(N__13166),
            .sr(N__12771));
    defparam \receive_module.rx_counter.Y__i5_LC_13_9_5 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i5_LC_13_9_5 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i5_LC_13_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i5_LC_13_9_5  (
            .in0(_gnd_net_),
            .in1(N__13211),
            .in2(_gnd_net_),
            .in3(N__13196),
            .lcout(\receive_module.rx_counter.Y_5 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3121 ),
            .carryout(\receive_module.rx_counter.n3122 ),
            .clk(N__24592),
            .ce(N__13166),
            .sr(N__12771));
    defparam \receive_module.rx_counter.Y__i6_LC_13_9_6 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i6_LC_13_9_6 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i6_LC_13_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i6_LC_13_9_6  (
            .in0(_gnd_net_),
            .in1(N__13193),
            .in2(_gnd_net_),
            .in3(N__13175),
            .lcout(\receive_module.rx_counter.Y_6 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3122 ),
            .carryout(\receive_module.rx_counter.n3123 ),
            .clk(N__24592),
            .ce(N__13166),
            .sr(N__12771));
    defparam \receive_module.rx_counter.Y__i7_LC_13_9_7 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i7_LC_13_9_7 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i7_LC_13_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i7_LC_13_9_7  (
            .in0(_gnd_net_),
            .in1(N__13867),
            .in2(_gnd_net_),
            .in3(N__13172),
            .lcout(\receive_module.rx_counter.Y_7 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3123 ),
            .carryout(\receive_module.rx_counter.n3124 ),
            .clk(N__24592),
            .ce(N__13166),
            .sr(N__12771));
    defparam \receive_module.rx_counter.Y__i8_LC_13_10_0 .C_ON=1'b0;
    defparam \receive_module.rx_counter.Y__i8_LC_13_10_0 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i8_LC_13_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i8_LC_13_10_0  (
            .in0(_gnd_net_),
            .in1(N__13763),
            .in2(_gnd_net_),
            .in3(N__13169),
            .lcout(\receive_module.rx_counter.Y_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24596),
            .ce(N__13165),
            .sr(N__12760));
    defparam \receive_module.BRAM_ADDR__i2_LC_13_11_0 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i2_LC_13_11_0 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i2_LC_13_11_0 .LUT_INIT=16'b1010110010101010;
    LogicCell40 \receive_module.BRAM_ADDR__i2_LC_13_11_0  (
            .in0(N__13148),
            .in1(N__12830),
            .in2(N__14669),
            .in3(N__13095),
            .lcout(RX_ADDR_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24600),
            .ce(),
            .sr(N__12772));
    defparam \transmit_module.video_signal_controller.VGA_Y_i0_LC_13_12_0 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i0_LC_13_12_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i0_LC_13_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i0_LC_13_12_0  (
            .in0(_gnd_net_),
            .in1(N__14873),
            .in2(_gnd_net_),
            .in3(N__12731),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_0 ),
            .ltout(),
            .carryin(bfn_13_12_0_),
            .carryout(\transmit_module.video_signal_controller.n3136 ),
            .clk(N__23501),
            .ce(N__14247),
            .sr(N__14203));
    defparam \transmit_module.video_signal_controller.VGA_Y_i1_LC_13_12_1 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i1_LC_13_12_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i1_LC_13_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i1_LC_13_12_1  (
            .in0(_gnd_net_),
            .in1(N__14896),
            .in2(_gnd_net_),
            .in3(N__13247),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_1 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3136 ),
            .carryout(\transmit_module.video_signal_controller.n3137 ),
            .clk(N__23501),
            .ce(N__14247),
            .sr(N__14203));
    defparam \transmit_module.video_signal_controller.VGA_Y_i2_LC_13_12_2 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i2_LC_13_12_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i2_LC_13_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i2_LC_13_12_2  (
            .in0(_gnd_net_),
            .in1(N__15381),
            .in2(_gnd_net_),
            .in3(N__13244),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_2 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3137 ),
            .carryout(\transmit_module.video_signal_controller.n3138 ),
            .clk(N__23501),
            .ce(N__14247),
            .sr(N__14203));
    defparam \transmit_module.video_signal_controller.VGA_Y_i3_LC_13_12_3 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i3_LC_13_12_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i3_LC_13_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i3_LC_13_12_3  (
            .in0(_gnd_net_),
            .in1(N__14922),
            .in2(_gnd_net_),
            .in3(N__13241),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_3 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3138 ),
            .carryout(\transmit_module.video_signal_controller.n3139 ),
            .clk(N__23501),
            .ce(N__14247),
            .sr(N__14203));
    defparam \transmit_module.video_signal_controller.VGA_Y_i4_LC_13_12_4 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i4_LC_13_12_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i4_LC_13_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i4_LC_13_12_4  (
            .in0(_gnd_net_),
            .in1(N__15528),
            .in2(_gnd_net_),
            .in3(N__13238),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_4 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3139 ),
            .carryout(\transmit_module.video_signal_controller.n3140 ),
            .clk(N__23501),
            .ce(N__14247),
            .sr(N__14203));
    defparam \transmit_module.video_signal_controller.VGA_Y_i5_LC_13_12_5 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i5_LC_13_12_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i5_LC_13_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i5_LC_13_12_5  (
            .in0(_gnd_net_),
            .in1(N__14955),
            .in2(_gnd_net_),
            .in3(N__13235),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_5 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3140 ),
            .carryout(\transmit_module.video_signal_controller.n3141 ),
            .clk(N__23501),
            .ce(N__14247),
            .sr(N__14203));
    defparam \transmit_module.video_signal_controller.VGA_Y_i6_LC_13_12_6 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i6_LC_13_12_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i6_LC_13_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i6_LC_13_12_6  (
            .in0(_gnd_net_),
            .in1(N__15012),
            .in2(_gnd_net_),
            .in3(N__13232),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_6 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3141 ),
            .carryout(\transmit_module.video_signal_controller.n3142 ),
            .clk(N__23501),
            .ce(N__14247),
            .sr(N__14203));
    defparam \transmit_module.video_signal_controller.VGA_Y_i7_LC_13_12_7 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i7_LC_13_12_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i7_LC_13_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i7_LC_13_12_7  (
            .in0(_gnd_net_),
            .in1(N__15048),
            .in2(_gnd_net_),
            .in3(N__13229),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_7 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3142 ),
            .carryout(\transmit_module.video_signal_controller.n3143 ),
            .clk(N__23501),
            .ce(N__14247),
            .sr(N__14203));
    defparam \transmit_module.video_signal_controller.VGA_Y_i8_LC_13_13_0 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i8_LC_13_13_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i8_LC_13_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i8_LC_13_13_0  (
            .in0(_gnd_net_),
            .in1(N__15073),
            .in2(_gnd_net_),
            .in3(N__13226),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_8 ),
            .ltout(),
            .carryin(bfn_13_13_0_),
            .carryout(\transmit_module.video_signal_controller.n3144 ),
            .clk(N__23364),
            .ce(N__14246),
            .sr(N__14207));
    defparam \transmit_module.video_signal_controller.VGA_Y_i9_LC_13_13_1 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i9_LC_13_13_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i9_LC_13_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i9_LC_13_13_1  (
            .in0(_gnd_net_),
            .in1(N__15488),
            .in2(_gnd_net_),
            .in3(N__13223),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_9 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3144 ),
            .carryout(\transmit_module.video_signal_controller.n3145 ),
            .clk(N__23364),
            .ce(N__14246),
            .sr(N__14207));
    defparam \transmit_module.video_signal_controller.VGA_Y_i10_LC_13_13_2 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i10_LC_13_13_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i10_LC_13_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i10_LC_13_13_2  (
            .in0(_gnd_net_),
            .in1(N__15429),
            .in2(_gnd_net_),
            .in3(N__13406),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_10 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3145 ),
            .carryout(\transmit_module.video_signal_controller.n3146 ),
            .clk(N__23364),
            .ce(N__14246),
            .sr(N__14207));
    defparam \transmit_module.video_signal_controller.VGA_Y_i11_LC_13_13_3 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.VGA_Y_i11_LC_13_13_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i11_LC_13_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i11_LC_13_13_3  (
            .in0(_gnd_net_),
            .in1(N__14983),
            .in2(_gnd_net_),
            .in3(N__13403),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23364),
            .ce(N__14246),
            .sr(N__14207));
    defparam \transmit_module.video_signal_controller.i485_4_lut_LC_13_14_0 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i485_4_lut_LC_13_14_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i485_4_lut_LC_13_14_0 .LUT_INIT=16'b1111100000000000;
    LogicCell40 \transmit_module.video_signal_controller.i485_4_lut_LC_13_14_0  (
            .in0(N__13349),
            .in1(N__13256),
            .in2(N__13274),
            .in3(N__15352),
            .lcout(\transmit_module.video_signal_controller.n18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_17_LC_13_14_1 .C_ON=1'b0;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_17_LC_13_14_1 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_17_LC_13_14_1 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \line_buffer.i1_2_lut_3_lut_4_lut_adj_17_LC_13_14_1  (
            .in0(N__14653),
            .in1(N__14803),
            .in2(N__14565),
            .in3(N__14456),
            .lcout(\line_buffer.n564 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_2_lut_adj_26_LC_13_14_2 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_2_lut_adj_26_LC_13_14_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_2_lut_adj_26_LC_13_14_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \transmit_module.video_signal_controller.i1_2_lut_adj_26_LC_13_14_2  (
            .in0(_gnd_net_),
            .in1(N__13511),
            .in2(_gnd_net_),
            .in3(N__13655),
            .lcout(\transmit_module.video_signal_controller.n3313 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_2_lut_3_lut_LC_13_14_3 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_2_lut_3_lut_LC_13_14_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_2_lut_3_lut_LC_13_14_3 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \transmit_module.video_signal_controller.i1_2_lut_3_lut_LC_13_14_3  (
            .in0(N__15304),
            .in1(N__13631),
            .in2(_gnd_net_),
            .in3(N__13538),
            .lcout(\transmit_module.video_signal_controller.n2001 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1585_2_lut_rep_18_LC_13_14_4 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1585_2_lut_rep_18_LC_13_14_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1585_2_lut_rep_18_LC_13_14_4 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \transmit_module.video_signal_controller.i1585_2_lut_rep_18_LC_13_14_4  (
            .in0(N__13310),
            .in1(_gnd_net_),
            .in2(N__13342),
            .in3(_gnd_net_),
            .lcout(\transmit_module.video_signal_controller.n3624 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1669_2_lut_3_lut_LC_13_14_5 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1669_2_lut_3_lut_LC_13_14_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1669_2_lut_3_lut_LC_13_14_5 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \transmit_module.video_signal_controller.i1669_2_lut_3_lut_LC_13_14_5  (
            .in0(N__13343),
            .in1(N__13311),
            .in2(_gnd_net_),
            .in3(N__13290),
            .lcout(),
            .ltout(\transmit_module.video_signal_controller.n2917_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1699_4_lut_LC_13_14_6 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1699_4_lut_LC_13_14_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1699_4_lut_LC_13_14_6 .LUT_INIT=16'b1100100010001000;
    LogicCell40 \transmit_module.video_signal_controller.i1699_4_lut_LC_13_14_6  (
            .in0(N__13270),
            .in1(N__15351),
            .in2(N__13259),
            .in3(N__13255),
            .lcout(),
            .ltout(\transmit_module.video_signal_controller.n2947_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1705_4_lut_LC_13_14_7 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1705_4_lut_LC_13_14_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1705_4_lut_LC_13_14_7 .LUT_INIT=16'b1111111010101010;
    LogicCell40 \transmit_module.video_signal_controller.i1705_4_lut_LC_13_14_7  (
            .in0(N__16717),
            .in1(N__13604),
            .in2(N__13697),
            .in3(N__13577),
            .lcout(\transmit_module.video_signal_controller.n2036 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n3591_bdd_4_lut_LC_13_15_0 .C_ON=1'b0;
    defparam \line_buffer.n3591_bdd_4_lut_LC_13_15_0 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3591_bdd_4_lut_LC_13_15_0 .LUT_INIT=16'b1101110010011000;
    LogicCell40 \line_buffer.n3591_bdd_4_lut_LC_13_15_0  (
            .in0(N__23806),
            .in1(N__13412),
            .in2(N__13694),
            .in3(N__13676),
            .lcout(\line_buffer.n3594 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_4_lut_adj_25_LC_13_15_2 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_4_lut_adj_25_LC_13_15_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_4_lut_adj_25_LC_13_15_2 .LUT_INIT=16'b1111111010101010;
    LogicCell40 \transmit_module.video_signal_controller.i1_4_lut_adj_25_LC_13_15_2  (
            .in0(N__13541),
            .in1(N__13512),
            .in2(N__13661),
            .in3(N__13633),
            .lcout(\transmit_module.video_signal_controller.n4_adj_617 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i2_4_lut_4_lut_LC_13_15_3 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i2_4_lut_4_lut_LC_13_15_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i2_4_lut_4_lut_LC_13_15_3 .LUT_INIT=16'b0101011101010110;
    LogicCell40 \transmit_module.video_signal_controller.i2_4_lut_4_lut_LC_13_15_3  (
            .in0(N__13572),
            .in1(N__13610),
            .in2(N__13603),
            .in3(N__16711),
            .lcout(\transmit_module.video_signal_controller.n7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i2_3_lut_rep_19_LC_13_15_5 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i2_3_lut_rep_19_LC_13_15_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i2_3_lut_rep_19_LC_13_15_5 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \transmit_module.video_signal_controller.i2_3_lut_rep_19_LC_13_15_5  (
            .in0(N__13595),
            .in1(N__13568),
            .in2(_gnd_net_),
            .in3(N__16712),
            .lcout(),
            .ltout(\transmit_module.video_signal_controller.n3625_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i2128_4_lut_LC_13_15_6 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i2128_4_lut_LC_13_15_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i2128_4_lut_LC_13_15_6 .LUT_INIT=16'b1111110011111000;
    LogicCell40 \transmit_module.video_signal_controller.i2128_4_lut_LC_13_15_6  (
            .in0(N__13547),
            .in1(N__13540),
            .in2(N__13517),
            .in3(N__13513),
            .lcout(\transmit_module.video_signal_controller.n3471 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_12_LC_13_15_7 .C_ON=1'b0;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_12_LC_13_15_7 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_12_LC_13_15_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \line_buffer.i1_2_lut_3_lut_4_lut_adj_12_LC_13_15_7  (
            .in0(N__14654),
            .in1(N__14799),
            .in2(N__14566),
            .in3(N__14460),
            .lcout(\line_buffer.n597 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2245_LC_13_16_1 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2245_LC_13_16_1 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2245_LC_13_16_1 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_2245_LC_13_16_1  (
            .in0(N__24339),
            .in1(N__13445),
            .in2(N__23841),
            .in3(N__13427),
            .lcout(\line_buffer.n3591 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_22_LC_13_16_7 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_22_LC_13_16_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_22_LC_13_16_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \transmit_module.video_signal_controller.i1_2_lut_rep_22_LC_13_16_7  (
            .in0(_gnd_net_),
            .in1(N__14900),
            .in2(_gnd_net_),
            .in3(N__15385),
            .lcout(\transmit_module.video_signal_controller.n3628 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_16_LC_13_17_0 .C_ON=1'b0;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_16_LC_13_17_0 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_16_LC_13_17_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \line_buffer.i1_2_lut_3_lut_4_lut_adj_16_LC_13_17_0  (
            .in0(N__14811),
            .in1(N__14655),
            .in2(N__14574),
            .in3(N__14472),
            .lcout(\line_buffer.n468 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i4_3_lut_LC_13_18_6 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i4_3_lut_LC_13_18_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i4_3_lut_LC_13_18_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_12_i4_3_lut_LC_13_18_6  (
            .in0(N__20635),
            .in1(N__13916),
            .in2(_gnd_net_),
            .in3(N__16501),
            .lcout(\transmit_module.n113 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1612_4_lut_LC_13_19_3 .C_ON=1'b0;
    defparam \transmit_module.i1612_4_lut_LC_13_19_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1612_4_lut_LC_13_19_3 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \transmit_module.i1612_4_lut_LC_13_19_3  (
            .in0(N__20763),
            .in1(N__20016),
            .in2(N__14857),
            .in3(N__15268),
            .lcout(n25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.ADDR_Y_COMPONENT__i3_LC_13_19_6 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i3_LC_13_19_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i3_LC_13_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i3_LC_13_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16505),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22976),
            .ce(N__20454),
            .sr(N__20240));
    defparam \tvp_video_buffer.BUFFER_0__i11_LC_14_4_0 .C_ON=1'b0;
    defparam \tvp_video_buffer.BUFFER_0__i11_LC_14_4_0 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.BUFFER_0__i11_LC_14_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.BUFFER_0__i11_LC_14_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13910),
            .lcout(\tvp_video_buffer.BUFFER_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24565),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i2_2_lut_LC_14_8_0 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i2_2_lut_LC_14_8_0 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i2_2_lut_LC_14_8_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \receive_module.rx_counter.i2_2_lut_LC_14_8_0  (
            .in0(_gnd_net_),
            .in1(N__13891),
            .in2(_gnd_net_),
            .in3(N__13863),
            .lcout(\receive_module.rx_counter.n10_adj_610 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i6_4_lut_LC_14_8_5 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i6_4_lut_LC_14_8_5 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i6_4_lut_LC_14_8_5 .LUT_INIT=16'b1111111110111111;
    LogicCell40 \receive_module.rx_counter.i6_4_lut_LC_14_8_5  (
            .in0(N__13840),
            .in1(N__13814),
            .in2(N__13793),
            .in3(N__13764),
            .lcout(),
            .ltout(\receive_module.rx_counter.n14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.SYNC_46_LC_14_8_6 .C_ON=1'b0;
    defparam \receive_module.rx_counter.SYNC_46_LC_14_8_6 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.SYNC_46_LC_14_8_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \receive_module.rx_counter.SYNC_46_LC_14_8_6  (
            .in0(N__13742),
            .in1(N__13734),
            .in2(N__13712),
            .in3(N__13709),
            .lcout(RX_TX_SYNC),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24584),
            .ce(),
            .sr(_gnd_net_));
    defparam \sync_buffer.BUFFER_0__i2_LC_14_9_2 .C_ON=1'b0;
    defparam \sync_buffer.BUFFER_0__i2_LC_14_9_2 .SEQ_MODE=4'b1000;
    defparam \sync_buffer.BUFFER_0__i2_LC_14_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sync_buffer.BUFFER_0__i2_LC_14_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14819),
            .lcout(\sync_buffer.BUFFER_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23507),
            .ce(),
            .sr(_gnd_net_));
    defparam \sync_buffer.BUFFER_0__i1_LC_14_9_3 .C_ON=1'b0;
    defparam \sync_buffer.BUFFER_0__i1_LC_14_9_3 .SEQ_MODE=4'b1000;
    defparam \sync_buffer.BUFFER_0__i1_LC_14_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sync_buffer.BUFFER_0__i1_LC_14_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14825),
            .lcout(\sync_buffer.BUFFER_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23507),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_11_LC_14_9_4 .C_ON=1'b0;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_11_LC_14_9_4 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_11_LC_14_9_4 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \line_buffer.i1_2_lut_3_lut_4_lut_adj_11_LC_14_9_4  (
            .in0(N__14813),
            .in1(N__14621),
            .in2(N__14576),
            .in3(N__14473),
            .lcout(\line_buffer.n532 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.WIRE_OUT_i1_LC_14_11_5 .C_ON=1'b0;
    defparam \tvp_video_buffer.WIRE_OUT_i1_LC_14_11_5 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.WIRE_OUT_i1_LC_14_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.WIRE_OUT_i1_LC_14_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14360),
            .lcout(RX_DATA_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24597),
            .ce(),
            .sr(_gnd_net_));
    defparam \sync_buffer.WIRE_OUT_0__9_LC_14_12_3 .C_ON=1'b0;
    defparam \sync_buffer.WIRE_OUT_0__9_LC_14_12_3 .SEQ_MODE=4'b1000;
    defparam \sync_buffer.WIRE_OUT_0__9_LC_14_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sync_buffer.WIRE_OUT_0__9_LC_14_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14267),
            .lcout(RX_TX_SYNC_BUFF),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23463),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1138_2_lut_LC_14_12_7 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1138_2_lut_LC_14_12_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1138_2_lut_LC_14_12_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \transmit_module.video_signal_controller.i1138_2_lut_LC_14_12_7  (
            .in0(_gnd_net_),
            .in1(N__14258),
            .in2(_gnd_net_),
            .in3(N__14239),
            .lcout(\transmit_module.video_signal_controller.n2378 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_2_lut_3_lut_adj_28_LC_14_13_0 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_2_lut_3_lut_adj_28_LC_14_13_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_2_lut_3_lut_adj_28_LC_14_13_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \transmit_module.video_signal_controller.i1_2_lut_3_lut_adj_28_LC_14_13_0  (
            .in0(N__14916),
            .in1(N__14891),
            .in2(_gnd_net_),
            .in3(N__15377),
            .lcout(),
            .ltout(\transmit_module.video_signal_controller.n49_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i2_4_lut_LC_14_13_1 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i2_4_lut_LC_14_13_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i2_4_lut_LC_14_13_1 .LUT_INIT=16'b1100100000000000;
    LogicCell40 \transmit_module.video_signal_controller.i2_4_lut_LC_14_13_1  (
            .in0(N__15527),
            .in1(N__14954),
            .in2(N__14186),
            .in3(N__15005),
            .lcout(\transmit_module.video_signal_controller.n3412 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i0_LC_14_13_3 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i0_LC_14_13_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i0_LC_14_13_3 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \transmit_module.BRAM_ADDR__i0_LC_14_13_3  (
            .in0(N__20855),
            .in1(N__16097),
            .in2(N__20288),
            .in3(N__16081),
            .lcout(\transmit_module.TX_ADDR_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23485),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_2_lut_adj_23_LC_14_13_5 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_2_lut_adj_23_LC_14_13_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_2_lut_adj_23_LC_14_13_5 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \transmit_module.video_signal_controller.i1_2_lut_adj_23_LC_14_13_5  (
            .in0(N__14892),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14872),
            .lcout(\transmit_module.video_signal_controller.n45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i1_LC_14_13_7 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i1_LC_14_13_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i1_LC_14_13_7 .LUT_INIT=16'b0000000010101100;
    LogicCell40 \transmit_module.BRAM_ADDR__i1_LC_14_13_7  (
            .in0(N__15851),
            .in1(N__15826),
            .in2(N__20875),
            .in3(N__20259),
            .lcout(\transmit_module.TX_ADDR_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23485),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_14_i2_3_lut_LC_14_14_0 .C_ON=1'b0;
    defparam \transmit_module.mux_14_i2_3_lut_LC_14_14_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_14_i2_3_lut_LC_14_14_0 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \transmit_module.mux_14_i2_3_lut_LC_14_14_0  (
            .in0(N__21612),
            .in1(_gnd_net_),
            .in2(N__16520),
            .in3(N__18282),
            .lcout(\transmit_module.n146 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i2124_2_lut_rep_16_3_lut_LC_14_14_2 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i2124_2_lut_rep_16_3_lut_LC_14_14_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i2124_2_lut_rep_16_3_lut_LC_14_14_2 .LUT_INIT=16'b1111111111111010;
    LogicCell40 \transmit_module.video_signal_controller.i2124_2_lut_rep_16_3_lut_LC_14_14_2  (
            .in0(N__15052),
            .in1(_gnd_net_),
            .in2(N__15017),
            .in3(N__15072),
            .lcout(\transmit_module.video_signal_controller.n3622 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i3_LC_14_14_3 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i3_LC_14_14_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i3_LC_14_14_3 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \transmit_module.BRAM_ADDR__i3_LC_14_14_3  (
            .in0(N__20869),
            .in1(N__14861),
            .in2(N__20258),
            .in3(N__15275),
            .lcout(\transmit_module.TX_ADDR_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23379),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_14_i6_3_lut_LC_14_14_4 .C_ON=1'b0;
    defparam \transmit_module.mux_14_i6_3_lut_LC_14_14_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_14_i6_3_lut_LC_14_14_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \transmit_module.mux_14_i6_3_lut_LC_14_14_4  (
            .in0(N__21613),
            .in1(N__16451),
            .in2(_gnd_net_),
            .in3(N__17015),
            .lcout(\transmit_module.n142 ),
            .ltout(\transmit_module.n142_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i5_LC_14_14_5 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i5_LC_14_14_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i5_LC_14_14_5 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \transmit_module.BRAM_ADDR__i5_LC_14_14_5  (
            .in0(N__20870),
            .in1(N__20189),
            .in2(N__14840),
            .in3(N__16991),
            .lcout(\transmit_module.TX_ADDR_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23379),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_14_i1_3_lut_LC_14_14_6 .C_ON=1'b0;
    defparam \transmit_module.mux_14_i1_3_lut_LC_14_14_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_14_i1_3_lut_LC_14_14_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \transmit_module.mux_14_i1_3_lut_LC_14_14_6  (
            .in0(N__21611),
            .in1(N__16526),
            .in2(_gnd_net_),
            .in3(N__16551),
            .lcout(\transmit_module.n147 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i6_4_lut_LC_14_14_7 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i6_4_lut_LC_14_14_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i6_4_lut_LC_14_14_7 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \transmit_module.video_signal_controller.i6_4_lut_LC_14_14_7  (
            .in0(N__15532),
            .in1(N__14959),
            .in2(N__14837),
            .in3(N__14982),
            .lcout(\transmit_module.video_signal_controller.n16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_4_lut_LC_14_15_0 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_4_lut_LC_14_15_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_4_lut_LC_14_15_0 .LUT_INIT=16'b1111110011101100;
    LogicCell40 \transmit_module.video_signal_controller.i1_4_lut_LC_14_15_0  (
            .in0(N__15026),
            .in1(N__15460),
            .in2(N__15496),
            .in3(N__15083),
            .lcout(\transmit_module.video_signal_controller.n3333 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1608_2_lut_rep_20_LC_14_15_2 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1608_2_lut_rep_20_LC_14_15_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1608_2_lut_rep_20_LC_14_15_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \transmit_module.video_signal_controller.i1608_2_lut_rep_20_LC_14_15_2  (
            .in0(_gnd_net_),
            .in1(N__15074),
            .in2(_gnd_net_),
            .in3(N__15053),
            .lcout(\transmit_module.video_signal_controller.n3626 ),
            .ltout(\transmit_module.video_signal_controller.n3626_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i2134_3_lut_4_lut_LC_14_15_3 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i2134_3_lut_4_lut_LC_14_15_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i2134_3_lut_4_lut_LC_14_15_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \transmit_module.video_signal_controller.i2134_3_lut_4_lut_LC_14_15_3  (
            .in0(N__15492),
            .in1(N__15016),
            .in2(N__14987),
            .in3(N__14930),
            .lcout(\transmit_module.video_signal_controller.n3477 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_2_lut_LC_14_15_4 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_2_lut_LC_14_15_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_2_lut_LC_14_15_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \transmit_module.video_signal_controller.i1_2_lut_LC_14_15_4  (
            .in0(_gnd_net_),
            .in1(N__14984),
            .in2(_gnd_net_),
            .in3(N__15430),
            .lcout(\transmit_module.video_signal_controller.n3331 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_14_i11_3_lut_LC_14_15_5 .C_ON=1'b0;
    defparam \transmit_module.mux_14_i11_3_lut_LC_14_15_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_14_i11_3_lut_LC_14_15_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_14_i11_3_lut_LC_14_15_5  (
            .in0(N__21585),
            .in1(N__16665),
            .in2(_gnd_net_),
            .in3(N__16610),
            .lcout(\transmit_module.n137 ),
            .ltout(\transmit_module.n137_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i10_LC_14_15_6 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i10_LC_14_15_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i10_LC_14_15_6 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \transmit_module.BRAM_ADDR__i10_LC_14_15_6  (
            .in0(N__20123),
            .in1(N__20824),
            .in2(N__14963),
            .in3(N__16642),
            .lcout(\transmit_module.TX_ADDR_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23131),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.ADDR_Y_COMPONENT__i0_LC_14_16_0 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i0_LC_14_16_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i0_LC_14_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i0_LC_14_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16553),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23397),
            .ce(N__20444),
            .sr(N__20186));
    defparam \transmit_module.ADDR_Y_COMPONENT__i10_LC_14_16_2 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i10_LC_14_16_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i10_LC_14_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i10_LC_14_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16667),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23397),
            .ce(N__20444),
            .sr(N__20186));
    defparam \transmit_module.ADDR_Y_COMPONENT__i5_LC_14_16_7 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i5_LC_14_16_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i5_LC_14_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i5_LC_14_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17021),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23397),
            .ce(N__20444),
            .sr(N__20186));
    defparam \transmit_module.video_signal_controller.i1_4_lut_adj_27_LC_14_17_0 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_4_lut_adj_27_LC_14_17_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_4_lut_adj_27_LC_14_17_0 .LUT_INIT=16'b1111101011101010;
    LogicCell40 \transmit_module.video_signal_controller.i1_4_lut_adj_27_LC_14_17_0  (
            .in0(N__14960),
            .in1(N__14929),
            .in2(N__15536),
            .in3(N__15503),
            .lcout(),
            .ltout(\transmit_module.video_signal_controller.n7_adj_618_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i5_4_lut_LC_14_17_1 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i5_4_lut_LC_14_17_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i5_4_lut_LC_14_17_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \transmit_module.video_signal_controller.i5_4_lut_LC_14_17_1  (
            .in0(N__15497),
            .in1(N__15464),
            .in2(N__15449),
            .in3(N__15446),
            .lcout(\transmit_module.video_signal_controller.VGA_VISIBLE_N_580 ),
            .ltout(\transmit_module.video_signal_controller.VGA_VISIBLE_N_580_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.VGA_VISIBLE_Y_64_LC_14_17_2 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.VGA_VISIBLE_Y_64_LC_14_17_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_VISIBLE_Y_64_LC_14_17_2 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \transmit_module.video_signal_controller.VGA_VISIBLE_Y_64_LC_14_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15437),
            .in3(N__16736),
            .lcout(\transmit_module.VGA_VISIBLE_Y ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23335),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.VGA_VS_67_LC_14_17_3 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.VGA_VS_67_LC_14_17_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_VS_67_LC_14_17_3 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \transmit_module.video_signal_controller.VGA_VS_67_LC_14_17_3  (
            .in0(N__15434),
            .in1(N__15410),
            .in2(N__15401),
            .in3(N__15389),
            .lcout(ADV_VSYNC_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23335),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i123_2_lut_4_lut_LC_14_17_4 .C_ON=1'b0;
    defparam \transmit_module.i123_2_lut_4_lut_LC_14_17_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i123_2_lut_4_lut_LC_14_17_4 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \transmit_module.i123_2_lut_4_lut_LC_14_17_4  (
            .in0(N__16423),
            .in1(N__16399),
            .in2(N__20121),
            .in3(N__16361),
            .lcout(\transmit_module.n2167 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.old_VGA_HS_40_LC_14_17_5 .C_ON=1'b0;
    defparam \transmit_module.old_VGA_HS_40_LC_14_17_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.old_VGA_HS_40_LC_14_17_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \transmit_module.old_VGA_HS_40_LC_14_17_5  (
            .in0(N__16362),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.old_VGA_HS ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23335),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.VGA_HS_66_LC_14_17_6 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.VGA_HS_66_LC_14_17_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_HS_66_LC_14_17_6 .LUT_INIT=16'b1110111011101111;
    LogicCell40 \transmit_module.video_signal_controller.VGA_HS_66_LC_14_17_6  (
            .in0(N__15356),
            .in1(N__15329),
            .in2(N__15320),
            .in3(N__15308),
            .lcout(ADV_HSYNC_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23335),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_14_i4_3_lut_LC_14_18_2 .C_ON=1'b0;
    defparam \transmit_module.mux_14_i4_3_lut_LC_14_18_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_14_i4_3_lut_LC_14_18_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \transmit_module.mux_14_i4_3_lut_LC_14_18_2  (
            .in0(N__21607),
            .in1(N__16469),
            .in2(_gnd_net_),
            .in3(N__16494),
            .lcout(\transmit_module.n144 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i123_2_lut_4_lut_rep_30_LC_14_18_5 .C_ON=1'b0;
    defparam \transmit_module.i123_2_lut_4_lut_rep_30_LC_14_18_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i123_2_lut_4_lut_rep_30_LC_14_18_5 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \transmit_module.i123_2_lut_4_lut_rep_30_LC_14_18_5  (
            .in0(N__16422),
            .in1(N__16398),
            .in2(N__20122),
            .in3(N__16360),
            .lcout(\transmit_module.n3636 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i1_3_lut_LC_14_18_6 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i1_3_lut_LC_14_18_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i1_3_lut_LC_14_18_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_12_i1_3_lut_LC_14_18_6  (
            .in0(N__20634),
            .in1(N__16439),
            .in2(_gnd_net_),
            .in3(N__16552),
            .lcout(\transmit_module.n116 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i2_3_lut_rep_21_LC_14_18_7 .C_ON=1'b0;
    defparam \transmit_module.i2_3_lut_rep_21_LC_14_18_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i2_3_lut_rep_21_LC_14_18_7 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \transmit_module.i2_3_lut_rep_21_LC_14_18_7  (
            .in0(N__16421),
            .in1(N__16397),
            .in2(_gnd_net_),
            .in3(N__16359),
            .lcout(\transmit_module.n3627 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1619_4_lut_LC_14_19_0 .C_ON=1'b0;
    defparam \transmit_module.i1619_4_lut_LC_14_19_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1619_4_lut_LC_14_19_0 .LUT_INIT=16'b0010001100100000;
    LogicCell40 \transmit_module.i1619_4_lut_LC_14_19_0  (
            .in0(N__16643),
            .in1(N__20015),
            .in2(N__20817),
            .in3(N__16334),
            .lcout(n18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1603_4_lut_LC_14_19_1 .C_ON=1'b0;
    defparam \transmit_module.i1603_4_lut_LC_14_19_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1603_4_lut_LC_14_19_1 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \transmit_module.i1603_4_lut_LC_14_19_1  (
            .in0(N__20769),
            .in1(N__16093),
            .in2(N__20163),
            .in3(N__16082),
            .lcout(n28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i2_3_lut_LC_14_20_7 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i2_3_lut_LC_14_20_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i2_3_lut_LC_14_20_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_12_i2_3_lut_LC_14_20_7  (
            .in0(N__20655),
            .in1(N__18263),
            .in2(_gnd_net_),
            .in3(N__18295),
            .lcout(\transmit_module.n115 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1610_4_lut_LC_14_31_7 .C_ON=1'b0;
    defparam \transmit_module.i1610_4_lut_LC_14_31_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1610_4_lut_LC_14_31_7 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \transmit_module.i1610_4_lut_LC_14_31_7  (
            .in0(N__20878),
            .in1(N__15850),
            .in2(N__20328),
            .in3(N__15830),
            .lcout(n27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.BUFFER_0__i4_LC_15_5_2 .C_ON=1'b0;
    defparam \tvp_video_buffer.BUFFER_0__i4_LC_15_5_2 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.BUFFER_0__i4_LC_15_5_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \tvp_video_buffer.BUFFER_0__i4_LC_15_5_2  (
            .in0(N__15602),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\tvp_video_buffer.BUFFER_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24566),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.BUFFER_0__i5_LC_15_7_1 .C_ON=1'b0;
    defparam \tvp_video_buffer.BUFFER_0__i5_LC_15_7_1 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.BUFFER_0__i5_LC_15_7_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.BUFFER_0__i5_LC_15_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15565),
            .lcout(\tvp_video_buffer.BUFFER_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24571),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.BUFFER_0__i14_LC_15_8_3 .C_ON=1'b0;
    defparam \tvp_video_buffer.BUFFER_0__i14_LC_15_8_3 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.BUFFER_0__i14_LC_15_8_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.BUFFER_0__i14_LC_15_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16559),
            .lcout(\tvp_video_buffer.BUFFER_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24577),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.BUFFER_0__i6_LC_15_8_7 .C_ON=1'b0;
    defparam \tvp_video_buffer.BUFFER_0__i6_LC_15_8_7 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.BUFFER_0__i6_LC_15_8_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.BUFFER_0__i6_LC_15_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16576),
            .lcout(\tvp_video_buffer.BUFFER_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24577),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_2_lut_LC_15_13_0 .C_ON=1'b1;
    defparam \transmit_module.add_13_2_lut_LC_15_13_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_2_lut_LC_15_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_2_lut_LC_15_13_0  (
            .in0(_gnd_net_),
            .in1(N__16544),
            .in2(N__19673),
            .in3(_gnd_net_),
            .lcout(\transmit_module.n132 ),
            .ltout(),
            .carryin(bfn_15_13_0_),
            .carryout(\transmit_module.n3104 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_3_lut_LC_15_13_1 .C_ON=1'b1;
    defparam \transmit_module.add_13_3_lut_LC_15_13_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_3_lut_LC_15_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_3_lut_LC_15_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18288),
            .in3(N__16511),
            .lcout(\transmit_module.n131 ),
            .ltout(),
            .carryin(\transmit_module.n3104 ),
            .carryout(\transmit_module.n3105 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_4_lut_LC_15_13_2 .C_ON=1'b1;
    defparam \transmit_module.add_13_4_lut_LC_15_13_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_4_lut_LC_15_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_4_lut_LC_15_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19215),
            .in3(N__16508),
            .lcout(\transmit_module.n130 ),
            .ltout(),
            .carryin(\transmit_module.n3105 ),
            .carryout(\transmit_module.n3106 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_5_lut_LC_15_13_3 .C_ON=1'b1;
    defparam \transmit_module.add_13_5_lut_LC_15_13_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_5_lut_LC_15_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_5_lut_LC_15_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16493),
            .in3(N__16457),
            .lcout(\transmit_module.n129 ),
            .ltout(),
            .carryin(\transmit_module.n3106 ),
            .carryout(\transmit_module.n3107 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_6_lut_LC_15_13_4 .C_ON=1'b1;
    defparam \transmit_module.add_13_6_lut_LC_15_13_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_6_lut_LC_15_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_6_lut_LC_15_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20523),
            .in3(N__16454),
            .lcout(\transmit_module.n128 ),
            .ltout(),
            .carryin(\transmit_module.n3107 ),
            .carryout(\transmit_module.n3108 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_7_lut_LC_15_13_5 .C_ON=1'b1;
    defparam \transmit_module.add_13_7_lut_LC_15_13_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_7_lut_LC_15_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_7_lut_LC_15_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17020),
            .in3(N__16445),
            .lcout(\transmit_module.n127 ),
            .ltout(),
            .carryin(\transmit_module.n3108 ),
            .carryout(\transmit_module.n3109 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_8_lut_LC_15_13_6 .C_ON=1'b1;
    defparam \transmit_module.add_13_8_lut_LC_15_13_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_8_lut_LC_15_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_8_lut_LC_15_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19262),
            .in3(N__16442),
            .lcout(\transmit_module.n126 ),
            .ltout(),
            .carryin(\transmit_module.n3109 ),
            .carryout(\transmit_module.n3110 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_9_lut_LC_15_13_7 .C_ON=1'b1;
    defparam \transmit_module.add_13_9_lut_LC_15_13_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_9_lut_LC_15_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_9_lut_LC_15_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19328),
            .in3(N__16619),
            .lcout(\transmit_module.n125 ),
            .ltout(),
            .carryin(\transmit_module.n3110 ),
            .carryout(\transmit_module.n3111 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_10_lut_LC_15_14_0 .C_ON=1'b1;
    defparam \transmit_module.add_13_10_lut_LC_15_14_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_10_lut_LC_15_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_10_lut_LC_15_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17271),
            .in3(N__16616),
            .lcout(\transmit_module.n124 ),
            .ltout(),
            .carryin(bfn_15_14_0_),
            .carryout(\transmit_module.n3112 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_11_lut_LC_15_14_1 .C_ON=1'b1;
    defparam \transmit_module.add_13_11_lut_LC_15_14_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_11_lut_LC_15_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_11_lut_LC_15_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19169),
            .in3(N__16613),
            .lcout(\transmit_module.n123 ),
            .ltout(),
            .carryin(\transmit_module.n3112 ),
            .carryout(\transmit_module.n3113 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_12_lut_LC_15_14_2 .C_ON=1'b1;
    defparam \transmit_module.add_13_12_lut_LC_15_14_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_12_lut_LC_15_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_12_lut_LC_15_14_2  (
            .in0(_gnd_net_),
            .in1(N__16664),
            .in2(_gnd_net_),
            .in3(N__16604),
            .lcout(\transmit_module.n122 ),
            .ltout(),
            .carryin(\transmit_module.n3113 ),
            .carryout(\transmit_module.n3114 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_13_lut_LC_15_14_3 .C_ON=1'b1;
    defparam \transmit_module.add_13_13_lut_LC_15_14_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_13_lut_LC_15_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_13_lut_LC_15_14_3  (
            .in0(_gnd_net_),
            .in1(N__24310),
            .in2(_gnd_net_),
            .in3(N__16601),
            .lcout(\transmit_module.n121 ),
            .ltout(),
            .carryin(\transmit_module.n3114 ),
            .carryout(\transmit_module.n3115 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_14_lut_LC_15_14_4 .C_ON=1'b1;
    defparam \transmit_module.add_13_14_lut_LC_15_14_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_14_lut_LC_15_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_14_lut_LC_15_14_4  (
            .in0(_gnd_net_),
            .in1(N__23783),
            .in2(_gnd_net_),
            .in3(N__16598),
            .lcout(\transmit_module.n120 ),
            .ltout(),
            .carryin(\transmit_module.n3115 ),
            .carryout(\transmit_module.n3116 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_15_lut_LC_15_14_5 .C_ON=1'b0;
    defparam \transmit_module.add_13_15_lut_LC_15_14_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_15_lut_LC_15_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_15_lut_LC_15_14_5  (
            .in0(_gnd_net_),
            .in1(N__23950),
            .in2(_gnd_net_),
            .in3(N__16595),
            .lcout(\transmit_module.n119 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.ADDR_Y_COMPONENT__i8_LC_15_14_7 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i8_LC_15_14_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i8_LC_15_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i8_LC_15_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17264),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23393),
            .ce(N__20455),
            .sr(N__20352));
    defparam \transmit_module.BRAM_ADDR__i9_LC_15_15_1 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i9_LC_15_15_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i9_LC_15_15_1 .LUT_INIT=16'b0000101100001000;
    LogicCell40 \transmit_module.BRAM_ADDR__i9_LC_15_15_1  (
            .in0(N__19142),
            .in1(N__20821),
            .in2(N__20286),
            .in3(N__19127),
            .lcout(\transmit_module.TX_ADDR_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23227),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i4_LC_15_15_2 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i4_LC_15_15_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i4_LC_15_15_2 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \transmit_module.BRAM_ADDR__i4_LC_15_15_2  (
            .in0(N__20819),
            .in1(N__20171),
            .in2(N__20558),
            .in3(N__18238),
            .lcout(\transmit_module.TX_ADDR_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23227),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i8_LC_15_15_4 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i8_LC_15_15_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i8_LC_15_15_4 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \transmit_module.BRAM_ADDR__i8_LC_15_15_4  (
            .in0(N__20820),
            .in1(N__20172),
            .in2(N__19601),
            .in3(N__19580),
            .lcout(\transmit_module.TX_ADDR_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23227),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i6_3_lut_LC_15_15_6 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i6_3_lut_LC_15_15_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i6_3_lut_LC_15_15_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \transmit_module.mux_12_i6_3_lut_LC_15_15_6  (
            .in0(N__17027),
            .in1(N__20656),
            .in2(_gnd_net_),
            .in3(N__17016),
            .lcout(\transmit_module.n111 ),
            .ltout(\transmit_module.n111_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1614_4_lut_LC_15_15_7 .C_ON=1'b0;
    defparam \transmit_module.i1614_4_lut_LC_15_15_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1614_4_lut_LC_15_15_7 .LUT_INIT=16'b0101000101000000;
    LogicCell40 \transmit_module.i1614_4_lut_LC_15_15_7  (
            .in0(N__20170),
            .in1(N__20818),
            .in2(N__16985),
            .in3(N__16982),
            .lcout(n23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.VGA_VISIBLE_65_LC_15_16_3 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.VGA_VISIBLE_65_LC_15_16_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_VISIBLE_65_LC_15_16_3 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \transmit_module.video_signal_controller.VGA_VISIBLE_65_LC_15_16_3  (
            .in0(N__16742),
            .in1(N__16735),
            .in2(N__16721),
            .in3(N__16685),
            .lcout(\transmit_module.VGA_VISIBLE ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23218),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i11_3_lut_LC_15_16_4 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i11_3_lut_LC_15_16_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i11_3_lut_LC_15_16_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_12_i11_3_lut_LC_15_16_4  (
            .in0(N__20652),
            .in1(N__16673),
            .in2(_gnd_net_),
            .in3(N__16666),
            .lcout(\transmit_module.n106 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1_3_lut_LC_15_16_6 .C_ON=1'b0;
    defparam \transmit_module.i1_3_lut_LC_15_16_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1_3_lut_LC_15_16_6 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \transmit_module.i1_3_lut_LC_15_16_6  (
            .in0(N__20654),
            .in1(N__20179),
            .in2(_gnd_net_),
            .in3(N__20822),
            .lcout(\transmit_module.n2069 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1625_4_lut_LC_15_16_7 .C_ON=1'b0;
    defparam \transmit_module.i1625_4_lut_LC_15_16_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1625_4_lut_LC_15_16_7 .LUT_INIT=16'b1111011111110010;
    LogicCell40 \transmit_module.i1625_4_lut_LC_15_16_7  (
            .in0(N__20823),
            .in1(N__20653),
            .in2(N__20287),
            .in3(N__21602),
            .lcout(\transmit_module.n2057 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i12_LC_15_17_0 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i12_LC_15_17_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i12_LC_15_17_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \transmit_module.BRAM_ADDR__i12_LC_15_17_0  (
            .in0(N__18584),
            .in1(N__20770),
            .in2(_gnd_net_),
            .in3(N__16628),
            .lcout(TX_ADDR_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22937),
            .ce(N__17558),
            .sr(N__20356));
    defparam \transmit_module.BRAM_ADDR__rep_1_i0_LC_15_17_2 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__rep_1_i0_LC_15_17_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__rep_1_i0_LC_15_17_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \transmit_module.BRAM_ADDR__rep_1_i0_LC_15_17_2  (
            .in0(N__18578),
            .in1(N__20772),
            .in2(_gnd_net_),
            .in3(N__17576),
            .lcout(TX_ADDR_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22937),
            .ce(N__17558),
            .sr(N__20356));
    defparam \transmit_module.BRAM_ADDR__i13_LC_15_17_4 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i13_LC_15_17_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i13_LC_15_17_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \transmit_module.BRAM_ADDR__i13_LC_15_17_4  (
            .in0(N__18593),
            .in1(N__20771),
            .in2(_gnd_net_),
            .in3(N__17567),
            .lcout(TX_ADDR_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22937),
            .ce(N__17558),
            .sr(N__20356));
    defparam \transmit_module.mux_14_i9_3_lut_LC_15_18_1 .C_ON=1'b0;
    defparam \transmit_module.mux_14_i9_3_lut_LC_15_18_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_14_i9_3_lut_LC_15_18_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_14_i9_3_lut_LC_15_18_1  (
            .in0(N__21606),
            .in1(N__17272),
            .in2(_gnd_net_),
            .in3(N__17549),
            .lcout(\transmit_module.n139 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_14_i7_3_lut_LC_15_18_5 .C_ON=1'b0;
    defparam \transmit_module.mux_14_i7_3_lut_LC_15_18_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_14_i7_3_lut_LC_15_18_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_14_i7_3_lut_LC_15_18_5  (
            .in0(N__21604),
            .in1(N__19272),
            .in2(_gnd_net_),
            .in3(N__17540),
            .lcout(\transmit_module.n141 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_14_i10_3_lut_LC_15_18_6 .C_ON=1'b0;
    defparam \transmit_module.mux_14_i10_3_lut_LC_15_18_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_14_i10_3_lut_LC_15_18_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_14_i10_3_lut_LC_15_18_6  (
            .in0(N__21603),
            .in1(N__19170),
            .in2(_gnd_net_),
            .in3(N__17531),
            .lcout(\transmit_module.n138 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_14_i8_3_lut_LC_15_18_7 .C_ON=1'b0;
    defparam \transmit_module.mux_14_i8_3_lut_LC_15_18_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_14_i8_3_lut_LC_15_18_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_14_i8_3_lut_LC_15_18_7  (
            .in0(N__21605),
            .in1(N__19334),
            .in2(_gnd_net_),
            .in3(N__17522),
            .lcout(\transmit_module.n140 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1615_4_lut_LC_15_19_0 .C_ON=1'b0;
    defparam \transmit_module.i1615_4_lut_LC_15_19_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1615_4_lut_LC_15_19_0 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \transmit_module.i1615_4_lut_LC_15_19_0  (
            .in0(N__20764),
            .in1(N__19237),
            .in2(N__20187),
            .in3(N__18418),
            .lcout(n22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i9_3_lut_LC_15_19_1 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i9_3_lut_LC_15_19_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i9_3_lut_LC_15_19_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_12_i9_3_lut_LC_15_19_1  (
            .in0(N__20621),
            .in1(N__17285),
            .in2(_gnd_net_),
            .in3(N__17276),
            .lcout(\transmit_module.n108 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1616_4_lut_LC_15_19_6 .C_ON=1'b0;
    defparam \transmit_module.i1616_4_lut_LC_15_19_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1616_4_lut_LC_15_19_6 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \transmit_module.i1616_4_lut_LC_15_19_6  (
            .in0(N__20765),
            .in1(N__19294),
            .in2(N__20188),
            .in3(N__18331),
            .lcout(n21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.ADDR_Y_COMPONENT__i6_LC_15_20_0 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i6_LC_15_20_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i6_LC_15_20_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i6_LC_15_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19277),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22779),
            .ce(N__20479),
            .sr(N__20168));
    defparam \transmit_module.ADDR_Y_COMPONENT__i1_LC_15_20_5 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i1_LC_15_20_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i1_LC_15_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i1_LC_15_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18299),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22779),
            .ce(N__20479),
            .sr(N__20168));
    defparam \transmit_module.mux_14_i5_3_lut_LC_15_21_5 .C_ON=1'b0;
    defparam \transmit_module.mux_14_i5_3_lut_LC_15_21_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_14_i5_3_lut_LC_15_21_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \transmit_module.mux_14_i5_3_lut_LC_15_21_5  (
            .in0(N__18257),
            .in1(N__21618),
            .in2(_gnd_net_),
            .in3(N__20516),
            .lcout(\transmit_module.n143 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_15_26_1.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_15_26_1.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_15_26_1.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_15_26_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.WIRE_OUT_i3_LC_16_5_1 .C_ON=1'b0;
    defparam \tvp_video_buffer.WIRE_OUT_i3_LC_16_5_1 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.WIRE_OUT_i3_LC_16_5_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.WIRE_OUT_i3_LC_16_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17807),
            .lcout(RX_DATA_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24564),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.BUFFER_0__i12_LC_16_5_2 .C_ON=1'b0;
    defparam \tvp_video_buffer.BUFFER_0__i12_LC_16_5_2 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.BUFFER_0__i12_LC_16_5_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.BUFFER_0__i12_LC_16_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17813),
            .lcout(\tvp_video_buffer.BUFFER_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24564),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.BUFFER_0__i13_LC_16_7_3 .C_ON=1'b0;
    defparam \tvp_video_buffer.BUFFER_0__i13_LC_16_7_3 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.BUFFER_0__i13_LC_16_7_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.BUFFER_0__i13_LC_16_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17801),
            .lcout(\tvp_video_buffer.BUFFER_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24570),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.WIRE_OUT_i4_LC_16_7_7 .C_ON=1'b0;
    defparam \tvp_video_buffer.WIRE_OUT_i4_LC_16_7_7 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.WIRE_OUT_i4_LC_16_7_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.WIRE_OUT_i4_LC_16_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17795),
            .lcout(RX_DATA_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24570),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.WIRE_OUT_i5_LC_16_8_6 .C_ON=1'b0;
    defparam \tvp_video_buffer.WIRE_OUT_i5_LC_16_8_6 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.WIRE_OUT_i5_LC_16_8_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.WIRE_OUT_i5_LC_16_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17693),
            .lcout(RX_DATA_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24572),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.WIRE_OUT_i6_LC_16_11_0 .C_ON=1'b0;
    defparam \tvp_video_buffer.WIRE_OUT_i6_LC_16_11_0 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.WIRE_OUT_i6_LC_16_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.WIRE_OUT_i6_LC_16_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18431),
            .lcout(RX_DATA_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24588),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.BUFFER_0__i7_LC_16_11_2 .C_ON=1'b0;
    defparam \tvp_video_buffer.BUFFER_0__i7_LC_16_11_2 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.BUFFER_0__i7_LC_16_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.BUFFER_0__i7_LC_16_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18454),
            .lcout(\tvp_video_buffer.BUFFER_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24588),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.BUFFER_0__i15_LC_16_11_5 .C_ON=1'b0;
    defparam \tvp_video_buffer.BUFFER_0__i15_LC_16_11_5 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.BUFFER_0__i15_LC_16_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.BUFFER_0__i15_LC_16_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18437),
            .lcout(\tvp_video_buffer.BUFFER_1_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24588),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i6_LC_16_12_2 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i6_LC_16_12_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i6_LC_16_12_2 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \transmit_module.BRAM_ADDR__i6_LC_16_12_2  (
            .in0(N__20868),
            .in1(N__19241),
            .in2(N__20353),
            .in3(N__18425),
            .lcout(\transmit_module.TX_ADDR_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23302),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.X_DELTA_PATTERN_i0_LC_16_13_0 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i0_LC_16_13_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i0_LC_16_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i0_LC_16_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21179),
            .lcout(\transmit_module.X_DELTA_PATTERN_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23130),
            .ce(N__21129),
            .sr(N__18382));
    defparam \transmit_module.BRAM_ADDR__i7_LC_16_14_0 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i7_LC_16_14_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i7_LC_16_14_0 .LUT_INIT=16'b0010001100100000;
    LogicCell40 \transmit_module.BRAM_ADDR__i7_LC_16_14_0  (
            .in0(N__19298),
            .in1(N__20237),
            .in2(N__20879),
            .in3(N__18338),
            .lcout(\transmit_module.TX_ADDR_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23392),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_14_i3_3_lut_LC_16_14_4 .C_ON=1'b0;
    defparam \transmit_module.mux_14_i3_3_lut_LC_16_14_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_14_i3_3_lut_LC_16_14_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \transmit_module.mux_14_i3_3_lut_LC_16_14_4  (
            .in0(N__19208),
            .in1(N__21614),
            .in2(_gnd_net_),
            .in3(N__18320),
            .lcout(\transmit_module.n145 ),
            .ltout(\transmit_module.n145_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i2_LC_16_14_5 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i2_LC_16_14_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i2_LC_16_14_5 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \transmit_module.BRAM_ADDR__i2_LC_16_14_5  (
            .in0(N__20236),
            .in1(N__20871),
            .in2(N__18314),
            .in3(N__18889),
            .lcout(\transmit_module.TX_ADDR_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23392),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.Y_DELTA_PATTERN_i16_LC_16_15_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i16_LC_16_15_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i16_LC_16_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i16_LC_16_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18626),
            .lcout(\transmit_module.Y_DELTA_PATTERN_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22700),
            .ce(N__21062),
            .sr(N__20239));
    defparam \transmit_module.Y_DELTA_PATTERN_i17_LC_16_15_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i17_LC_16_15_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i17_LC_16_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i17_LC_16_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18599),
            .lcout(\transmit_module.Y_DELTA_PATTERN_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22700),
            .ce(N__21062),
            .sr(N__20239));
    defparam \transmit_module.Y_DELTA_PATTERN_i19_LC_16_16_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i19_LC_16_16_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i19_LC_16_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i19_LC_16_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18620),
            .lcout(\transmit_module.Y_DELTA_PATTERN_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23194),
            .ce(N__21056),
            .sr(N__20250));
    defparam \transmit_module.Y_DELTA_PATTERN_i18_LC_16_16_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i18_LC_16_16_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i18_LC_16_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i18_LC_16_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18605),
            .lcout(\transmit_module.Y_DELTA_PATTERN_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23194),
            .ce(N__21056),
            .sr(N__20250));
    defparam \transmit_module.ADDR_Y_COMPONENT__i9_LC_16_17_0 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i9_LC_16_17_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i9_LC_16_17_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i9_LC_16_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19178),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22936),
            .ce(N__20472),
            .sr(N__20238));
    defparam \transmit_module.ADDR_Y_COMPONENT__i2_LC_16_17_2 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i2_LC_16_17_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i2_LC_16_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i2_LC_16_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19217),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22936),
            .ce(N__20472),
            .sr(N__20238));
    defparam \transmit_module.ADDR_Y_COMPONENT__i13_LC_16_17_3 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i13_LC_16_17_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i13_LC_16_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i13_LC_16_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23949),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22936),
            .ce(N__20472),
            .sr(N__20238));
    defparam \transmit_module.ADDR_Y_COMPONENT__i12_LC_16_17_4 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i12_LC_16_17_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i12_LC_16_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i12_LC_16_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23733),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22936),
            .ce(N__20472),
            .sr(N__20238));
    defparam \transmit_module.ADDR_Y_COMPONENT__i11_LC_16_17_5 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i11_LC_16_17_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i11_LC_16_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i11_LC_16_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24261),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22936),
            .ce(N__20472),
            .sr(N__20238));
    defparam \transmit_module.ADDR_Y_COMPONENT__i7_LC_16_17_7 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i7_LC_16_17_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i7_LC_16_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i7_LC_16_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19333),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22936),
            .ce(N__20472),
            .sr(N__20238));
    defparam \transmit_module.Y_DELTA_PATTERN_i0_LC_16_18_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i0_LC_16_18_2 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i0_LC_16_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i0_LC_16_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19610),
            .lcout(\transmit_module.Y_DELTA_PATTERN_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23031),
            .ce(N__21061),
            .sr(N__20268));
    defparam \transmit_module.i1617_4_lut_LC_16_19_0 .C_ON=1'b0;
    defparam \transmit_module.i1617_4_lut_LC_16_19_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1617_4_lut_LC_16_19_0 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \transmit_module.i1617_4_lut_LC_16_19_0  (
            .in0(N__20839),
            .in1(N__19591),
            .in2(N__20355),
            .in3(N__19576),
            .lcout(n20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i8_3_lut_LC_16_19_1 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i8_3_lut_LC_16_19_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i8_3_lut_LC_16_19_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_12_i8_3_lut_LC_16_19_1  (
            .in0(N__20611),
            .in1(N__19343),
            .in2(_gnd_net_),
            .in3(N__19332),
            .lcout(\transmit_module.n109 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i7_3_lut_LC_16_19_2 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i7_3_lut_LC_16_19_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i7_3_lut_LC_16_19_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_12_i7_3_lut_LC_16_19_2  (
            .in0(N__20613),
            .in1(N__19283),
            .in2(_gnd_net_),
            .in3(N__19273),
            .lcout(\transmit_module.n110 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i3_3_lut_LC_16_19_3 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i3_3_lut_LC_16_19_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i3_3_lut_LC_16_19_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_12_i3_3_lut_LC_16_19_3  (
            .in0(N__20610),
            .in1(N__19226),
            .in2(_gnd_net_),
            .in3(N__19216),
            .lcout(\transmit_module.n114 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i10_3_lut_LC_16_19_5 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i10_3_lut_LC_16_19_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i10_3_lut_LC_16_19_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_12_i10_3_lut_LC_16_19_5  (
            .in0(N__20612),
            .in1(N__19187),
            .in2(_gnd_net_),
            .in3(N__19177),
            .lcout(\transmit_module.n107 ),
            .ltout(\transmit_module.n107_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1618_4_lut_LC_16_19_6 .C_ON=1'b0;
    defparam \transmit_module.i1618_4_lut_LC_16_19_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1618_4_lut_LC_16_19_6 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \transmit_module.i1618_4_lut_LC_16_19_6  (
            .in0(N__20840),
            .in1(N__20305),
            .in2(N__19130),
            .in3(N__19123),
            .lcout(n19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1611_4_lut_LC_16_31_2 .C_ON=1'b0;
    defparam \transmit_module.i1611_4_lut_LC_16_31_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1611_4_lut_LC_16_31_2 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \transmit_module.i1611_4_lut_LC_16_31_2  (
            .in0(N__20876),
            .in1(N__18890),
            .in2(N__20407),
            .in3(N__18869),
            .lcout(n26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.WIRE_OUT_i2_LC_17_11_7 .C_ON=1'b0;
    defparam \tvp_video_buffer.WIRE_OUT_i2_LC_17_11_7 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.WIRE_OUT_i2_LC_17_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.WIRE_OUT_i2_LC_17_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18641),
            .lcout(RX_DATA_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24580),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.X_DELTA_PATTERN_i15_LC_17_14_5 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i15_LC_17_14_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i15_LC_17_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i15_LC_17_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19672),
            .lcout(\transmit_module.X_DELTA_PATTERN_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23378),
            .ce(N__21119),
            .sr(N__21063));
    defparam \transmit_module.X_DELTA_PATTERN_i9_LC_17_15_0 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i9_LC_17_15_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i9_LC_17_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i9_LC_17_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19658),
            .lcout(\transmit_module.X_DELTA_PATTERN_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23125),
            .ce(N__21111),
            .sr(N__21057));
    defparam \transmit_module.X_DELTA_PATTERN_i10_LC_17_15_2 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i10_LC_17_15_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.X_DELTA_PATTERN_i10_LC_17_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i10_LC_17_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19628),
            .lcout(\transmit_module.X_DELTA_PATTERN_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23125),
            .ce(N__21111),
            .sr(N__21057));
    defparam \transmit_module.X_DELTA_PATTERN_i13_LC_17_15_4 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i13_LC_17_15_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i13_LC_17_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i13_LC_17_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19646),
            .lcout(\transmit_module.X_DELTA_PATTERN_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23125),
            .ce(N__21111),
            .sr(N__21057));
    defparam \transmit_module.X_DELTA_PATTERN_i14_LC_17_15_5 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i14_LC_17_15_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.X_DELTA_PATTERN_i14_LC_17_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i14_LC_17_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19652),
            .lcout(\transmit_module.X_DELTA_PATTERN_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23125),
            .ce(N__21111),
            .sr(N__21057));
    defparam \transmit_module.X_DELTA_PATTERN_i12_LC_17_15_6 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i12_LC_17_15_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.X_DELTA_PATTERN_i12_LC_17_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i12_LC_17_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19640),
            .lcout(\transmit_module.X_DELTA_PATTERN_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23125),
            .ce(N__21111),
            .sr(N__21057));
    defparam \transmit_module.X_DELTA_PATTERN_i11_LC_17_15_7 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i11_LC_17_15_7 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i11_LC_17_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i11_LC_17_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19634),
            .lcout(\transmit_module.X_DELTA_PATTERN_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23125),
            .ce(N__21111),
            .sr(N__21057));
    defparam \transmit_module.X_DELTA_PATTERN_i7_LC_17_16_3 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i7_LC_17_16_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i7_LC_17_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i7_LC_17_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19616),
            .lcout(\transmit_module.X_DELTA_PATTERN_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23391),
            .ce(N__21118),
            .sr(N__21054));
    defparam \transmit_module.X_DELTA_PATTERN_i8_LC_17_16_4 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i8_LC_17_16_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.X_DELTA_PATTERN_i8_LC_17_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i8_LC_17_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19622),
            .lcout(\transmit_module.X_DELTA_PATTERN_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23391),
            .ce(N__21118),
            .sr(N__21054));
    defparam \transmit_module.X_DELTA_PATTERN_i5_LC_17_16_7 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i5_LC_17_16_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.X_DELTA_PATTERN_i5_LC_17_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i5_LC_17_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21137),
            .lcout(\transmit_module.X_DELTA_PATTERN_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23391),
            .ce(N__21118),
            .sr(N__21054));
    defparam \transmit_module.i2_3_lut_LC_17_17_1 .C_ON=1'b0;
    defparam \transmit_module.i2_3_lut_LC_17_17_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i2_3_lut_LC_17_17_1 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \transmit_module.i2_3_lut_LC_17_17_1  (
            .in0(N__20229),
            .in1(N__20841),
            .in2(_gnd_net_),
            .in3(N__21622),
            .lcout(\transmit_module.n2115 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2176_3_lut_LC_17_18_0 .C_ON=1'b0;
    defparam \line_buffer.i2176_3_lut_LC_17_18_0 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2176_3_lut_LC_17_18_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \line_buffer.i2176_3_lut_LC_17_18_0  (
            .in0(N__20687),
            .in1(N__20669),
            .in2(_gnd_net_),
            .in3(N__24335),
            .lcout(\line_buffer.n3519 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i5_3_lut_LC_17_19_5 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i5_3_lut_LC_17_19_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i5_3_lut_LC_17_19_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \transmit_module.mux_12_i5_3_lut_LC_17_19_5  (
            .in0(N__20524),
            .in1(N__20620),
            .in2(_gnd_net_),
            .in3(N__20486),
            .lcout(\transmit_module.n112 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.ADDR_Y_COMPONENT__i4_LC_17_20_7 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i4_LC_17_20_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i4_LC_17_20_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i4_LC_17_20_7  (
            .in0(N__20528),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23262),
            .ce(N__20480),
            .sr(N__20169));
    defparam \line_buffer.i2157_3_lut_LC_17_21_3 .C_ON=1'b0;
    defparam \line_buffer.i2157_3_lut_LC_17_21_3 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2157_3_lut_LC_17_21_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \line_buffer.i2157_3_lut_LC_17_21_3  (
            .in0(N__24373),
            .in1(N__19826),
            .in2(_gnd_net_),
            .in3(N__19811),
            .lcout(),
            .ltout(\line_buffer.n3500_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_2210_LC_17_21_4 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_2210_LC_17_21_4 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_2210_LC_17_21_4 .LUT_INIT=16'b1110101001100010;
    LogicCell40 \line_buffer.TX_ADDR_12__bdd_4_lut_2210_LC_17_21_4  (
            .in0(N__23827),
            .in1(N__24010),
            .in2(N__19796),
            .in3(N__19793),
            .lcout(),
            .ltout(\line_buffer.n3537_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i6_LC_17_21_5 .C_ON=1'b0;
    defparam \line_buffer.dout_i6_LC_17_21_5 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i6_LC_17_21_5 .LUT_INIT=16'b1111000011001010;
    LogicCell40 \line_buffer.dout_i6_LC_17_21_5  (
            .in0(N__21239),
            .in1(N__21461),
            .in2(N__19781),
            .in3(N__24011),
            .lcout(TX_DATA_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23015),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2154_3_lut_LC_17_22_0 .C_ON=1'b0;
    defparam \line_buffer.i2154_3_lut_LC_17_22_0 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2154_3_lut_LC_17_22_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \line_buffer.i2154_3_lut_LC_17_22_0  (
            .in0(N__21272),
            .in1(N__21257),
            .in2(_gnd_net_),
            .in3(N__24385),
            .lcout(\line_buffer.n3497 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2178_3_lut_LC_18_11_2 .C_ON=1'b0;
    defparam \line_buffer.i2178_3_lut_LC_18_11_2 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2178_3_lut_LC_18_11_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \line_buffer.i2178_3_lut_LC_18_11_2  (
            .in0(N__24384),
            .in1(N__21233),
            .in2(_gnd_net_),
            .in3(N__21215),
            .lcout(\line_buffer.n3521 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2182_3_lut_LC_18_13_2 .C_ON=1'b0;
    defparam \line_buffer.i2182_3_lut_LC_18_13_2 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2182_3_lut_LC_18_13_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \line_buffer.i2182_3_lut_LC_18_13_2  (
            .in0(N__21206),
            .in1(N__21188),
            .in2(_gnd_net_),
            .in3(N__24357),
            .lcout(\line_buffer.n3525 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.X_DELTA_PATTERN_i1_LC_18_14_0 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i1_LC_18_14_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.X_DELTA_PATTERN_i1_LC_18_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i1_LC_18_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21167),
            .lcout(\transmit_module.X_DELTA_PATTERN_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23389),
            .ce(N__21131),
            .sr(N__21064));
    defparam \transmit_module.X_DELTA_PATTERN_i2_LC_18_14_1 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i2_LC_18_14_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i2_LC_18_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i2_LC_18_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21161),
            .lcout(\transmit_module.X_DELTA_PATTERN_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23389),
            .ce(N__21131),
            .sr(N__21064));
    defparam \transmit_module.X_DELTA_PATTERN_i3_LC_18_14_2 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i3_LC_18_14_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.X_DELTA_PATTERN_i3_LC_18_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i3_LC_18_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21149),
            .lcout(\transmit_module.X_DELTA_PATTERN_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23389),
            .ce(N__21131),
            .sr(N__21064));
    defparam \transmit_module.X_DELTA_PATTERN_i4_LC_18_15_6 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i4_LC_18_15_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i4_LC_18_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i4_LC_18_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21155),
            .lcout(\transmit_module.X_DELTA_PATTERN_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23147),
            .ce(N__21117),
            .sr(N__21065));
    defparam \transmit_module.X_DELTA_PATTERN_i6_LC_18_16_6 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i6_LC_18_16_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i6_LC_18_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i6_LC_18_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21143),
            .lcout(\transmit_module.X_DELTA_PATTERN_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23464),
            .ce(N__21130),
            .sr(N__21055));
    defparam \line_buffer.i2181_3_lut_LC_18_17_0 .C_ON=1'b0;
    defparam \line_buffer.i2181_3_lut_LC_18_17_0 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2181_3_lut_LC_18_17_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \line_buffer.i2181_3_lut_LC_18_17_0  (
            .in0(N__20909),
            .in1(N__20894),
            .in2(_gnd_net_),
            .in3(N__24367),
            .lcout(),
            .ltout(\line_buffer.n3524_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i5_LC_18_17_1 .C_ON=1'b0;
    defparam \line_buffer.dout_i5_LC_18_17_1 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i5_LC_18_17_1 .LUT_INIT=16'b1110111001010000;
    LogicCell40 \line_buffer.dout_i5_LC_18_17_1  (
            .in0(N__23974),
            .in1(N__21530),
            .in2(N__21521),
            .in3(N__21725),
            .lcout(TX_DATA_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23433),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_2215_LC_18_19_1 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_2215_LC_18_19_1 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_2215_LC_18_19_1 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \line_buffer.TX_ADDR_12__bdd_4_lut_2215_LC_18_19_1  (
            .in0(N__23826),
            .in1(N__22343),
            .in2(N__24009),
            .in3(N__21518),
            .lcout(),
            .ltout(\line_buffer.n3555_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i1_LC_18_19_2 .C_ON=1'b0;
    defparam \line_buffer.dout_i1_LC_18_19_2 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i1_LC_18_19_2 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \line_buffer.dout_i1_LC_18_19_2  (
            .in0(N__23997),
            .in1(N__24161),
            .in2(N__21509),
            .in3(N__21506),
            .lcout(TX_DATA_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22969),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2155_3_lut_LC_18_20_0 .C_ON=1'b0;
    defparam \line_buffer.i2155_3_lut_LC_18_20_0 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2155_3_lut_LC_18_20_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \line_buffer.i2155_3_lut_LC_18_20_0  (
            .in0(N__24341),
            .in1(N__21500),
            .in2(_gnd_net_),
            .in3(N__21482),
            .lcout(\line_buffer.n3498 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2250_LC_18_20_2 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2250_LC_18_20_2 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2250_LC_18_20_2 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_2250_LC_18_20_2  (
            .in0(N__24340),
            .in1(N__21455),
            .in2(N__23846),
            .in3(N__21446),
            .lcout(\line_buffer.n3597 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.VGA_R__i1_LC_18_21_0 .C_ON=1'b0;
    defparam \transmit_module.VGA_R__i1_LC_18_21_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.VGA_R__i1_LC_18_21_0 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \transmit_module.VGA_R__i1_LC_18_21_0  (
            .in0(_gnd_net_),
            .in1(N__21629),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n1814),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23019),
            .ce(),
            .sr(N__24784));
    defparam \transmit_module.VGA_R__i2_LC_18_22_3 .C_ON=1'b0;
    defparam \transmit_module.VGA_R__i2_LC_18_22_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.VGA_R__i2_LC_18_22_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.VGA_R__i2_LC_18_22_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21386),
            .lcout(n1813),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23061),
            .ce(),
            .sr(N__24796));
    defparam \transmit_module.VGA_R__i6_LC_18_23_6 .C_ON=1'b0;
    defparam \transmit_module.VGA_R__i6_LC_18_23_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.VGA_R__i6_LC_18_23_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.VGA_R__i6_LC_18_23_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21326),
            .lcout(n1809),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22772),
            .ce(),
            .sr(N__24798));
    defparam \transmit_module.VGA_R__i7_LC_18_24_1 .C_ON=1'b0;
    defparam \transmit_module.VGA_R__i7_LC_18_24_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.VGA_R__i7_LC_18_24_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.VGA_R__i7_LC_18_24_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21878),
            .lcout(n1808),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22911),
            .ce(),
            .sr(N__24797));
    defparam \line_buffer.i2145_3_lut_LC_19_9_3 .C_ON=1'b0;
    defparam \line_buffer.i2145_3_lut_LC_19_9_3 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2145_3_lut_LC_19_9_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \line_buffer.i2145_3_lut_LC_19_9_3  (
            .in0(N__24378),
            .in1(N__21815),
            .in2(_gnd_net_),
            .in3(N__21800),
            .lcout(\line_buffer.n3488 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i7_LC_19_15_5 .C_ON=1'b0;
    defparam \line_buffer.dout_i7_LC_19_15_5 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i7_LC_19_15_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \line_buffer.dout_i7_LC_19_15_5  (
            .in0(N__23998),
            .in1(N__21785),
            .in2(_gnd_net_),
            .in3(N__22037),
            .lcout(TX_DATA_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23129),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2146_3_lut_LC_19_16_1 .C_ON=1'b0;
    defparam \line_buffer.i2146_3_lut_LC_19_16_1 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2146_3_lut_LC_19_16_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \line_buffer.i2146_3_lut_LC_19_16_1  (
            .in0(N__24369),
            .in1(N__21776),
            .in2(_gnd_net_),
            .in3(N__21761),
            .lcout(\line_buffer.n3489 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_2220_LC_19_17_3 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_2220_LC_19_17_3 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_2220_LC_19_17_3 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \line_buffer.TX_ADDR_12__bdd_4_lut_2220_LC_19_17_3  (
            .in0(N__23819),
            .in1(N__21740),
            .in2(N__24008),
            .in3(N__21734),
            .lcout(\line_buffer.n3561 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2230_LC_19_17_4 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2230_LC_19_17_4 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2230_LC_19_17_4 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_2230_LC_19_17_4  (
            .in0(N__24290),
            .in1(N__21719),
            .in2(N__23842),
            .in3(N__21704),
            .lcout(\line_buffer.n3573 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n3597_bdd_4_lut_LC_19_20_0 .C_ON=1'b0;
    defparam \line_buffer.n3597_bdd_4_lut_LC_19_20_0 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3597_bdd_4_lut_LC_19_20_0 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \line_buffer.n3597_bdd_4_lut_LC_19_20_0  (
            .in0(N__21683),
            .in1(N__23833),
            .in2(N__21659),
            .in3(N__21638),
            .lcout(),
            .ltout(\line_buffer.n3600_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i0_LC_19_20_1 .C_ON=1'b0;
    defparam \line_buffer.dout_i0_LC_19_20_1 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i0_LC_19_20_1 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \line_buffer.dout_i0_LC_19_20_1  (
            .in0(_gnd_net_),
            .in1(N__23996),
            .in2(N__21632),
            .in3(N__22286),
            .lcout(TX_DATA_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23263),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1118_1_lut_LC_19_21_1 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1118_1_lut_LC_19_21_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1118_1_lut_LC_19_21_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \transmit_module.video_signal_controller.i1118_1_lut_LC_19_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21623),
            .lcout(\transmit_module.n2367 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.VGA_R__i8_LC_19_22_6 .C_ON=1'b0;
    defparam \transmit_module.VGA_R__i8_LC_19_22_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.VGA_R__i8_LC_19_22_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.VGA_R__i8_LC_19_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22220),
            .lcout(ADV_B_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23123),
            .ce(),
            .sr(N__24792));
    defparam \tvp_video_buffer.WIRE_OUT_i7_LC_20_4_5 .C_ON=1'b0;
    defparam \tvp_video_buffer.WIRE_OUT_i7_LC_20_4_5 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.WIRE_OUT_i7_LC_20_4_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.WIRE_OUT_i7_LC_20_4_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24728),
            .lcout(RX_DATA_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24567),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n3585_bdd_4_lut_LC_20_15_2 .C_ON=1'b0;
    defparam \line_buffer.n3585_bdd_4_lut_LC_20_15_2 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3585_bdd_4_lut_LC_20_15_2 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \line_buffer.n3585_bdd_4_lut_LC_20_15_2  (
            .in0(N__22073),
            .in1(N__23840),
            .in2(N__22055),
            .in3(N__24056),
            .lcout(\line_buffer.n3588 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2225_LC_20_15_3 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2225_LC_20_15_3 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2225_LC_20_15_3 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_2225_LC_20_15_3  (
            .in0(N__24337),
            .in1(N__22031),
            .in2(N__23849),
            .in3(N__22019),
            .lcout(\line_buffer.n3549 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n3549_bdd_4_lut_LC_20_17_1 .C_ON=1'b0;
    defparam \line_buffer.n3549_bdd_4_lut_LC_20_17_1 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3549_bdd_4_lut_LC_20_17_1 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \line_buffer.n3549_bdd_4_lut_LC_20_17_1  (
            .in0(N__22004),
            .in1(N__23816),
            .in2(N__21989),
            .in3(N__21965),
            .lcout(),
            .ltout(\line_buffer.n3552_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i2_LC_20_17_2 .C_ON=1'b0;
    defparam \line_buffer.dout_i2_LC_20_17_2 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i2_LC_20_17_2 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \line_buffer.dout_i2_LC_20_17_2  (
            .in0(_gnd_net_),
            .in1(N__23986),
            .in2(N__21956),
            .in3(N__22469),
            .lcout(TX_DATA_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23390),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n3573_bdd_4_lut_LC_20_17_3 .C_ON=1'b0;
    defparam \line_buffer.n3573_bdd_4_lut_LC_20_17_3 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3573_bdd_4_lut_LC_20_17_3 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \line_buffer.n3573_bdd_4_lut_LC_20_17_3  (
            .in0(N__21953),
            .in1(N__23817),
            .in2(N__21938),
            .in3(N__21917),
            .lcout(\line_buffer.n3576 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_LC_20_17_6 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_LC_20_17_6 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_LC_20_17_6 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_LC_20_17_6  (
            .in0(N__24344),
            .in1(N__21911),
            .in2(N__23844),
            .in3(N__21896),
            .lcout(),
            .ltout(\line_buffer.n3603_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n3603_bdd_4_lut_LC_20_17_7 .C_ON=1'b0;
    defparam \line_buffer.n3603_bdd_4_lut_LC_20_17_7 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3603_bdd_4_lut_LC_20_17_7 .LUT_INIT=16'b1111000011001010;
    LogicCell40 \line_buffer.n3603_bdd_4_lut_LC_20_17_7  (
            .in0(N__22502),
            .in1(N__22487),
            .in2(N__22472),
            .in3(N__23818),
            .lcout(\line_buffer.n3606 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n3543_bdd_4_lut_LC_20_18_3 .C_ON=1'b0;
    defparam \line_buffer.n3543_bdd_4_lut_LC_20_18_3 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3543_bdd_4_lut_LC_20_18_3 .LUT_INIT=16'b1110111001010000;
    LogicCell40 \line_buffer.n3543_bdd_4_lut_LC_20_18_3  (
            .in0(N__23831),
            .in1(N__22463),
            .in2(N__22448),
            .in3(N__23657),
            .lcout(),
            .ltout(\line_buffer.n3546_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i4_LC_20_18_4 .C_ON=1'b0;
    defparam \line_buffer.dout_i4_LC_20_18_4 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i4_LC_20_18_4 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \line_buffer.dout_i4_LC_20_18_4  (
            .in0(_gnd_net_),
            .in1(N__24016),
            .in2(N__22430),
            .in3(N__22427),
            .lcout(TX_DATA_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23183),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2235_LC_20_18_7 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2235_LC_20_18_7 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2235_LC_20_18_7 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_2235_LC_20_18_7  (
            .in0(N__24368),
            .in1(N__22421),
            .in2(N__23847),
            .in3(N__22409),
            .lcout(\line_buffer.n3579 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2139_3_lut_LC_20_19_0 .C_ON=1'b0;
    defparam \line_buffer.i2139_3_lut_LC_20_19_0 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2139_3_lut_LC_20_19_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \line_buffer.i2139_3_lut_LC_20_19_0  (
            .in0(N__22400),
            .in1(N__22385),
            .in2(_gnd_net_),
            .in3(N__24380),
            .lcout(\line_buffer.n3482 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2179_3_lut_LC_20_19_3 .C_ON=1'b0;
    defparam \line_buffer.i2179_3_lut_LC_20_19_3 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2179_3_lut_LC_20_19_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \line_buffer.i2179_3_lut_LC_20_19_3  (
            .in0(N__24379),
            .in1(N__22370),
            .in2(_gnd_net_),
            .in3(N__22358),
            .lcout(\line_buffer.n3522 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n3579_bdd_4_lut_LC_20_20_1 .C_ON=1'b0;
    defparam \line_buffer.n3579_bdd_4_lut_LC_20_20_1 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3579_bdd_4_lut_LC_20_20_1 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \line_buffer.n3579_bdd_4_lut_LC_20_20_1  (
            .in0(N__22334),
            .in1(N__23832),
            .in2(N__22319),
            .in3(N__22295),
            .lcout(\line_buffer.n3582 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.VGA_R__i3_LC_20_21_4 .C_ON=1'b0;
    defparam \transmit_module.VGA_R__i3_LC_20_21_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.VGA_R__i3_LC_20_21_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.VGA_R__i3_LC_20_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22280),
            .lcout(n1812),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22932),
            .ce(),
            .sr(N__24785));
    defparam \transmit_module.VGA_R__i5_LC_20_24_1 .C_ON=1'b0;
    defparam \transmit_module.VGA_R__i5_LC_20_24_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.VGA_R__i5_LC_20_24_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.VGA_R__i5_LC_20_24_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24152),
            .lcout(n1810),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23092),
            .ce(),
            .sr(N__24799));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2240_LC_21_15_7 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2240_LC_21_15_7 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2240_LC_21_15_7 .LUT_INIT=16'b1110101001001010;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_2240_LC_21_15_7  (
            .in0(N__24336),
            .in1(N__24086),
            .in2(N__23848),
            .in3(N__24071),
            .lcout(\line_buffer.n3585 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2140_3_lut_LC_21_16_1 .C_ON=1'b0;
    defparam \line_buffer.i2140_3_lut_LC_21_16_1 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2140_3_lut_LC_21_16_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \line_buffer.i2140_3_lut_LC_21_16_1  (
            .in0(N__24377),
            .in1(N__24050),
            .in2(_gnd_net_),
            .in3(N__24032),
            .lcout(\line_buffer.n3483 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_LC_21_16_3 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_LC_21_16_3 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_LC_21_16_3 .LUT_INIT=16'b1110101001001010;
    LogicCell40 \line_buffer.TX_ADDR_12__bdd_4_lut_LC_21_16_3  (
            .in0(N__23845),
            .in1(N__24689),
            .in2(N__24017),
            .in3(N__23624),
            .lcout(),
            .ltout(\line_buffer.n3567_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i3_LC_21_16_4 .C_ON=1'b0;
    defparam \line_buffer.dout_i3_LC_21_16_4 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i3_LC_21_16_4 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \line_buffer.dout_i3_LC_21_16_4  (
            .in0(N__24015),
            .in1(N__23888),
            .in2(N__23879),
            .in3(N__23876),
            .lcout(TX_DATA_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23499),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2205_LC_21_17_1 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2205_LC_21_17_1 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2205_LC_21_17_1 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_2205_LC_21_17_1  (
            .in0(N__24342),
            .in1(N__23870),
            .in2(N__23843),
            .in3(N__23669),
            .lcout(\line_buffer.n3543 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2137_3_lut_LC_21_17_7 .C_ON=1'b0;
    defparam \line_buffer.i2137_3_lut_LC_21_17_7 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2137_3_lut_LC_21_17_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \line_buffer.i2137_3_lut_LC_21_17_7  (
            .in0(N__24343),
            .in1(N__23651),
            .in2(_gnd_net_),
            .in3(N__23636),
            .lcout(\line_buffer.n3480 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.VGA_R__i4_LC_21_21_4 .C_ON=1'b0;
    defparam \transmit_module.VGA_R__i4_LC_21_21_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.VGA_R__i4_LC_21_21_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.VGA_R__i4_LC_21_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23618),
            .lcout(n1811),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23184),
            .ce(),
            .sr(N__24803));
    defparam \tvp_video_buffer.BUFFER_0__i16_LC_22_4_7 .C_ON=1'b0;
    defparam \tvp_video_buffer.BUFFER_0__i16_LC_22_4_7 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.BUFFER_0__i16_LC_22_4_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.BUFFER_0__i16_LC_22_4_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24647),
            .lcout(\tvp_video_buffer.BUFFER_1_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24573),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2136_3_lut_LC_22_15_0 .C_ON=1'b0;
    defparam \line_buffer.i2136_3_lut_LC_22_15_0 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2136_3_lut_LC_22_15_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \line_buffer.i2136_3_lut_LC_22_15_0  (
            .in0(N__24719),
            .in1(N__24338),
            .in2(_gnd_net_),
            .in3(N__24704),
            .lcout(\line_buffer.n3479 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.BUFFER_0__i8_LC_23_4_6 .C_ON=1'b0;
    defparam \tvp_video_buffer.BUFFER_0__i8_LC_23_4_6 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.BUFFER_0__i8_LC_23_4_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \tvp_video_buffer.BUFFER_0__i8_LC_23_4_6  (
            .in0(N__24664),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\tvp_video_buffer.BUFFER_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24578),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2175_3_lut_LC_24_19_2 .C_ON=1'b0;
    defparam \line_buffer.i2175_3_lut_LC_24_19_2 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2175_3_lut_LC_24_19_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \line_buffer.i2175_3_lut_LC_24_19_2  (
            .in0(N__24413),
            .in1(N__24401),
            .in2(_gnd_net_),
            .in3(N__24386),
            .lcout(\line_buffer.n3518 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // main
