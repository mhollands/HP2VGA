// Verilog netlist produced by program LSE :  version Diamond Version 0.0.0
// Netlist written on Sat Sep 15 01:57:52 2018
//
// Verilog Description of module main
//

module main (DEBUG, TVP_CLK, TVP_HSYNC, TVP_VSYNC, TVP_VIDEO, LED, 
            ADV_HSYNC, ADV_VSYNC, ADV_R, ADV_G, ADV_B, ADV_CLK, 
            ADV_SYNC_N, ADV_BLANK_N) /* synthesis syn_module_defined=1 */ ;   // ../main.v(1[8:12])
    output [7:0]DEBUG;   // ../main.v(2[19:24])
    input TVP_CLK;   // ../main.v(3[13:20])
    input TVP_HSYNC;   // ../main.v(4[13:22])
    input TVP_VSYNC;   // ../main.v(5[13:22])
    input [9:0]TVP_VIDEO;   // ../main.v(6[19:28])
    output LED;   // ../main.v(7[14:17])
    output ADV_HSYNC;   // ../main.v(8[14:23])
    output ADV_VSYNC;   // ../main.v(9[14:23])
    output [7:0]ADV_R;   // ../main.v(10[19:24])
    output [7:0]ADV_G;   // ../main.v(11[19:24])
    output [7:0]ADV_B;   // ../main.v(12[19:24])
    output ADV_CLK;   // ../main.v(13[14:21])
    output ADV_SYNC_N;   // ../main.v(14[14:24])
    output ADV_BLANK_N;   // ../main.v(15[14:25])
    
    wire TVP_CLK_c /* synthesis SET_AS_NETWORK=TVP_CLK_c, is_clock=1 */ ;   // ../main.v(3[13:20])
    wire ADV_CLK_c /* synthesis SET_AS_NETWORK=ADV_CLK_c, is_clock=1 */ ;   // ../main.v(13[14:21])
    
    wire GND_net, VCC_net, DEBUG_c_6, DEBUG_c_5, DEBUG_c_3, DEBUG_c_2, 
        TVP_HSYNC_c, TVP_VSYNC_c, TVP_VIDEO_c_9, TVP_VIDEO_c_8, TVP_VIDEO_c_7, 
        TVP_VIDEO_c_6, TVP_VIDEO_c_5, TVP_VIDEO_c_4, TVP_VIDEO_c_3, 
        TVP_VIDEO_c_2, LED_c, ADV_HSYNC_c, ADV_VSYNC_c, ADV_B_c, n1844, 
        n1845, n1846, n1847, n1848, n1849, n1850;
    wire [13:0]RX_ADDR;   // ../main.v(28[14:21])
    wire [13:0]TX_ADDR;   // ../main.v(47[14:21])
    wire [7:0]TX_DATA;   // ../main.v(48[13:20])
    
    wire n2057, old_HS, n21, n20, n19, n22, n18, n28, n26, 
        n27, n2404, n25, n24, n23, n3860, n3852;
    
    VCC i2 (.Y(VCC_net));
    RX receive_module (.\RX_ADDR[6] (RX_ADDR[6]), .GND_net(GND_net), .\RX_ADDR[5] (RX_ADDR[5]), 
       .\RX_ADDR[11] (RX_ADDR[11]), .\RX_ADDR[2] (RX_ADDR[2]), .DEBUG_c_5(DEBUG_c_5), 
       .TVP_VSYNC_c(TVP_VSYNC_c), .\RX_ADDR[4] (RX_ADDR[4]), .\RX_ADDR[3] (RX_ADDR[3]), 
       .\RX_ADDR[0] (RX_ADDR[0]), .\RX_ADDR[10] (RX_ADDR[10]), .VCC_net(VCC_net), 
       .\RX_ADDR[1] (RX_ADDR[1]), .\RX_ADDR[9] (RX_ADDR[9]), .\RX_ADDR[12] (RX_ADDR[12]), 
       .TVP_CLK_c(TVP_CLK_c), .\RX_ADDR[8] (RX_ADDR[8]), .DEBUG_c_3(DEBUG_c_3), 
       .\RX_ADDR[7] (RX_ADDR[7]), .TVP_HSYNC_c(TVP_HSYNC_c), .old_HS(old_HS), 
       .DEBUG_c_6(DEBUG_c_6), .n3860(n3860), .n2057(n2057), .LED_c(LED_c)) /* synthesis syn_module_defined=1 */ ;   // ../main.v(33[5] 44[29])
    TX transmit_module (.GND_net(GND_net), .ADV_HSYNC_c(ADV_HSYNC_c), .ADV_CLK_c(ADV_CLK_c), 
       .ADV_VSYNC_c(ADV_VSYNC_c), .n23(n23), .DEBUG_c_2(DEBUG_c_2), .\TX_ADDR[12] (TX_ADDR[12]), 
       .n22(n22), .n18(n18), .n19(n19), .n20(n20), .n21(n21), .n24(n24), 
       .n25(n25), .n26(n26), .n27(n27), .\TX_ADDR[11] (TX_ADDR[11]), 
       .n3852(n3852), .n28(n28), .VCC_net(VCC_net), .DEBUG_c_6(DEBUG_c_6), 
       .n2404(n2404)) /* synthesis syn_module_defined=1 */ ;   // ../main.v(51[5] 63[34])
    SB_IO ADV_R_pad_7 (.PACKAGE_PIN(ADV_R[7]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(ADV_B_c));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_R_pad_7.PIN_TYPE = 6'b011001;
    defparam ADV_R_pad_7.PULLUP = 1'b0;
    defparam ADV_R_pad_7.NEG_TRIGGER = 1'b0;
    defparam ADV_R_pad_7.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_pad_4 (.PACKAGE_PIN(DEBUG[4]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n3852));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_pad_4.PIN_TYPE = 6'b011001;
    defparam DEBUG_pad_4.PULLUP = 1'b0;
    defparam DEBUG_pad_4.NEG_TRIGGER = 1'b0;
    defparam DEBUG_pad_4.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_pad_2 (.PACKAGE_PIN(DEBUG[2]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(DEBUG_c_2));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_pad_2.PIN_TYPE = 6'b011001;
    defparam DEBUG_pad_2.PULLUP = 1'b0;
    defparam DEBUG_pad_2.NEG_TRIGGER = 1'b0;
    defparam DEBUG_pad_2.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_pad_5 (.PACKAGE_PIN(DEBUG[5]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(DEBUG_c_5));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_pad_5.PIN_TYPE = 6'b011001;
    defparam DEBUG_pad_5.PULLUP = 1'b0;
    defparam DEBUG_pad_5.NEG_TRIGGER = 1'b0;
    defparam DEBUG_pad_5.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_HSYNC_pad (.PACKAGE_PIN(ADV_HSYNC), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(ADV_HSYNC_c));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_HSYNC_pad.PIN_TYPE = 6'b011001;
    defparam ADV_HSYNC_pad.PULLUP = 1'b0;
    defparam ADV_HSYNC_pad.NEG_TRIGGER = 1'b0;
    defparam ADV_HSYNC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_R_pad_6 (.PACKAGE_PIN(ADV_R[6]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1844));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_R_pad_6.PIN_TYPE = 6'b011001;
    defparam ADV_R_pad_6.PULLUP = 1'b0;
    defparam ADV_R_pad_6.NEG_TRIGGER = 1'b0;
    defparam ADV_R_pad_6.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_pad_3 (.PACKAGE_PIN(DEBUG[3]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(DEBUG_c_3));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_pad_3.PIN_TYPE = 6'b011001;
    defparam DEBUG_pad_3.PULLUP = 1'b0;
    defparam DEBUG_pad_3.NEG_TRIGGER = 1'b0;
    defparam DEBUG_pad_3.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_pad_6 (.PACKAGE_PIN(DEBUG[6]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(DEBUG_c_6));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_pad_6.PIN_TYPE = 6'b011001;
    defparam DEBUG_pad_6.PULLUP = 1'b0;
    defparam DEBUG_pad_6.NEG_TRIGGER = 1'b0;
    defparam DEBUG_pad_6.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_pad_7 (.PACKAGE_PIN(DEBUG[7]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(GND_net));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_pad_7.PIN_TYPE = 6'b011001;
    defparam DEBUG_pad_7.PULLUP = 1'b0;
    defparam DEBUG_pad_7.NEG_TRIGGER = 1'b0;
    defparam DEBUG_pad_7.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_VSYNC_pad (.PACKAGE_PIN(ADV_VSYNC), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(ADV_VSYNC_c));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_VSYNC_pad.PIN_TYPE = 6'b011001;
    defparam ADV_VSYNC_pad.PULLUP = 1'b0;
    defparam ADV_VSYNC_pad.NEG_TRIGGER = 1'b0;
    defparam ADV_VSYNC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_pad_1 (.PACKAGE_PIN(DEBUG[1]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(GND_net));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_pad_1.PIN_TYPE = 6'b011001;
    defparam DEBUG_pad_1.PULLUP = 1'b0;
    defparam DEBUG_pad_1.NEG_TRIGGER = 1'b0;
    defparam DEBUG_pad_1.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_R_pad_5 (.PACKAGE_PIN(ADV_R[5]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1845));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_R_pad_5.PIN_TYPE = 6'b011001;
    defparam ADV_R_pad_5.PULLUP = 1'b0;
    defparam ADV_R_pad_5.NEG_TRIGGER = 1'b0;
    defparam ADV_R_pad_5.IO_STANDARD = "SB_LVCMOS";
    SB_IO LED_pad (.PACKAGE_PIN(LED), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(LED_c));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam LED_pad.PIN_TYPE = 6'b011001;
    defparam LED_pad.PULLUP = 1'b0;
    defparam LED_pad.NEG_TRIGGER = 1'b0;
    defparam LED_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_R_pad_4 (.PACKAGE_PIN(ADV_R[4]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1846));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_R_pad_4.PIN_TYPE = 6'b011001;
    defparam ADV_R_pad_4.PULLUP = 1'b0;
    defparam ADV_R_pad_4.NEG_TRIGGER = 1'b0;
    defparam ADV_R_pad_4.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_R_pad_3 (.PACKAGE_PIN(ADV_R[3]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1847));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_R_pad_3.PIN_TYPE = 6'b011001;
    defparam ADV_R_pad_3.PULLUP = 1'b0;
    defparam ADV_R_pad_3.NEG_TRIGGER = 1'b0;
    defparam ADV_R_pad_3.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_R_pad_2 (.PACKAGE_PIN(ADV_R[2]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1848));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_R_pad_2.PIN_TYPE = 6'b011001;
    defparam ADV_R_pad_2.PULLUP = 1'b0;
    defparam ADV_R_pad_2.NEG_TRIGGER = 1'b0;
    defparam ADV_R_pad_2.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_R_pad_1 (.PACKAGE_PIN(ADV_R[1]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1849));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_R_pad_1.PIN_TYPE = 6'b011001;
    defparam ADV_R_pad_1.PULLUP = 1'b0;
    defparam ADV_R_pad_1.NEG_TRIGGER = 1'b0;
    defparam ADV_R_pad_1.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_R_pad_0 (.PACKAGE_PIN(ADV_R[0]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1850));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_R_pad_0.PIN_TYPE = 6'b011001;
    defparam ADV_R_pad_0.PULLUP = 1'b0;
    defparam ADV_R_pad_0.NEG_TRIGGER = 1'b0;
    defparam ADV_R_pad_0.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_G_pad_7 (.PACKAGE_PIN(ADV_G[7]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(ADV_B_c));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_G_pad_7.PIN_TYPE = 6'b011001;
    defparam ADV_G_pad_7.PULLUP = 1'b0;
    defparam ADV_G_pad_7.NEG_TRIGGER = 1'b0;
    defparam ADV_G_pad_7.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_G_pad_6 (.PACKAGE_PIN(ADV_G[6]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1844));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_G_pad_6.PIN_TYPE = 6'b011001;
    defparam ADV_G_pad_6.PULLUP = 1'b0;
    defparam ADV_G_pad_6.NEG_TRIGGER = 1'b0;
    defparam ADV_G_pad_6.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_G_pad_5 (.PACKAGE_PIN(ADV_G[5]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1845));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_G_pad_5.PIN_TYPE = 6'b011001;
    defparam ADV_G_pad_5.PULLUP = 1'b0;
    defparam ADV_G_pad_5.NEG_TRIGGER = 1'b0;
    defparam ADV_G_pad_5.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_G_pad_4 (.PACKAGE_PIN(ADV_G[4]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1846));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_G_pad_4.PIN_TYPE = 6'b011001;
    defparam ADV_G_pad_4.PULLUP = 1'b0;
    defparam ADV_G_pad_4.NEG_TRIGGER = 1'b0;
    defparam ADV_G_pad_4.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_G_pad_3 (.PACKAGE_PIN(ADV_G[3]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1847));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_G_pad_3.PIN_TYPE = 6'b011001;
    defparam ADV_G_pad_3.PULLUP = 1'b0;
    defparam ADV_G_pad_3.NEG_TRIGGER = 1'b0;
    defparam ADV_G_pad_3.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_G_pad_2 (.PACKAGE_PIN(ADV_G[2]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1848));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_G_pad_2.PIN_TYPE = 6'b011001;
    defparam ADV_G_pad_2.PULLUP = 1'b0;
    defparam ADV_G_pad_2.NEG_TRIGGER = 1'b0;
    defparam ADV_G_pad_2.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_G_pad_1 (.PACKAGE_PIN(ADV_G[1]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1849));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_G_pad_1.PIN_TYPE = 6'b011001;
    defparam ADV_G_pad_1.PULLUP = 1'b0;
    defparam ADV_G_pad_1.NEG_TRIGGER = 1'b0;
    defparam ADV_G_pad_1.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_G_pad_0 (.PACKAGE_PIN(ADV_G[0]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1850));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_G_pad_0.PIN_TYPE = 6'b011001;
    defparam ADV_G_pad_0.PULLUP = 1'b0;
    defparam ADV_G_pad_0.NEG_TRIGGER = 1'b0;
    defparam ADV_G_pad_0.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_B_pad_7 (.PACKAGE_PIN(ADV_B[7]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(ADV_B_c));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_B_pad_7.PIN_TYPE = 6'b011001;
    defparam ADV_B_pad_7.PULLUP = 1'b0;
    defparam ADV_B_pad_7.NEG_TRIGGER = 1'b0;
    defparam ADV_B_pad_7.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_B_pad_6 (.PACKAGE_PIN(ADV_B[6]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1844));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_B_pad_6.PIN_TYPE = 6'b011001;
    defparam ADV_B_pad_6.PULLUP = 1'b0;
    defparam ADV_B_pad_6.NEG_TRIGGER = 1'b0;
    defparam ADV_B_pad_6.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_B_pad_5 (.PACKAGE_PIN(ADV_B[5]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1845));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_B_pad_5.PIN_TYPE = 6'b011001;
    defparam ADV_B_pad_5.PULLUP = 1'b0;
    defparam ADV_B_pad_5.NEG_TRIGGER = 1'b0;
    defparam ADV_B_pad_5.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_B_pad_4 (.PACKAGE_PIN(ADV_B[4]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1846));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_B_pad_4.PIN_TYPE = 6'b011001;
    defparam ADV_B_pad_4.PULLUP = 1'b0;
    defparam ADV_B_pad_4.NEG_TRIGGER = 1'b0;
    defparam ADV_B_pad_4.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_B_pad_3 (.PACKAGE_PIN(ADV_B[3]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1847));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_B_pad_3.PIN_TYPE = 6'b011001;
    defparam ADV_B_pad_3.PULLUP = 1'b0;
    defparam ADV_B_pad_3.NEG_TRIGGER = 1'b0;
    defparam ADV_B_pad_3.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_B_pad_2 (.PACKAGE_PIN(ADV_B[2]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1848));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_B_pad_2.PIN_TYPE = 6'b011001;
    defparam ADV_B_pad_2.PULLUP = 1'b0;
    defparam ADV_B_pad_2.NEG_TRIGGER = 1'b0;
    defparam ADV_B_pad_2.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_B_pad_1 (.PACKAGE_PIN(ADV_B[1]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1849));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_B_pad_1.PIN_TYPE = 6'b011001;
    defparam ADV_B_pad_1.PULLUP = 1'b0;
    defparam ADV_B_pad_1.NEG_TRIGGER = 1'b0;
    defparam ADV_B_pad_1.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_B_pad_0 (.PACKAGE_PIN(ADV_B[0]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(n1850));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_B_pad_0.PIN_TYPE = 6'b011001;
    defparam ADV_B_pad_0.PULLUP = 1'b0;
    defparam ADV_B_pad_0.NEG_TRIGGER = 1'b0;
    defparam ADV_B_pad_0.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_CLK_pad (.PACKAGE_PIN(ADV_CLK), .OUTPUT_ENABLE(VCC_net), .D_OUT_0(ADV_CLK_c));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_CLK_pad.PIN_TYPE = 6'b011001;
    defparam ADV_CLK_pad.PULLUP = 1'b0;
    defparam ADV_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam ADV_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_SYNC_N_pad (.PACKAGE_PIN(ADV_SYNC_N), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(GND_net));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_SYNC_N_pad.PIN_TYPE = 6'b011001;
    defparam ADV_SYNC_N_pad.PULLUP = 1'b0;
    defparam ADV_SYNC_N_pad.NEG_TRIGGER = 1'b0;
    defparam ADV_SYNC_N_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO ADV_BLANK_N_pad (.PACKAGE_PIN(ADV_BLANK_N), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(VCC_net));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam ADV_BLANK_N_pad.PIN_TYPE = 6'b011001;
    defparam ADV_BLANK_N_pad.PULLUP = 1'b0;
    defparam ADV_BLANK_N_pad.NEG_TRIGGER = 1'b0;
    defparam ADV_BLANK_N_pad.IO_STANDARD = "SB_LVCMOS";
    SB_GB_IO TVP_CLK_pad (.PACKAGE_PIN(TVP_CLK), .OUTPUT_ENABLE(VCC_net), 
            .GLOBAL_BUFFER_OUTPUT(TVP_CLK_c));   // ../main.v(3[13:20])
    defparam TVP_CLK_pad.PIN_TYPE = 6'b000001;
    defparam TVP_CLK_pad.PULLUP = 1'b0;
    defparam TVP_CLK_pad.NEG_TRIGGER = 1'b0;
    defparam TVP_CLK_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO TVP_HSYNC_pad (.PACKAGE_PIN(TVP_HSYNC), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(TVP_HSYNC_c));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam TVP_HSYNC_pad.PIN_TYPE = 6'b000001;
    defparam TVP_HSYNC_pad.PULLUP = 1'b0;
    defparam TVP_HSYNC_pad.NEG_TRIGGER = 1'b0;
    defparam TVP_HSYNC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO TVP_VSYNC_pad (.PACKAGE_PIN(TVP_VSYNC), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(TVP_VSYNC_c));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam TVP_VSYNC_pad.PIN_TYPE = 6'b000001;
    defparam TVP_VSYNC_pad.PULLUP = 1'b0;
    defparam TVP_VSYNC_pad.NEG_TRIGGER = 1'b0;
    defparam TVP_VSYNC_pad.IO_STANDARD = "SB_LVCMOS";
    SB_IO TVP_VIDEO_pad_9 (.PACKAGE_PIN(TVP_VIDEO[9]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(TVP_VIDEO_c_9));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam TVP_VIDEO_pad_9.PIN_TYPE = 6'b000001;
    defparam TVP_VIDEO_pad_9.PULLUP = 1'b0;
    defparam TVP_VIDEO_pad_9.NEG_TRIGGER = 1'b0;
    defparam TVP_VIDEO_pad_9.IO_STANDARD = "SB_LVCMOS";
    SB_IO TVP_VIDEO_pad_8 (.PACKAGE_PIN(TVP_VIDEO[8]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(TVP_VIDEO_c_8));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam TVP_VIDEO_pad_8.PIN_TYPE = 6'b000001;
    defparam TVP_VIDEO_pad_8.PULLUP = 1'b0;
    defparam TVP_VIDEO_pad_8.NEG_TRIGGER = 1'b0;
    defparam TVP_VIDEO_pad_8.IO_STANDARD = "SB_LVCMOS";
    SB_IO TVP_VIDEO_pad_7 (.PACKAGE_PIN(TVP_VIDEO[7]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(TVP_VIDEO_c_7));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam TVP_VIDEO_pad_7.PIN_TYPE = 6'b000001;
    defparam TVP_VIDEO_pad_7.PULLUP = 1'b0;
    defparam TVP_VIDEO_pad_7.NEG_TRIGGER = 1'b0;
    defparam TVP_VIDEO_pad_7.IO_STANDARD = "SB_LVCMOS";
    SB_IO TVP_VIDEO_pad_6 (.PACKAGE_PIN(TVP_VIDEO[6]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(TVP_VIDEO_c_6));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam TVP_VIDEO_pad_6.PIN_TYPE = 6'b000001;
    defparam TVP_VIDEO_pad_6.PULLUP = 1'b0;
    defparam TVP_VIDEO_pad_6.NEG_TRIGGER = 1'b0;
    defparam TVP_VIDEO_pad_6.IO_STANDARD = "SB_LVCMOS";
    SB_IO TVP_VIDEO_pad_5 (.PACKAGE_PIN(TVP_VIDEO[5]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(TVP_VIDEO_c_5));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam TVP_VIDEO_pad_5.PIN_TYPE = 6'b000001;
    defparam TVP_VIDEO_pad_5.PULLUP = 1'b0;
    defparam TVP_VIDEO_pad_5.NEG_TRIGGER = 1'b0;
    defparam TVP_VIDEO_pad_5.IO_STANDARD = "SB_LVCMOS";
    SB_IO TVP_VIDEO_pad_4 (.PACKAGE_PIN(TVP_VIDEO[4]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(TVP_VIDEO_c_4));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam TVP_VIDEO_pad_4.PIN_TYPE = 6'b000001;
    defparam TVP_VIDEO_pad_4.PULLUP = 1'b0;
    defparam TVP_VIDEO_pad_4.NEG_TRIGGER = 1'b0;
    defparam TVP_VIDEO_pad_4.IO_STANDARD = "SB_LVCMOS";
    SB_IO TVP_VIDEO_pad_3 (.PACKAGE_PIN(TVP_VIDEO[3]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(TVP_VIDEO_c_3));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam TVP_VIDEO_pad_3.PIN_TYPE = 6'b000001;
    defparam TVP_VIDEO_pad_3.PULLUP = 1'b0;
    defparam TVP_VIDEO_pad_3.NEG_TRIGGER = 1'b0;
    defparam TVP_VIDEO_pad_3.IO_STANDARD = "SB_LVCMOS";
    SB_IO TVP_VIDEO_pad_2 (.PACKAGE_PIN(TVP_VIDEO[2]), .OUTPUT_ENABLE(VCC_net), 
          .D_IN_0(TVP_VIDEO_c_2));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam TVP_VIDEO_pad_2.PIN_TYPE = 6'b000001;
    defparam TVP_VIDEO_pad_2.PULLUP = 1'b0;
    defparam TVP_VIDEO_pad_2.NEG_TRIGGER = 1'b0;
    defparam TVP_VIDEO_pad_2.IO_STANDARD = "SB_LVCMOS";
    SB_IO DEBUG_pad_0 (.PACKAGE_PIN(DEBUG[0]), .OUTPUT_ENABLE(VCC_net), 
          .D_OUT_0(GND_net));   // C:/lscc/iCEcube2.2017.08/LSE/userware/NT/SYNTHESIS_HEADERS/sb_ice40.v(502[8:13])
    defparam DEBUG_pad_0.PIN_TYPE = 6'b011001;
    defparam DEBUG_pad_0.PULLUP = 1'b0;
    defparam DEBUG_pad_0.NEG_TRIGGER = 1'b0;
    defparam DEBUG_pad_0.IO_STANDARD = "SB_LVCMOS";
    SB_DFFNSR ADV_R__i2 (.Q(n1849), .C(ADV_CLK_c), .D(TX_DATA[1]), .R(n2404));   // ../main.v(65[9] 69[5])
    SB_DFFNSR ADV_R__i3 (.Q(n1848), .C(ADV_CLK_c), .D(TX_DATA[2]), .R(n2404));   // ../main.v(65[9] 69[5])
    SB_DFFNSR ADV_R__i4 (.Q(n1847), .C(ADV_CLK_c), .D(TX_DATA[3]), .R(n2404));   // ../main.v(65[9] 69[5])
    SB_DFFNSR ADV_R__i5 (.Q(n1846), .C(ADV_CLK_c), .D(TX_DATA[4]), .R(n2404));   // ../main.v(65[9] 69[5])
    SB_DFFNSR ADV_R__i6 (.Q(n1845), .C(ADV_CLK_c), .D(TX_DATA[5]), .R(n2404));   // ../main.v(65[9] 69[5])
    SB_DFFNSR ADV_R__i7 (.Q(n1844), .C(ADV_CLK_c), .D(TX_DATA[6]), .R(n2404));   // ../main.v(65[9] 69[5])
    SB_DFFNSR ADV_R__i8 (.Q(ADV_B_c), .C(ADV_CLK_c), .D(TX_DATA[7]), .R(n2404));   // ../main.v(65[9] 69[5])
    SB_LUT4 i272_3_lut_3_lut (.I0(TVP_HSYNC_c), .I1(TVP_VSYNC_c), .I2(old_HS), 
            .I3(GND_net), .O(n2057));   // ../main.v(4[13:22])
    defparam i272_3_lut_3_lut.LUT_INIT = 16'h7373;
    SB_LUT4 i26_1_lut_rep_24 (.I0(TVP_HSYNC_c), .I1(GND_net), .I2(GND_net), 
            .I3(GND_net), .O(n3860));   // ../main.v(4[13:22])
    defparam i26_1_lut_rep_24.LUT_INIT = 16'h5555;
    SB_DFFNSR ADV_R__i1 (.Q(n1850), .C(ADV_CLK_c), .D(TX_DATA[0]), .R(n2404));   // ../main.v(65[9] 69[5])
    GND i1 (.Y(GND_net));
    TX_PLL tx_pll (.TVP_CLK_c(TVP_CLK_c), .VCC_net(VCC_net), .GND_net(GND_net), 
           .ADV_CLK_c(ADV_CLK_c)) /* synthesis syn_module_defined=1 */ ;   // ../main.v(20[9] 24[27])
    RAM line_buffer (.\TX_ADDR[11] (TX_ADDR[11]), .\TX_ADDR[12] (TX_ADDR[12]), 
        .TX_DATA({TX_DATA}), .ADV_CLK_c(ADV_CLK_c), .DEBUG_c_2(DEBUG_c_2), 
        .\RX_ADDR[0] (RX_ADDR[0]), .\RX_ADDR[1] (RX_ADDR[1]), .\RX_ADDR[2] (RX_ADDR[2]), 
        .\RX_ADDR[3] (RX_ADDR[3]), .\RX_ADDR[4] (RX_ADDR[4]), .\RX_ADDR[5] (RX_ADDR[5]), 
        .\RX_ADDR[6] (RX_ADDR[6]), .\RX_ADDR[7] (RX_ADDR[7]), .\RX_ADDR[8] (RX_ADDR[8]), 
        .\RX_ADDR[9] (RX_ADDR[9]), .\RX_ADDR[10] (RX_ADDR[10]), .n28(n28), 
        .n27(n27), .n26(n26), .n25(n25), .n24(n24), .n23(n23), .n22(n22), 
        .n21(n21), .n20(n20), .n19(n19), .n18(n18), .TVP_VIDEO_c_8(TVP_VIDEO_c_8), 
        .TVP_VIDEO_c_9(TVP_VIDEO_c_9), .TVP_CLK_c(TVP_CLK_c), .VCC_net(VCC_net), 
        .TVP_VIDEO_c_6(TVP_VIDEO_c_6), .TVP_VIDEO_c_7(TVP_VIDEO_c_7), .TVP_VIDEO_c_4(TVP_VIDEO_c_4), 
        .TVP_VIDEO_c_5(TVP_VIDEO_c_5), .TVP_VIDEO_c_2(TVP_VIDEO_c_2), .TVP_VIDEO_c_3(TVP_VIDEO_c_3), 
        .\RX_ADDR[11] (RX_ADDR[11]), .\RX_ADDR[12] (RX_ADDR[12]), .DEBUG_c_3(DEBUG_c_3), 
        .DEBUG_c_5(DEBUG_c_5), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // ../main.v(72[6] 78[21])
    
endmodule
//
// Verilog Description of module RX
//

module RX (\RX_ADDR[6] , GND_net, \RX_ADDR[5] , \RX_ADDR[11] , \RX_ADDR[2] , 
           DEBUG_c_5, TVP_VSYNC_c, \RX_ADDR[4] , \RX_ADDR[3] , \RX_ADDR[0] , 
           \RX_ADDR[10] , VCC_net, \RX_ADDR[1] , \RX_ADDR[9] , \RX_ADDR[12] , 
           TVP_CLK_c, \RX_ADDR[8] , DEBUG_c_3, \RX_ADDR[7] , TVP_HSYNC_c, 
           old_HS, DEBUG_c_6, n3860, n2057, LED_c) /* synthesis syn_module_defined=1 */ ;
    output \RX_ADDR[6] ;
    input GND_net;
    output \RX_ADDR[5] ;
    output \RX_ADDR[11] ;
    output \RX_ADDR[2] ;
    output DEBUG_c_5;
    input TVP_VSYNC_c;
    output \RX_ADDR[4] ;
    output \RX_ADDR[3] ;
    output \RX_ADDR[0] ;
    output \RX_ADDR[10] ;
    input VCC_net;
    output \RX_ADDR[1] ;
    output \RX_ADDR[9] ;
    output \RX_ADDR[12] ;
    input TVP_CLK_c;
    output \RX_ADDR[8] ;
    output DEBUG_c_3;
    output \RX_ADDR[7] ;
    input TVP_HSYNC_c;
    output old_HS;
    output DEBUG_c_6;
    input n3860;
    input n2057;
    output LED_c;
    
    wire TVP_CLK_c /* synthesis SET_AS_NETWORK=TVP_CLK_c, is_clock=1 */ ;   // ../main.v(3[13:20])
    
    wire n3328, n3329;
    wire [13:0]n122;
    
    wire n3327, n3333, n3324, n3325, n3334, n2773, n2753, n2777, 
        n3332, n3323, n3331, n3854, n3326, BRAM_ADDR_13__N_31, n3330, 
        n3335, n2755, n2757, n2759, n2761, n2771, n2769, n2763, 
        n2767, n2765;
    
    SB_CARRY add_12_8 (.CI(n3328), .I0(\RX_ADDR[6] ), .I1(GND_net), .CO(n3329));
    SB_LUT4 add_12_7_lut (.I0(GND_net), .I1(\RX_ADDR[5] ), .I2(GND_net), 
            .I3(n3327), .O(n122[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_13_lut (.I0(GND_net), .I1(\RX_ADDR[11] ), .I2(GND_net), 
            .I3(n3333), .O(n122[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_13_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_4 (.CI(n3324), .I0(\RX_ADDR[2] ), .I1(GND_net), .CO(n3325));
    SB_CARRY add_12_13 (.CI(n3333), .I0(\RX_ADDR[11] ), .I1(GND_net), 
            .CO(n3334));
    SB_LUT4 i1502_3_lut_4_lut (.I0(DEBUG_c_5), .I1(TVP_VSYNC_c), .I2(n122[4]), 
            .I3(\RX_ADDR[4] ), .O(n2773));
    defparam i1502_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i1482_3_lut_4_lut (.I0(DEBUG_c_5), .I1(TVP_VSYNC_c), .I2(n122[3]), 
            .I3(\RX_ADDR[3] ), .O(n2753));
    defparam i1482_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i1506_3_lut_4_lut (.I0(DEBUG_c_5), .I1(TVP_VSYNC_c), .I2(n122[0]), 
            .I3(\RX_ADDR[0] ), .O(n2777));
    defparam i1506_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 add_12_12_lut (.I0(GND_net), .I1(\RX_ADDR[10] ), .I2(GND_net), 
            .I3(n3332), .O(n122[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_7 (.CI(n3327), .I0(\RX_ADDR[5] ), .I1(GND_net), .CO(n3328));
    SB_CARRY add_12_2 (.CI(VCC_net), .I0(\RX_ADDR[0] ), .I1(GND_net), 
            .CO(n3323));
    SB_CARRY add_12_12 (.CI(n3332), .I0(\RX_ADDR[10] ), .I1(GND_net), 
            .CO(n3333));
    SB_LUT4 add_12_3_lut (.I0(GND_net), .I1(\RX_ADDR[1] ), .I2(GND_net), 
            .I3(n3323), .O(n122[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_3_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_11_lut (.I0(GND_net), .I1(\RX_ADDR[9] ), .I2(GND_net), 
            .I3(n3331), .O(n122[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2393_2_lut_rep_18 (.I0(DEBUG_c_5), .I1(TVP_VSYNC_c), .I2(GND_net), 
            .I3(GND_net), .O(n3854));
    defparam i2393_2_lut_rep_18.LUT_INIT = 16'hbbbb;
    SB_CARRY add_12_11 (.CI(n3331), .I0(\RX_ADDR[9] ), .I1(GND_net), .CO(n3332));
    SB_CARRY add_12_3 (.CI(n3323), .I0(\RX_ADDR[1] ), .I1(GND_net), .CO(n3324));
    SB_LUT4 add_12_6_lut (.I0(GND_net), .I1(\RX_ADDR[4] ), .I2(GND_net), 
            .I3(n3326), .O(n122[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_6 (.CI(n3326), .I0(\RX_ADDR[4] ), .I1(GND_net), .CO(n3327));
    SB_DFFESR BRAM_ADDR__i12 (.Q(\RX_ADDR[12] ), .C(TVP_CLK_c), .E(n3854), 
            .D(n122[12]), .R(BRAM_ADDR_13__N_31));   // ../rx.v(51[12] 60[8])
    SB_DFFESR BRAM_ADDR__i11 (.Q(\RX_ADDR[11] ), .C(TVP_CLK_c), .E(n3854), 
            .D(n122[11]), .R(BRAM_ADDR_13__N_31));   // ../rx.v(51[12] 60[8])
    SB_LUT4 add_12_5_lut (.I0(GND_net), .I1(\RX_ADDR[3] ), .I2(GND_net), 
            .I3(n3325), .O(n122[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_10_lut (.I0(GND_net), .I1(\RX_ADDR[8] ), .I2(GND_net), 
            .I3(n3330), .O(n122[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_2_lut (.I0(GND_net), .I1(\RX_ADDR[0] ), .I2(GND_net), 
            .I3(VCC_net), .O(n122[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_12_15_lut (.I0(GND_net), .I1(DEBUG_c_3), .I2(GND_net), 
            .I3(n3335), .O(n122[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_15_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_10 (.CI(n3330), .I0(\RX_ADDR[8] ), .I1(GND_net), .CO(n3331));
    SB_LUT4 add_12_9_lut (.I0(GND_net), .I1(\RX_ADDR[7] ), .I2(GND_net), 
            .I3(n3329), .O(n122[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_12_5 (.CI(n3325), .I0(\RX_ADDR[3] ), .I1(GND_net), .CO(n3326));
    SB_CARRY add_12_9 (.CI(n3329), .I0(\RX_ADDR[7] ), .I1(GND_net), .CO(n3330));
    SB_LUT4 add_12_14_lut (.I0(GND_net), .I1(\RX_ADDR[12] ), .I2(GND_net), 
            .I3(n3334), .O(n122[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_14_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1484_3_lut_4_lut (.I0(DEBUG_c_5), .I1(TVP_VSYNC_c), .I2(n122[2]), 
            .I3(\RX_ADDR[2] ), .O(n2755));
    defparam i1484_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_CARRY add_12_14 (.CI(n3334), .I0(\RX_ADDR[12] ), .I1(GND_net), 
            .CO(n3335));
    SB_DFFSR BRAM_ADDR__i0 (.Q(\RX_ADDR[0] ), .C(TVP_CLK_c), .D(n2777), 
            .R(BRAM_ADDR_13__N_31));   // ../rx.v(51[12] 60[8])
    SB_LUT4 i1486_3_lut_4_lut (.I0(DEBUG_c_5), .I1(TVP_VSYNC_c), .I2(n122[1]), 
            .I3(\RX_ADDR[1] ), .O(n2757));
    defparam i1486_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_LUT4 i1488_3_lut_4_lut (.I0(DEBUG_c_5), .I1(TVP_VSYNC_c), .I2(n122[13]), 
            .I3(DEBUG_c_3), .O(n2759));
    defparam i1488_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_DFFSR BRAM_ADDR__i4 (.Q(\RX_ADDR[4] ), .C(TVP_CLK_c), .D(n2773), 
            .R(BRAM_ADDR_13__N_31));   // ../rx.v(51[12] 60[8])
    SB_LUT4 i1490_3_lut_4_lut (.I0(DEBUG_c_5), .I1(TVP_VSYNC_c), .I2(n122[10]), 
            .I3(\RX_ADDR[10] ), .O(n2761));
    defparam i1490_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_DFFSR BRAM_ADDR__i5 (.Q(\RX_ADDR[5] ), .C(TVP_CLK_c), .D(n2771), 
            .R(BRAM_ADDR_13__N_31));   // ../rx.v(51[12] 60[8])
    SB_LUT4 add_12_8_lut (.I0(GND_net), .I1(\RX_ADDR[6] ), .I2(GND_net), 
            .I3(n3328), .O(n122[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_8_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR BRAM_ADDR__i6 (.Q(\RX_ADDR[6] ), .C(TVP_CLK_c), .D(n2769), 
            .R(BRAM_ADDR_13__N_31));   // ../rx.v(51[12] 60[8])
    SB_LUT4 i1492_3_lut_4_lut (.I0(DEBUG_c_5), .I1(TVP_VSYNC_c), .I2(n122[9]), 
            .I3(\RX_ADDR[9] ), .O(n2763));
    defparam i1492_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_DFFSR BRAM_ADDR__i7 (.Q(\RX_ADDR[7] ), .C(TVP_CLK_c), .D(n2767), 
            .R(BRAM_ADDR_13__N_31));   // ../rx.v(51[12] 60[8])
    SB_DFFSR BRAM_ADDR__i8 (.Q(\RX_ADDR[8] ), .C(TVP_CLK_c), .D(n2765), 
            .R(BRAM_ADDR_13__N_31));   // ../rx.v(51[12] 60[8])
    SB_DFFSR BRAM_ADDR__i9 (.Q(\RX_ADDR[9] ), .C(TVP_CLK_c), .D(n2763), 
            .R(BRAM_ADDR_13__N_31));   // ../rx.v(51[12] 60[8])
    SB_LUT4 i1494_3_lut_4_lut (.I0(DEBUG_c_5), .I1(TVP_VSYNC_c), .I2(n122[8]), 
            .I3(\RX_ADDR[8] ), .O(n2765));
    defparam i1494_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_DFFSR BRAM_ADDR__i10 (.Q(\RX_ADDR[10] ), .C(TVP_CLK_c), .D(n2761), 
            .R(BRAM_ADDR_13__N_31));   // ../rx.v(51[12] 60[8])
    SB_LUT4 i1496_3_lut_4_lut (.I0(DEBUG_c_5), .I1(TVP_VSYNC_c), .I2(n122[7]), 
            .I3(\RX_ADDR[7] ), .O(n2767));
    defparam i1496_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_DFFSR BRAM_ADDR__i13 (.Q(DEBUG_c_3), .C(TVP_CLK_c), .D(n2759), 
            .R(BRAM_ADDR_13__N_31));   // ../rx.v(51[12] 60[8])
    SB_LUT4 i1498_3_lut_4_lut (.I0(DEBUG_c_5), .I1(TVP_VSYNC_c), .I2(n122[6]), 
            .I3(\RX_ADDR[6] ), .O(n2769));
    defparam i1498_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_DFFSR BRAM_ADDR__i1 (.Q(\RX_ADDR[1] ), .C(TVP_CLK_c), .D(n2757), 
            .R(BRAM_ADDR_13__N_31));   // ../rx.v(51[12] 60[8])
    SB_LUT4 i1500_3_lut_4_lut (.I0(DEBUG_c_5), .I1(TVP_VSYNC_c), .I2(n122[5]), 
            .I3(\RX_ADDR[5] ), .O(n2771));
    defparam i1500_3_lut_4_lut.LUT_INIT = 16'hf4b0;
    SB_DFFSR BRAM_ADDR__i2 (.Q(\RX_ADDR[2] ), .C(TVP_CLK_c), .D(n2755), 
            .R(BRAM_ADDR_13__N_31));   // ../rx.v(51[12] 60[8])
    SB_LUT4 add_12_4_lut (.I0(GND_net), .I1(\RX_ADDR[2] ), .I2(GND_net), 
            .I3(n3324), .O(n122[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_12_4_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR BRAM_ADDR__i3 (.Q(\RX_ADDR[3] ), .C(TVP_CLK_c), .D(n2753), 
            .R(BRAM_ADDR_13__N_31));   // ../rx.v(51[12] 60[8])
    O_COUNTER rx_counter (.TVP_CLK_c(TVP_CLK_c), .VCC_net(VCC_net), .GND_net(GND_net), 
            .TVP_HSYNC_c(TVP_HSYNC_c), .old_HS(old_HS), .TVP_VSYNC_c(TVP_VSYNC_c), 
            .DEBUG_c_6(DEBUG_c_6), .n3860(n3860), .n2057(n2057), .BRAM_ADDR_13__N_31(BRAM_ADDR_13__N_31), 
            .LED_c(LED_c), .DEBUG_c_5(DEBUG_c_5)) /* synthesis syn_module_defined=1 */ ;   // ../rx.v(41[15] 49[41])
    
endmodule
//
// Verilog Description of module O_COUNTER
//

module O_COUNTER (TVP_CLK_c, VCC_net, GND_net, TVP_HSYNC_c, old_HS, 
            TVP_VSYNC_c, DEBUG_c_6, n3860, n2057, BRAM_ADDR_13__N_31, 
            LED_c, DEBUG_c_5) /* synthesis syn_module_defined=1 */ ;
    input TVP_CLK_c;
    input VCC_net;
    input GND_net;
    input TVP_HSYNC_c;
    output old_HS;
    input TVP_VSYNC_c;
    output DEBUG_c_6;
    input n3860;
    input n2057;
    output BRAM_ADDR_13__N_31;
    output LED_c;
    output DEBUG_c_5;
    
    wire TVP_CLK_c /* synthesis SET_AS_NETWORK=TVP_CLK_c, is_clock=1 */ ;   // ../main.v(3[13:20])
    wire [5:0]n29;
    
    wire n3862;
    wire [5:0]FRAME_COUNTER;   // ../o_counter.v(46[19:32])
    
    wire n2562;
    wire [8:0]Y;   // ../o_counter.v(48[19:20])
    
    wire n3349, PULSE_1HZ_N_94, SYNC_N_96;
    wire [9:0]n45;
    wire [9:0]n79;
    
    wire n3387;
    wire [8:0]n303;
    
    wire PULSE_1HZ_N_92;
    wire [9:0]X;   // ../o_counter.v(47[19:20])
    
    wire n3365, n3364, n3363, n3362, n3361, n3360, n3359, n3547, 
        n14, n15, n3613, n3646, n4, n11, n3391, n3390, n3389, 
        n3388, n3358, n3357, n3861, n3657, n28, n3356, n3355, 
        n3619, n3648, n3354, n3353, n3352, n3351, n3350, n7, 
        n10_adj_570, n3693;
    
    SB_DFFESR FRAME_COUNTER_264__i2 (.Q(FRAME_COUNTER[2]), .C(TVP_CLK_c), 
            .E(n3862), .D(n29[2]), .R(n2562));   // ../o_counter.v(72[46:63])
    SB_CARRY add_65_2 (.CI(VCC_net), .I0(Y[0]), .I1(GND_net), .CO(n3349));
    SB_DFF old_HS_50 (.Q(old_HS), .C(TVP_CLK_c), .D(TVP_HSYNC_c));   // ../o_counter.v(51[16] 80[12])
    SB_DFFESR FRAME_COUNTER_264__i1 (.Q(FRAME_COUNTER[1]), .C(TVP_CLK_c), 
            .E(n3862), .D(n29[1]), .R(n2562));   // ../o_counter.v(72[46:63])
    SB_DFF old_VS_51 (.Q(PULSE_1HZ_N_94), .C(TVP_CLK_c), .D(TVP_VSYNC_c));   // ../o_counter.v(51[16] 80[12])
    SB_DFF SYNC_45 (.Q(DEBUG_c_6), .C(TVP_CLK_c), .D(SYNC_N_96));   // ../o_counter.v(51[16] 80[12])
    SB_DFFSR X_263__i0 (.Q(n79[0]), .C(TVP_CLK_c), .D(n45[0]), .R(n3860));   // ../o_counter.v(62[26:31])
    SB_CARRY FRAME_COUNTER_264_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(FRAME_COUNTER[0]), 
            .CO(n3387));
    SB_LUT4 FRAME_COUNTER_264_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(FRAME_COUNTER[0]), 
            .I3(VCC_net), .O(n29[0])) /* synthesis syn_instantiated=1 */ ;
    defparam FRAME_COUNTER_264_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR Y__i1 (.Q(Y[1]), .C(TVP_CLK_c), .E(n2057), .D(n303[1]), 
            .R(BRAM_ADDR_13__N_31));   // ../o_counter.v(51[16] 80[12])
    SB_DFFESR FRAME_COUNTER_264__i4 (.Q(FRAME_COUNTER[4]), .C(TVP_CLK_c), 
            .E(n3862), .D(n29[4]), .R(n2562));   // ../o_counter.v(72[46:63])
    SB_DFFESR Y__i2 (.Q(Y[2]), .C(TVP_CLK_c), .E(n2057), .D(n303[2]), 
            .R(BRAM_ADDR_13__N_31));   // ../o_counter.v(51[16] 80[12])
    SB_DFFESR Y__i3 (.Q(Y[3]), .C(TVP_CLK_c), .E(n2057), .D(n303[3]), 
            .R(BRAM_ADDR_13__N_31));   // ../o_counter.v(51[16] 80[12])
    SB_DFFESR Y__i4 (.Q(Y[4]), .C(TVP_CLK_c), .E(n2057), .D(n303[4]), 
            .R(BRAM_ADDR_13__N_31));   // ../o_counter.v(51[16] 80[12])
    SB_DFFESR FRAME_COUNTER_264__i3 (.Q(FRAME_COUNTER[3]), .C(TVP_CLK_c), 
            .E(n3862), .D(n29[3]), .R(n2562));   // ../o_counter.v(72[46:63])
    SB_DFFESR Y__i5 (.Q(Y[5]), .C(TVP_CLK_c), .E(n2057), .D(n303[5]), 
            .R(BRAM_ADDR_13__N_31));   // ../o_counter.v(51[16] 80[12])
    SB_DFFE PULSE_1HZ_48 (.Q(LED_c), .C(TVP_CLK_c), .E(n3862), .D(PULSE_1HZ_N_92));   // ../o_counter.v(51[16] 80[12])
    SB_LUT4 X_263_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(X[9]), 
            .I3(n3365), .O(n45[9])) /* synthesis syn_instantiated=1 */ ;
    defparam X_263_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 X_263_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(X[8]), 
            .I3(n3364), .O(n45[8])) /* synthesis syn_instantiated=1 */ ;
    defparam X_263_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY X_263_add_4_10 (.CI(n3364), .I0(GND_net), .I1(X[8]), .CO(n3365));
    SB_LUT4 X_263_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(X[7]), 
            .I3(n3363), .O(n45[7])) /* synthesis syn_instantiated=1 */ ;
    defparam X_263_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY X_263_add_4_9 (.CI(n3363), .I0(GND_net), .I1(X[7]), .CO(n3364));
    SB_LUT4 X_263_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(X[6]), 
            .I3(n3362), .O(n45[6])) /* synthesis syn_instantiated=1 */ ;
    defparam X_263_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY X_263_add_4_8 (.CI(n3362), .I0(GND_net), .I1(X[6]), .CO(n3363));
    SB_LUT4 X_263_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(X[5]), 
            .I3(n3361), .O(n45[5])) /* synthesis syn_instantiated=1 */ ;
    defparam X_263_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY X_263_add_4_7 (.CI(n3361), .I0(GND_net), .I1(X[5]), .CO(n3362));
    SB_LUT4 X_263_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(X[4]), 
            .I3(n3360), .O(n45[4])) /* synthesis syn_instantiated=1 */ ;
    defparam X_263_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY X_263_add_4_6 (.CI(n3360), .I0(GND_net), .I1(X[4]), .CO(n3361));
    SB_LUT4 X_263_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(X[3]), 
            .I3(n3359), .O(n45[3])) /* synthesis syn_instantiated=1 */ ;
    defparam X_263_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY X_263_add_4_5 (.CI(n3359), .I0(GND_net), .I1(X[3]), .CO(n3360));
    SB_LUT4 i2_3_lut (.I0(X[4]), .I1(X[5]), .I2(X[3]), .I3(GND_net), 
            .O(n3547));   // ../o_counter.v(82[61:90])
    defparam i2_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1_2_lut (.I0(Y[0]), .I1(Y[1]), .I2(GND_net), .I3(GND_net), 
            .O(n14));   // ../o_counter.v(51[16] 80[12])
    defparam i1_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i1_4_lut (.I0(Y[4]), .I1(Y[2]), .I2(Y[3]), .I3(n14), .O(n15));   // ../o_counter.v(51[16] 80[12])
    defparam i1_4_lut.LUT_INIT = 16'haaa8;
    SB_LUT4 i2251_3_lut (.I0(X[6]), .I1(X[7]), .I2(n3547), .I3(GND_net), 
            .O(n3613));
    defparam i2251_3_lut.LUT_INIT = 16'hc8c8;
    SB_LUT4 i2_3_lut_adj_15 (.I0(X[6]), .I1(X[7]), .I2(n3547), .I3(GND_net), 
            .O(n3646));
    defparam i2_3_lut_adj_15.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_adj_16 (.I0(Y[0]), .I1(Y[2]), .I2(GND_net), .I3(GND_net), 
            .O(n4));
    defparam i1_2_lut_adj_16.LUT_INIT = 16'heeee;
    SB_LUT4 i1294_2_lut_3_lut (.I0(PULSE_1HZ_N_94), .I1(TVP_VSYNC_c), .I2(n11), 
            .I3(GND_net), .O(n2562));   // ../o_counter.v(65[16] 75[19])
    defparam i1294_2_lut_3_lut.LUT_INIT = 16'h0202;
    SB_LUT4 FRAME_COUNTER_264_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(FRAME_COUNTER[5]), 
            .I3(n3391), .O(n29[5])) /* synthesis syn_instantiated=1 */ ;
    defparam FRAME_COUNTER_264_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 FRAME_COUNTER_264_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(FRAME_COUNTER[4]), 
            .I3(n3390), .O(n29[4])) /* synthesis syn_instantiated=1 */ ;
    defparam FRAME_COUNTER_264_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY FRAME_COUNTER_264_add_4_6 (.CI(n3390), .I0(GND_net), .I1(FRAME_COUNTER[4]), 
            .CO(n3391));
    SB_LUT4 FRAME_COUNTER_264_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(FRAME_COUNTER[3]), 
            .I3(n3389), .O(n29[3])) /* synthesis syn_instantiated=1 */ ;
    defparam FRAME_COUNTER_264_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY FRAME_COUNTER_264_add_4_5 (.CI(n3389), .I0(GND_net), .I1(FRAME_COUNTER[3]), 
            .CO(n3390));
    SB_LUT4 FRAME_COUNTER_264_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(FRAME_COUNTER[2]), 
            .I3(n3388), .O(n29[2])) /* synthesis syn_instantiated=1 */ ;
    defparam FRAME_COUNTER_264_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY FRAME_COUNTER_264_add_4_4 (.CI(n3388), .I0(GND_net), .I1(FRAME_COUNTER[2]), 
            .CO(n3389));
    SB_LUT4 FRAME_COUNTER_264_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(FRAME_COUNTER[1]), 
            .I3(n3387), .O(n29[1])) /* synthesis syn_instantiated=1 */ ;
    defparam FRAME_COUNTER_264_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY FRAME_COUNTER_264_add_4_3 (.CI(n3387), .I0(GND_net), .I1(FRAME_COUNTER[1]), 
            .CO(n3388));
    SB_LUT4 X_263_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(n79[2]), 
            .I3(n3358), .O(n45[2])) /* synthesis syn_instantiated=1 */ ;
    defparam X_263_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY X_263_add_4_4 (.CI(n3358), .I0(GND_net), .I1(n79[2]), .CO(n3359));
    SB_LUT4 X_263_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(n79[1]), 
            .I3(n3357), .O(n45[1])) /* synthesis syn_instantiated=1 */ ;
    defparam X_263_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY X_263_add_4_3 (.CI(n3357), .I0(GND_net), .I1(n79[1]), .CO(n3358));
    SB_LUT4 X_263_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(n79[0]), 
            .I3(VCC_net), .O(n45[0])) /* synthesis syn_instantiated=1 */ ;
    defparam X_263_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i2_4_lut (.I0(Y[7]), .I1(Y[8]), .I2(n15), .I3(n3861), .O(n3657));   // ../o_counter.v(82[28:148])
    defparam i2_4_lut.LUT_INIT = 16'h8880;
    SB_DFFSR X_263__i1 (.Q(n79[1]), .C(TVP_CLK_c), .D(n45[1]), .R(n3860));   // ../o_counter.v(62[26:31])
    SB_DFFSR X_263__i2 (.Q(n79[2]), .C(TVP_CLK_c), .D(n45[2]), .R(n3860));   // ../o_counter.v(62[26:31])
    SB_LUT4 i35_4_lut (.I0(X[8]), .I1(n3646), .I2(X[9]), .I3(n3613), 
            .O(n28));   // ../o_counter.v(82[28:148])
    defparam i35_4_lut.LUT_INIT = 16'he0e5;
    SB_LUT4 i140_2_lut_rep_26 (.I0(PULSE_1HZ_N_94), .I1(TVP_VSYNC_c), .I2(GND_net), 
            .I3(GND_net), .O(n3862));   // ../o_counter.v(65[16] 75[19])
    defparam i140_2_lut_rep_26.LUT_INIT = 16'h2222;
    SB_CARRY X_263_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(n79[0]), .CO(n3357));
    SB_LUT4 add_65_10_lut (.I0(GND_net), .I1(Y[8]), .I2(GND_net), .I3(n3356), 
            .O(n303[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_65_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_65_9_lut (.I0(GND_net), .I1(Y[7]), .I2(GND_net), .I3(n3355), 
            .O(n303[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_65_9_lut.LUT_INIT = 16'hC33C;
    SB_DFFSR X_263__i3 (.Q(X[3]), .C(TVP_CLK_c), .D(n45[3]), .R(n3860));   // ../o_counter.v(62[26:31])
    SB_DFFSR X_263__i4 (.Q(X[4]), .C(TVP_CLK_c), .D(n45[4]), .R(n3860));   // ../o_counter.v(62[26:31])
    SB_DFFSR X_263__i5 (.Q(X[5]), .C(TVP_CLK_c), .D(n45[5]), .R(n3860));   // ../o_counter.v(62[26:31])
    SB_DFFSR X_263__i6 (.Q(X[6]), .C(TVP_CLK_c), .D(n45[6]), .R(n3860));   // ../o_counter.v(62[26:31])
    SB_DFFSR X_263__i7 (.Q(X[7]), .C(TVP_CLK_c), .D(n45[7]), .R(n3860));   // ../o_counter.v(62[26:31])
    SB_DFFSR X_263__i8 (.Q(X[8]), .C(TVP_CLK_c), .D(n45[8]), .R(n3860));   // ../o_counter.v(62[26:31])
    SB_DFFSR X_263__i9 (.Q(X[9]), .C(TVP_CLK_c), .D(n45[9]), .R(n3860));   // ../o_counter.v(62[26:31])
    SB_LUT4 i2_3_lut_4_lut (.I0(Y[6]), .I1(Y[5]), .I2(Y[7]), .I3(Y[8]), 
            .O(n3619));   // ../o_counter.v(51[16] 80[12])
    defparam i2_3_lut_4_lut.LUT_INIT = 16'hfffe;
    SB_LUT4 i1_2_lut_rep_25 (.I0(Y[6]), .I1(Y[5]), .I2(GND_net), .I3(GND_net), 
            .O(n3861));   // ../o_counter.v(51[16] 80[12])
    defparam i1_2_lut_rep_25.LUT_INIT = 16'heeee;
    SB_LUT4 i2_4_lut_adj_17 (.I0(Y[1]), .I1(Y[4]), .I2(n4), .I3(Y[3]), 
            .O(n3648));
    defparam i2_4_lut_adj_17.LUT_INIT = 16'hc800;
    SB_LUT4 i2397_4_lut (.I0(n3648), .I1(n28), .I2(n3619), .I3(n3657), 
            .O(DEBUG_c_5));   // ../o_counter.v(82[28:148])
    defparam i2397_4_lut.LUT_INIT = 16'h0032;
    SB_DFFESR Y__i6 (.Q(Y[6]), .C(TVP_CLK_c), .E(n2057), .D(n303[6]), 
            .R(BRAM_ADDR_13__N_31));   // ../o_counter.v(51[16] 80[12])
    SB_CARRY add_65_9 (.CI(n3355), .I0(Y[7]), .I1(GND_net), .CO(n3356));
    SB_DFFESR Y__i7 (.Q(Y[7]), .C(TVP_CLK_c), .E(n2057), .D(n303[7]), 
            .R(BRAM_ADDR_13__N_31));   // ../o_counter.v(51[16] 80[12])
    SB_DFFESR Y__i8 (.Q(Y[8]), .C(TVP_CLK_c), .E(n2057), .D(n303[8]), 
            .R(BRAM_ADDR_13__N_31));   // ../o_counter.v(51[16] 80[12])
    SB_LUT4 add_65_8_lut (.I0(GND_net), .I1(Y[6]), .I2(GND_net), .I3(n3354), 
            .O(n303[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_65_8_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR Y__i0 (.Q(Y[0]), .C(TVP_CLK_c), .E(n2057), .D(n303[0]), 
            .R(BRAM_ADDR_13__N_31));   // ../o_counter.v(51[16] 80[12])
    SB_DFFESR FRAME_COUNTER_264__i0 (.Q(FRAME_COUNTER[0]), .C(TVP_CLK_c), 
            .E(n3862), .D(n29[0]), .R(n2562));   // ../o_counter.v(72[46:63])
    SB_CARRY add_65_8 (.CI(n3354), .I0(Y[6]), .I1(GND_net), .CO(n3355));
    SB_LUT4 add_65_7_lut (.I0(GND_net), .I1(Y[5]), .I2(GND_net), .I3(n3353), 
            .O(n303[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_65_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_65_7 (.CI(n3353), .I0(Y[5]), .I1(GND_net), .CO(n3354));
    SB_LUT4 add_65_6_lut (.I0(GND_net), .I1(Y[4]), .I2(GND_net), .I3(n3352), 
            .O(n303[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_65_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_65_6 (.CI(n3352), .I0(Y[4]), .I1(GND_net), .CO(n3353));
    SB_LUT4 add_65_5_lut (.I0(GND_net), .I1(Y[3]), .I2(GND_net), .I3(n3351), 
            .O(n303[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_65_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_65_5 (.CI(n3351), .I0(Y[3]), .I1(GND_net), .CO(n3352));
    SB_LUT4 add_65_4_lut (.I0(GND_net), .I1(Y[2]), .I2(GND_net), .I3(n3350), 
            .O(n303[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_65_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_65_4 (.CI(n3350), .I0(Y[2]), .I1(GND_net), .CO(n3351));
    SB_LUT4 i1_2_lut_adj_18 (.I0(FRAME_COUNTER[2]), .I1(FRAME_COUNTER[4]), 
            .I2(GND_net), .I3(GND_net), .O(n7));
    defparam i1_2_lut_adj_18.LUT_INIT = 16'hbbbb;
    SB_LUT4 i4_4_lut (.I0(Y[3]), .I1(Y[4]), .I2(Y[1]), .I3(n3619), .O(n10_adj_570));
    defparam i4_4_lut.LUT_INIT = 16'h0002;
    SB_LUT4 i2331_2_lut (.I0(FRAME_COUNTER[1]), .I1(FRAME_COUNTER[5]), .I2(GND_net), 
            .I3(GND_net), .O(n3693));
    defparam i2331_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i5_4_lut (.I0(n3693), .I1(n7), .I2(FRAME_COUNTER[3]), .I3(FRAME_COUNTER[0]), 
            .O(n11));
    defparam i5_4_lut.LUT_INIT = 16'hdfff;
    SB_LUT4 i1_2_lut_adj_19 (.I0(LED_c), .I1(n11), .I2(GND_net), .I3(GND_net), 
            .O(PULSE_1HZ_N_92));
    defparam i1_2_lut_adj_19.LUT_INIT = 16'h9999;
    SB_LUT4 i23_1_lut (.I0(TVP_VSYNC_c), .I1(GND_net), .I2(GND_net), .I3(GND_net), 
            .O(BRAM_ADDR_13__N_31));   // ../main.v(5[13:22])
    defparam i23_1_lut.LUT_INIT = 16'h5555;
    SB_LUT4 i5_3_lut (.I0(Y[2]), .I1(n10_adj_570), .I2(Y[0]), .I3(GND_net), 
            .O(SYNC_N_96));
    defparam i5_3_lut.LUT_INIT = 16'h0808;
    SB_LUT4 add_65_3_lut (.I0(GND_net), .I1(Y[1]), .I2(GND_net), .I3(n3349), 
            .O(n303[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_65_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_65_3 (.CI(n3349), .I0(Y[1]), .I1(GND_net), .CO(n3350));
    SB_DFFESR FRAME_COUNTER_264__i5 (.Q(FRAME_COUNTER[5]), .C(TVP_CLK_c), 
            .E(n3862), .D(n29[5]), .R(n2562));   // ../o_counter.v(72[46:63])
    SB_LUT4 add_65_2_lut (.I0(GND_net), .I1(Y[0]), .I2(GND_net), .I3(VCC_net), 
            .O(n303[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_65_2_lut.LUT_INIT = 16'hC33C;
    
endmodule
//
// Verilog Description of module TX
//

module TX (GND_net, ADV_HSYNC_c, ADV_CLK_c, ADV_VSYNC_c, n23, DEBUG_c_2, 
           \TX_ADDR[12] , n22, n18, n19, n20, n21, n24, n25, 
           n26, n27, \TX_ADDR[11] , n3852, n28, VCC_net, DEBUG_c_6, 
           n2404) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output ADV_HSYNC_c;
    input ADV_CLK_c;
    output ADV_VSYNC_c;
    output n23;
    output DEBUG_c_2;
    output \TX_ADDR[12] ;
    output n22;
    output n18;
    output n19;
    output n20;
    output n21;
    output n24;
    output n25;
    output n26;
    output n27;
    output \TX_ADDR[11] ;
    output n3852;
    output n28;
    input VCC_net;
    input DEBUG_c_6;
    output n2404;
    
    wire ADV_CLK_c /* synthesis SET_AS_NETWORK=ADV_CLK_c, is_clock=1 */ ;   // ../main.v(13[14:21])
    wire [13:0]ADDR_Y_COMPONENT;   // ../tx.v(64[16:32])
    wire [13:0]TX_ADDR;   // ../main.v(47[14:21])
    wire [99:0]Y_DELTA_PATTERN;   // ../tx.v(63[16:31])
    wire [13:0]n174;
    
    wire old_VGA_HS, n3864, n2125;
    wire [13:0]n206;
    
    wire n3853;
    wire [13:0]n190;
    
    wire n3348, n3865;
    wire [15:0]X_DELTA_PATTERN;   // ../tx.v(62[16:31])
    
    wire n2099, n3342, n3347, n3343, n3338, n3339, n3337, n3336, 
        n3341, n2321, n3346, n3549, n3855, n3859, n3340;
    wire [13:0]BRAM_ADDR_13__N_256;
    
    wire n2039, n2775, n3345, n3344;
    
    SB_LUT4 mux_12_i6_3_lut (.I0(ADDR_Y_COMPONENT[5]), .I1(TX_ADDR[5]), 
            .I2(Y_DELTA_PATTERN[0]), .I3(GND_net), .O(n174[5]));   // ../tx.v(79[30:81])
    defparam mux_12_i6_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF old_VGA_HS_39 (.Q(old_VGA_HS), .C(ADV_CLK_c), .D(ADV_HSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i99 (.Q(Y_DELTA_PATTERN[99]), .C(ADV_CLK_c), 
            .E(n3864), .D(Y_DELTA_PATTERN[0]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESR Y_DELTA_PATTERN_i98 (.Q(Y_DELTA_PATTERN[98]), .C(ADV_CLK_c), 
            .E(n2125), .D(Y_DELTA_PATTERN[99]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i97 (.Q(Y_DELTA_PATTERN[97]), .C(ADV_CLK_c), 
            .E(n2125), .D(Y_DELTA_PATTERN[98]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i96 (.Q(Y_DELTA_PATTERN[96]), .C(ADV_CLK_c), 
            .E(n2125), .D(Y_DELTA_PATTERN[97]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESR Y_DELTA_PATTERN_i95 (.Q(Y_DELTA_PATTERN[95]), .C(ADV_CLK_c), 
            .E(n2125), .D(Y_DELTA_PATTERN[96]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_LUT4 i1680_4_lut (.I0(n206[5]), .I1(ADV_VSYNC_c), .I2(n174[5]), 
            .I3(n3853), .O(n23));   // ../tx.v(68[12] 91[8])
    defparam i1680_4_lut.LUT_INIT = 16'h3022;
    SB_DFFESS Y_DELTA_PATTERN_i94 (.Q(Y_DELTA_PATTERN[94]), .C(ADV_CLK_c), 
            .E(n2125), .D(Y_DELTA_PATTERN[95]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESR Y_DELTA_PATTERN_i93 (.Q(Y_DELTA_PATTERN[93]), .C(ADV_CLK_c), 
            .E(n2125), .D(Y_DELTA_PATTERN[94]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i92 (.Q(Y_DELTA_PATTERN[92]), .C(ADV_CLK_c), 
            .E(n2125), .D(Y_DELTA_PATTERN[93]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i91 (.Q(Y_DELTA_PATTERN[91]), .C(ADV_CLK_c), 
            .E(n2125), .D(Y_DELTA_PATTERN[92]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESR Y_DELTA_PATTERN_i90 (.Q(Y_DELTA_PATTERN[90]), .C(ADV_CLK_c), 
            .E(n2125), .D(Y_DELTA_PATTERN[91]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i89 (.Q(Y_DELTA_PATTERN[89]), .C(ADV_CLK_c), 
            .E(n2125), .D(Y_DELTA_PATTERN[90]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i88 (.Q(Y_DELTA_PATTERN[88]), .C(ADV_CLK_c), 
            .E(n2125), .D(Y_DELTA_PATTERN[89]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESR Y_DELTA_PATTERN_i87 (.Q(Y_DELTA_PATTERN[87]), .C(ADV_CLK_c), 
            .E(n2125), .D(Y_DELTA_PATTERN[88]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_LUT4 add_13_15_lut (.I0(GND_net), .I1(DEBUG_c_2), .I2(GND_net), 
            .I3(n3348), .O(n190[13])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_15_lut.LUT_INIT = 16'hC33C;
    SB_DFFESS Y_DELTA_PATTERN_i86 (.Q(Y_DELTA_PATTERN[86]), .C(ADV_CLK_c), 
            .E(n2125), .D(Y_DELTA_PATTERN[87]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESR Y_DELTA_PATTERN_i85 (.Q(Y_DELTA_PATTERN[85]), .C(ADV_CLK_c), 
            .E(n2125), .D(Y_DELTA_PATTERN[86]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_LUT4 mux_12_i11_3_lut (.I0(ADDR_Y_COMPONENT[10]), .I1(TX_ADDR[10]), 
            .I2(Y_DELTA_PATTERN[0]), .I3(GND_net), .O(n174[10]));   // ../tx.v(79[30:81])
    defparam mux_12_i11_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESS Y_DELTA_PATTERN_i84 (.Q(Y_DELTA_PATTERN[84]), .C(ADV_CLK_c), 
            .E(n2125), .D(Y_DELTA_PATTERN[85]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i83 (.Q(Y_DELTA_PATTERN[83]), .C(ADV_CLK_c), 
            .E(n2125), .D(Y_DELTA_PATTERN[84]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESR Y_DELTA_PATTERN_i82 (.Q(Y_DELTA_PATTERN[82]), .C(ADV_CLK_c), 
            .E(n3865), .D(Y_DELTA_PATTERN[83]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i81 (.Q(Y_DELTA_PATTERN[81]), .C(ADV_CLK_c), 
            .E(n3865), .D(Y_DELTA_PATTERN[82]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i80 (.Q(Y_DELTA_PATTERN[80]), .C(ADV_CLK_c), 
            .E(n3865), .D(Y_DELTA_PATTERN[81]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_LUT4 mux_12_i7_3_lut (.I0(ADDR_Y_COMPONENT[6]), .I1(TX_ADDR[6]), 
            .I2(Y_DELTA_PATTERN[0]), .I3(GND_net), .O(n174[6]));   // ../tx.v(79[30:81])
    defparam mux_12_i7_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR Y_DELTA_PATTERN_i79 (.Q(Y_DELTA_PATTERN[79]), .C(ADV_CLK_c), 
            .E(n3865), .D(Y_DELTA_PATTERN[80]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i78 (.Q(Y_DELTA_PATTERN[78]), .C(ADV_CLK_c), 
            .E(n3865), .D(Y_DELTA_PATTERN[79]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESR Y_DELTA_PATTERN_i77 (.Q(Y_DELTA_PATTERN[77]), .C(ADV_CLK_c), 
            .E(n3865), .D(Y_DELTA_PATTERN[78]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i76 (.Q(Y_DELTA_PATTERN[76]), .C(ADV_CLK_c), 
            .E(n3865), .D(Y_DELTA_PATTERN[77]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i75 (.Q(Y_DELTA_PATTERN[75]), .C(ADV_CLK_c), 
            .E(n3865), .D(Y_DELTA_PATTERN[76]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESR Y_DELTA_PATTERN_i74 (.Q(Y_DELTA_PATTERN[74]), .C(ADV_CLK_c), 
            .E(n3865), .D(Y_DELTA_PATTERN[75]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i73 (.Q(Y_DELTA_PATTERN[73]), .C(ADV_CLK_c), 
            .E(n3865), .D(Y_DELTA_PATTERN[74]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i2 (.Q(Y_DELTA_PATTERN[2]), .C(ADV_CLK_c), 
            .E(n3865), .D(Y_DELTA_PATTERN[3]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESR Y_DELTA_PATTERN_i1 (.Q(Y_DELTA_PATTERN[1]), .C(ADV_CLK_c), 
            .E(n3864), .D(Y_DELTA_PATTERN[2]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS X_DELTA_PATTERN_i15 (.Q(X_DELTA_PATTERN[15]), .C(ADV_CLK_c), 
            .E(n2099), .D(X_DELTA_PATTERN[0]), .S(n3864));   // ../tx.v(68[12] 91[8])
    SB_LUT4 add_13_9_lut (.I0(GND_net), .I1(TX_ADDR[7]), .I2(GND_net), 
            .I3(n3342), .O(n190[7])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_9_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 add_13_14_lut (.I0(GND_net), .I1(\TX_ADDR[12] ), .I2(GND_net), 
            .I3(n3347), .O(n190[12])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_14_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR X_DELTA_PATTERN_i14 (.Q(X_DELTA_PATTERN[14]), .C(ADV_CLK_c), 
            .E(n2099), .D(X_DELTA_PATTERN[15]), .R(n3864));   // ../tx.v(68[12] 91[8])
    SB_CARRY add_13_9 (.CI(n3342), .I0(TX_ADDR[7]), .I1(GND_net), .CO(n3343));
    SB_LUT4 i1681_4_lut (.I0(n206[6]), .I1(ADV_VSYNC_c), .I2(n174[6]), 
            .I3(n3853), .O(n22));   // ../tx.v(68[12] 91[8])
    defparam i1681_4_lut.LUT_INIT = 16'h3022;
    SB_DFFESS X_DELTA_PATTERN_i13 (.Q(X_DELTA_PATTERN[13]), .C(ADV_CLK_c), 
            .E(n2099), .D(X_DELTA_PATTERN[14]), .S(n3864));   // ../tx.v(68[12] 91[8])
    SB_DFFESR X_DELTA_PATTERN_i12 (.Q(X_DELTA_PATTERN[12]), .C(ADV_CLK_c), 
            .E(n2099), .D(X_DELTA_PATTERN[13]), .R(n3864));   // ../tx.v(68[12] 91[8])
    SB_CARRY add_13_5 (.CI(n3338), .I0(TX_ADDR[3]), .I1(GND_net), .CO(n3339));
    SB_LUT4 add_13_4_lut (.I0(GND_net), .I1(TX_ADDR[2]), .I2(GND_net), 
            .I3(n3337), .O(n190[2])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_4_lut.LUT_INIT = 16'hC33C;
    SB_DFFESS X_DELTA_PATTERN_i11 (.Q(X_DELTA_PATTERN[11]), .C(ADV_CLK_c), 
            .E(n2099), .D(X_DELTA_PATTERN[12]), .S(n3864));   // ../tx.v(68[12] 91[8])
    SB_CARRY add_13_4 (.CI(n3337), .I0(TX_ADDR[2]), .I1(GND_net), .CO(n3338));
    SB_DFFESR X_DELTA_PATTERN_i10 (.Q(X_DELTA_PATTERN[10]), .C(ADV_CLK_c), 
            .E(n2099), .D(X_DELTA_PATTERN[11]), .R(n3864));   // ../tx.v(68[12] 91[8])
    SB_LUT4 add_13_3_lut (.I0(GND_net), .I1(TX_ADDR[1]), .I2(GND_net), 
            .I3(n3336), .O(n190[1])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_3_lut.LUT_INIT = 16'hC33C;
    SB_DFFESS X_DELTA_PATTERN_i9 (.Q(X_DELTA_PATTERN[9]), .C(ADV_CLK_c), 
            .E(n2099), .D(X_DELTA_PATTERN[10]), .S(n3864));   // ../tx.v(68[12] 91[8])
    SB_DFFESR X_DELTA_PATTERN_i8 (.Q(X_DELTA_PATTERN[8]), .C(ADV_CLK_c), 
            .E(n2099), .D(X_DELTA_PATTERN[9]), .R(n3864));   // ../tx.v(68[12] 91[8])
    SB_DFF BRAM_ADDR__i10 (.Q(TX_ADDR[10]), .C(ADV_CLK_c), .D(n18));   // ../tx.v(68[12] 91[8])
    SB_LUT4 add_13_8_lut (.I0(GND_net), .I1(TX_ADDR[6]), .I2(GND_net), 
            .I3(n3341), .O(n190[6])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_8_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_12_i8_3_lut (.I0(ADDR_Y_COMPONENT[7]), .I1(TX_ADDR[7]), 
            .I2(Y_DELTA_PATTERN[0]), .I3(GND_net), .O(n174[7]));   // ../tx.v(79[30:81])
    defparam mux_12_i8_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF BRAM_ADDR__i9 (.Q(TX_ADDR[9]), .C(ADV_CLK_c), .D(n19));   // ../tx.v(68[12] 91[8])
    SB_DFF BRAM_ADDR__i8 (.Q(TX_ADDR[8]), .C(ADV_CLK_c), .D(n20));   // ../tx.v(68[12] 91[8])
    SB_DFF BRAM_ADDR__i7 (.Q(TX_ADDR[7]), .C(ADV_CLK_c), .D(n21));   // ../tx.v(68[12] 91[8])
    SB_DFF BRAM_ADDR__i6 (.Q(TX_ADDR[6]), .C(ADV_CLK_c), .D(n22));   // ../tx.v(68[12] 91[8])
    SB_DFF BRAM_ADDR__i5 (.Q(TX_ADDR[5]), .C(ADV_CLK_c), .D(n23));   // ../tx.v(68[12] 91[8])
    SB_DFF BRAM_ADDR__i4 (.Q(TX_ADDR[4]), .C(ADV_CLK_c), .D(n24));   // ../tx.v(68[12] 91[8])
    SB_CARRY add_13_14 (.CI(n3347), .I0(\TX_ADDR[12] ), .I1(GND_net), 
            .CO(n3348));
    SB_DFF BRAM_ADDR__i3 (.Q(TX_ADDR[3]), .C(ADV_CLK_c), .D(n25));   // ../tx.v(68[12] 91[8])
    SB_DFF BRAM_ADDR__i2 (.Q(TX_ADDR[2]), .C(ADV_CLK_c), .D(n26));   // ../tx.v(68[12] 91[8])
    SB_DFF BRAM_ADDR__i1 (.Q(TX_ADDR[1]), .C(ADV_CLK_c), .D(n27));   // ../tx.v(68[12] 91[8])
    SB_DFFESR ADDR_Y_COMPONENT__i3 (.Q(ADDR_Y_COMPONENT[3]), .C(ADV_CLK_c), 
            .E(n2321), .D(TX_ADDR[3]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_LUT4 add_13_13_lut (.I0(GND_net), .I1(\TX_ADDR[11] ), .I2(GND_net), 
            .I3(n3346), .O(n190[11])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_13_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1682_4_lut (.I0(n206[7]), .I1(ADV_VSYNC_c), .I2(n174[7]), 
            .I3(n3853), .O(n21));   // ../tx.v(68[12] 91[8])
    defparam i1682_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 i1685_4_lut (.I0(n206[10]), .I1(ADV_VSYNC_c), .I2(n174[10]), 
            .I3(n3853), .O(n18));   // ../tx.v(68[12] 91[8])
    defparam i1685_4_lut.LUT_INIT = 16'h3022;
    SB_DFFESS Y_DELTA_PATTERN_i72 (.Q(Y_DELTA_PATTERN[72]), .C(ADV_CLK_c), 
            .E(n3864), .D(Y_DELTA_PATTERN[73]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESR Y_DELTA_PATTERN_i71 (.Q(Y_DELTA_PATTERN[71]), .C(ADV_CLK_c), 
            .E(n3865), .D(Y_DELTA_PATTERN[72]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i70 (.Q(Y_DELTA_PATTERN[70]), .C(ADV_CLK_c), 
            .E(n3865), .D(Y_DELTA_PATTERN[71]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i69 (.Q(Y_DELTA_PATTERN[69]), .C(ADV_CLK_c), 
            .E(n3865), .D(Y_DELTA_PATTERN[70]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_LUT4 i2_4_lut (.I0(ADV_VSYNC_c), .I1(n3549), .I2(n3855), .I3(n3859), 
            .O(n2099));
    defparam i2_4_lut.LUT_INIT = 16'heeea;
    SB_LUT4 mux_12_i9_3_lut (.I0(ADDR_Y_COMPONENT[8]), .I1(TX_ADDR[8]), 
            .I2(Y_DELTA_PATTERN[0]), .I3(GND_net), .O(n174[8]));   // ../tx.v(79[30:81])
    defparam mux_12_i9_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESR Y_DELTA_PATTERN_i68 (.Q(Y_DELTA_PATTERN[68]), .C(ADV_CLK_c), 
            .E(n3865), .D(Y_DELTA_PATTERN[69]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i67 (.Q(Y_DELTA_PATTERN[67]), .C(ADV_CLK_c), 
            .E(n3865), .D(Y_DELTA_PATTERN[68]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESR Y_DELTA_PATTERN_i66 (.Q(Y_DELTA_PATTERN[66]), .C(ADV_CLK_c), 
            .E(n3865), .D(Y_DELTA_PATTERN[67]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i65 (.Q(Y_DELTA_PATTERN[65]), .C(ADV_CLK_c), 
            .E(n3865), .D(Y_DELTA_PATTERN[66]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i64 (.Q(Y_DELTA_PATTERN[64]), .C(ADV_CLK_c), 
            .E(n3865), .D(Y_DELTA_PATTERN[65]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESR Y_DELTA_PATTERN_i63 (.Q(Y_DELTA_PATTERN[63]), .C(ADV_CLK_c), 
            .E(n3865), .D(Y_DELTA_PATTERN[64]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i62 (.Q(Y_DELTA_PATTERN[62]), .C(ADV_CLK_c), 
            .E(n3865), .D(Y_DELTA_PATTERN[63]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i61 (.Q(Y_DELTA_PATTERN[61]), .C(ADV_CLK_c), 
            .E(n3865), .D(Y_DELTA_PATTERN[62]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_CARRY add_13_8 (.CI(n3341), .I0(TX_ADDR[6]), .I1(GND_net), .CO(n3342));
    SB_DFFESR Y_DELTA_PATTERN_i60 (.Q(Y_DELTA_PATTERN[60]), .C(ADV_CLK_c), 
            .E(n3865), .D(Y_DELTA_PATTERN[61]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i59 (.Q(Y_DELTA_PATTERN[59]), .C(ADV_CLK_c), 
            .E(n3865), .D(Y_DELTA_PATTERN[60]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESR Y_DELTA_PATTERN_i58 (.Q(Y_DELTA_PATTERN[58]), .C(ADV_CLK_c), 
            .E(n3865), .D(Y_DELTA_PATTERN[59]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i57 (.Q(Y_DELTA_PATTERN[57]), .C(ADV_CLK_c), 
            .E(n3865), .D(Y_DELTA_PATTERN[58]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i56 (.Q(Y_DELTA_PATTERN[56]), .C(ADV_CLK_c), 
            .E(n3865), .D(Y_DELTA_PATTERN[57]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESR Y_DELTA_PATTERN_i55 (.Q(Y_DELTA_PATTERN[55]), .C(ADV_CLK_c), 
            .E(n3865), .D(Y_DELTA_PATTERN[56]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_LUT4 i1683_4_lut (.I0(n206[8]), .I1(ADV_VSYNC_c), .I2(n174[8]), 
            .I3(n3853), .O(n20));   // ../tx.v(68[12] 91[8])
    defparam i1683_4_lut.LUT_INIT = 16'h3022;
    SB_DFFESS X_DELTA_PATTERN_i7 (.Q(X_DELTA_PATTERN[7]), .C(ADV_CLK_c), 
            .E(n2099), .D(X_DELTA_PATTERN[8]), .S(n3864));   // ../tx.v(68[12] 91[8])
    SB_LUT4 mux_12_i10_3_lut (.I0(ADDR_Y_COMPONENT[9]), .I1(TX_ADDR[9]), 
            .I2(Y_DELTA_PATTERN[0]), .I3(GND_net), .O(n174[9]));   // ../tx.v(79[30:81])
    defparam mux_12_i10_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESS Y_DELTA_PATTERN_i54 (.Q(Y_DELTA_PATTERN[54]), .C(ADV_CLK_c), 
            .E(n3865), .D(Y_DELTA_PATTERN[55]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_LUT4 i1684_4_lut (.I0(n206[9]), .I1(ADV_VSYNC_c), .I2(n174[9]), 
            .I3(n3853), .O(n19));   // ../tx.v(68[12] 91[8])
    defparam i1684_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 add_13_7_lut (.I0(GND_net), .I1(TX_ADDR[5]), .I2(GND_net), 
            .I3(n3340), .O(n190[5])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_7 (.CI(n3340), .I0(TX_ADDR[5]), .I1(GND_net), .CO(n3341));
    SB_CARRY add_13_3 (.CI(n3336), .I0(TX_ADDR[1]), .I1(GND_net), .CO(n3337));
    SB_DFFESS Y_DELTA_PATTERN_i53 (.Q(Y_DELTA_PATTERN[53]), .C(ADV_CLK_c), 
            .E(n3865), .D(Y_DELTA_PATTERN[54]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESR Y_DELTA_PATTERN_i52 (.Q(Y_DELTA_PATTERN[52]), .C(ADV_CLK_c), 
            .E(n3865), .D(Y_DELTA_PATTERN[53]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i51 (.Q(Y_DELTA_PATTERN[51]), .C(ADV_CLK_c), 
            .E(n3865), .D(Y_DELTA_PATTERN[52]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i50 (.Q(Y_DELTA_PATTERN[50]), .C(ADV_CLK_c), 
            .E(n3865), .D(Y_DELTA_PATTERN[51]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESR Y_DELTA_PATTERN_i49 (.Q(Y_DELTA_PATTERN[49]), .C(ADV_CLK_c), 
            .E(n3865), .D(Y_DELTA_PATTERN[50]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i48 (.Q(Y_DELTA_PATTERN[48]), .C(ADV_CLK_c), 
            .E(n3865), .D(Y_DELTA_PATTERN[49]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESR Y_DELTA_PATTERN_i47 (.Q(Y_DELTA_PATTERN[47]), .C(ADV_CLK_c), 
            .E(n3865), .D(Y_DELTA_PATTERN[48]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i46 (.Q(Y_DELTA_PATTERN[46]), .C(ADV_CLK_c), 
            .E(n3865), .D(Y_DELTA_PATTERN[47]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i45 (.Q(Y_DELTA_PATTERN[45]), .C(ADV_CLK_c), 
            .E(n3865), .D(Y_DELTA_PATTERN[46]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESR Y_DELTA_PATTERN_i44 (.Q(Y_DELTA_PATTERN[44]), .C(ADV_CLK_c), 
            .E(n3865), .D(Y_DELTA_PATTERN[45]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i43 (.Q(Y_DELTA_PATTERN[43]), .C(ADV_CLK_c), 
            .E(n3865), .D(Y_DELTA_PATTERN[44]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i42 (.Q(Y_DELTA_PATTERN[42]), .C(ADV_CLK_c), 
            .E(n3865), .D(Y_DELTA_PATTERN[43]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESR Y_DELTA_PATTERN_i41 (.Q(Y_DELTA_PATTERN[41]), .C(ADV_CLK_c), 
            .E(n3865), .D(Y_DELTA_PATTERN[42]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i40 (.Q(Y_DELTA_PATTERN[40]), .C(ADV_CLK_c), 
            .E(n3865), .D(Y_DELTA_PATTERN[41]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESR Y_DELTA_PATTERN_i39 (.Q(Y_DELTA_PATTERN[39]), .C(ADV_CLK_c), 
            .E(n3865), .D(Y_DELTA_PATTERN[40]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i38 (.Q(Y_DELTA_PATTERN[38]), .C(ADV_CLK_c), 
            .E(n3865), .D(Y_DELTA_PATTERN[39]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i37 (.Q(Y_DELTA_PATTERN[37]), .C(ADV_CLK_c), 
            .E(n3865), .D(Y_DELTA_PATTERN[38]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESR Y_DELTA_PATTERN_i36 (.Q(Y_DELTA_PATTERN[36]), .C(ADV_CLK_c), 
            .E(n3865), .D(Y_DELTA_PATTERN[37]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i35 (.Q(Y_DELTA_PATTERN[35]), .C(ADV_CLK_c), 
            .E(n3865), .D(Y_DELTA_PATTERN[36]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i34 (.Q(Y_DELTA_PATTERN[34]), .C(ADV_CLK_c), 
            .E(n3865), .D(Y_DELTA_PATTERN[35]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESR Y_DELTA_PATTERN_i33 (.Q(Y_DELTA_PATTERN[33]), .C(ADV_CLK_c), 
            .E(n3865), .D(Y_DELTA_PATTERN[34]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i32 (.Q(Y_DELTA_PATTERN[32]), .C(ADV_CLK_c), 
            .E(n3864), .D(Y_DELTA_PATTERN[33]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESR Y_DELTA_PATTERN_i31 (.Q(Y_DELTA_PATTERN[31]), .C(ADV_CLK_c), 
            .E(n3864), .D(Y_DELTA_PATTERN[32]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i30 (.Q(Y_DELTA_PATTERN[30]), .C(ADV_CLK_c), 
            .E(n3864), .D(Y_DELTA_PATTERN[31]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i29 (.Q(Y_DELTA_PATTERN[29]), .C(ADV_CLK_c), 
            .E(n3864), .D(Y_DELTA_PATTERN[30]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESR Y_DELTA_PATTERN_i28 (.Q(Y_DELTA_PATTERN[28]), .C(ADV_CLK_c), 
            .E(n3864), .D(Y_DELTA_PATTERN[29]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i27 (.Q(Y_DELTA_PATTERN[27]), .C(ADV_CLK_c), 
            .E(n3864), .D(Y_DELTA_PATTERN[28]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i26 (.Q(Y_DELTA_PATTERN[26]), .C(ADV_CLK_c), 
            .E(n3864), .D(Y_DELTA_PATTERN[27]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESR Y_DELTA_PATTERN_i25 (.Q(Y_DELTA_PATTERN[25]), .C(ADV_CLK_c), 
            .E(n3864), .D(Y_DELTA_PATTERN[26]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i24 (.Q(Y_DELTA_PATTERN[24]), .C(ADV_CLK_c), 
            .E(n3864), .D(Y_DELTA_PATTERN[25]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i23 (.Q(Y_DELTA_PATTERN[23]), .C(ADV_CLK_c), 
            .E(n3864), .D(Y_DELTA_PATTERN[24]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESR Y_DELTA_PATTERN_i22 (.Q(Y_DELTA_PATTERN[22]), .C(ADV_CLK_c), 
            .E(n3864), .D(Y_DELTA_PATTERN[23]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i21 (.Q(Y_DELTA_PATTERN[21]), .C(ADV_CLK_c), 
            .E(n3864), .D(Y_DELTA_PATTERN[22]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESR Y_DELTA_PATTERN_i20 (.Q(Y_DELTA_PATTERN[20]), .C(ADV_CLK_c), 
            .E(n3864), .D(Y_DELTA_PATTERN[21]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i19 (.Q(Y_DELTA_PATTERN[19]), .C(ADV_CLK_c), 
            .E(n3864), .D(Y_DELTA_PATTERN[20]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i18 (.Q(Y_DELTA_PATTERN[18]), .C(ADV_CLK_c), 
            .E(n3864), .D(Y_DELTA_PATTERN[19]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESR Y_DELTA_PATTERN_i17 (.Q(Y_DELTA_PATTERN[17]), .C(ADV_CLK_c), 
            .E(n3864), .D(Y_DELTA_PATTERN[18]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS X_DELTA_PATTERN_i6 (.Q(X_DELTA_PATTERN[6]), .C(ADV_CLK_c), 
            .E(n2099), .D(X_DELTA_PATTERN[7]), .S(n3864));   // ../tx.v(68[12] 91[8])
    SB_DFFESR X_DELTA_PATTERN_i5 (.Q(X_DELTA_PATTERN[5]), .C(ADV_CLK_c), 
            .E(n2099), .D(X_DELTA_PATTERN[6]), .R(n3864));   // ../tx.v(68[12] 91[8])
    SB_DFFESS X_DELTA_PATTERN_i4 (.Q(X_DELTA_PATTERN[4]), .C(ADV_CLK_c), 
            .E(n2099), .D(X_DELTA_PATTERN[5]), .S(n3864));   // ../tx.v(68[12] 91[8])
    SB_DFFESR X_DELTA_PATTERN_i3 (.Q(X_DELTA_PATTERN[3]), .C(ADV_CLK_c), 
            .E(n2099), .D(X_DELTA_PATTERN[4]), .R(n3864));   // ../tx.v(68[12] 91[8])
    SB_DFFESS X_DELTA_PATTERN_i2 (.Q(X_DELTA_PATTERN[2]), .C(ADV_CLK_c), 
            .E(n2099), .D(X_DELTA_PATTERN[3]), .S(n3864));   // ../tx.v(68[12] 91[8])
    SB_LUT4 i1504_3_lut (.I0(DEBUG_c_2), .I1(BRAM_ADDR_13__N_256[13]), .I2(n2039), 
            .I3(GND_net), .O(n2775));   // ../tx.v(68[12] 91[8])
    defparam i1504_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1716_4_lut (.I0(ADV_VSYNC_c), .I1(n3852), .I2(Y_DELTA_PATTERN[0]), 
            .I3(n3853), .O(n2039));
    defparam i1716_4_lut.LUT_INIT = 16'hafee;
    SB_CARRY add_13_13 (.CI(n3346), .I0(\TX_ADDR[11] ), .I1(GND_net), 
            .CO(n3347));
    SB_LUT4 add_13_2_lut (.I0(GND_net), .I1(TX_ADDR[0]), .I2(X_DELTA_PATTERN[0]), 
            .I3(GND_net), .O(n190[0])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_2_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR X_DELTA_PATTERN_i1 (.Q(X_DELTA_PATTERN[1]), .C(ADV_CLK_c), 
            .E(n2099), .D(X_DELTA_PATTERN[2]), .R(n3864));   // ../tx.v(68[12] 91[8])
    SB_LUT4 add_13_6_lut (.I0(GND_net), .I1(TX_ADDR[4]), .I2(GND_net), 
            .I3(n3339), .O(n190[4])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_2 (.CI(GND_net), .I0(TX_ADDR[0]), .I1(X_DELTA_PATTERN[0]), 
            .CO(n3336));
    SB_LUT4 add_13_12_lut (.I0(GND_net), .I1(TX_ADDR[10]), .I2(GND_net), 
            .I3(n3345), .O(n190[10])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_12 (.CI(n3345), .I0(TX_ADDR[10]), .I1(GND_net), .CO(n3346));
    SB_CARRY add_13_6 (.CI(n3339), .I0(TX_ADDR[4]), .I1(GND_net), .CO(n3340));
    SB_LUT4 add_13_11_lut (.I0(GND_net), .I1(TX_ADDR[9]), .I2(GND_net), 
            .I3(n3344), .O(n190[9])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY add_13_11 (.CI(n3344), .I0(TX_ADDR[9]), .I1(GND_net), .CO(n3345));
    SB_LUT4 add_13_10_lut (.I0(GND_net), .I1(TX_ADDR[8]), .I2(GND_net), 
            .I3(n3343), .O(n190[8])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_10_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR ADDR_Y_COMPONENT__i0 (.Q(ADDR_Y_COMPONENT[0]), .C(ADV_CLK_c), 
            .E(n2321), .D(TX_ADDR[0]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESR BRAM_ADDR__i12 (.Q(\TX_ADDR[12] ), .C(ADV_CLK_c), .E(n2039), 
            .D(BRAM_ADDR_13__N_256[12]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESR BRAM_ADDR__rep_1_i0 (.Q(\TX_ADDR[11] ), .C(ADV_CLK_c), .E(n2039), 
            .D(BRAM_ADDR_13__N_256[11]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i0 (.Q(Y_DELTA_PATTERN[0]), .C(ADV_CLK_c), 
            .E(n3864), .D(Y_DELTA_PATTERN[1]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS X_DELTA_PATTERN_i0 (.Q(X_DELTA_PATTERN[0]), .C(ADV_CLK_c), 
            .E(n2099), .D(X_DELTA_PATTERN[1]), .S(n3864));   // ../tx.v(68[12] 91[8])
    SB_DFF BRAM_ADDR__i0 (.Q(TX_ADDR[0]), .C(ADV_CLK_c), .D(n28));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i16 (.Q(Y_DELTA_PATTERN[16]), .C(ADV_CLK_c), 
            .E(n3864), .D(Y_DELTA_PATTERN[17]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i15 (.Q(Y_DELTA_PATTERN[15]), .C(ADV_CLK_c), 
            .E(n3864), .D(Y_DELTA_PATTERN[16]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESR Y_DELTA_PATTERN_i14 (.Q(Y_DELTA_PATTERN[14]), .C(ADV_CLK_c), 
            .E(n3864), .D(Y_DELTA_PATTERN[15]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i13 (.Q(Y_DELTA_PATTERN[13]), .C(ADV_CLK_c), 
            .E(n3864), .D(Y_DELTA_PATTERN[14]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESR Y_DELTA_PATTERN_i12 (.Q(Y_DELTA_PATTERN[12]), .C(ADV_CLK_c), 
            .E(n3864), .D(Y_DELTA_PATTERN[13]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_LUT4 mux_12_i1_3_lut (.I0(ADDR_Y_COMPONENT[0]), .I1(TX_ADDR[0]), 
            .I2(Y_DELTA_PATTERN[0]), .I3(GND_net), .O(n174[0]));   // ../tx.v(79[30:81])
    defparam mux_12_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_DFFESS Y_DELTA_PATTERN_i11 (.Q(Y_DELTA_PATTERN[11]), .C(ADV_CLK_c), 
            .E(n3864), .D(Y_DELTA_PATTERN[12]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i10 (.Q(Y_DELTA_PATTERN[10]), .C(ADV_CLK_c), 
            .E(n3864), .D(Y_DELTA_PATTERN[11]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESR Y_DELTA_PATTERN_i9 (.Q(Y_DELTA_PATTERN[9]), .C(ADV_CLK_c), 
            .E(n3864), .D(Y_DELTA_PATTERN[10]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i8 (.Q(Y_DELTA_PATTERN[8]), .C(ADV_CLK_c), 
            .E(n3864), .D(Y_DELTA_PATTERN[9]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i7 (.Q(Y_DELTA_PATTERN[7]), .C(ADV_CLK_c), 
            .E(n3864), .D(Y_DELTA_PATTERN[8]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_CARRY add_13_10 (.CI(n3343), .I0(TX_ADDR[8]), .I1(GND_net), .CO(n3344));
    SB_DFFESR Y_DELTA_PATTERN_i6 (.Q(Y_DELTA_PATTERN[6]), .C(ADV_CLK_c), 
            .E(n3864), .D(Y_DELTA_PATTERN[7]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i5 (.Q(Y_DELTA_PATTERN[5]), .C(ADV_CLK_c), 
            .E(n3864), .D(Y_DELTA_PATTERN[6]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESR Y_DELTA_PATTERN_i4 (.Q(Y_DELTA_PATTERN[4]), .C(ADV_CLK_c), 
            .E(n3864), .D(Y_DELTA_PATTERN[5]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESS Y_DELTA_PATTERN_i3 (.Q(Y_DELTA_PATTERN[3]), .C(ADV_CLK_c), 
            .E(n3864), .D(Y_DELTA_PATTERN[4]), .S(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESR ADDR_Y_COMPONENT__i13 (.Q(ADDR_Y_COMPONENT[13]), .C(ADV_CLK_c), 
            .E(n2321), .D(DEBUG_c_2), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_LUT4 add_13_5_lut (.I0(GND_net), .I1(TX_ADDR[3]), .I2(GND_net), 
            .I3(n3338), .O(n190[3])) /* synthesis syn_instantiated=1 */ ;
    defparam add_13_5_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i1670_4_lut (.I0(n206[0]), .I1(ADV_VSYNC_c), .I2(n174[0]), 
            .I3(n3853), .O(n28));   // ../tx.v(68[12] 91[8])
    defparam i1670_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 mux_12_i2_3_lut (.I0(ADDR_Y_COMPONENT[1]), .I1(TX_ADDR[1]), 
            .I2(Y_DELTA_PATTERN[0]), .I3(GND_net), .O(n174[1]));   // ../tx.v(79[30:81])
    defparam mux_12_i2_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1676_4_lut (.I0(n206[1]), .I1(ADV_VSYNC_c), .I2(n174[1]), 
            .I3(n3853), .O(n27));   // ../tx.v(68[12] 91[8])
    defparam i1676_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 mux_12_i3_3_lut (.I0(ADDR_Y_COMPONENT[2]), .I1(TX_ADDR[2]), 
            .I2(Y_DELTA_PATTERN[0]), .I3(GND_net), .O(n174[2]));   // ../tx.v(79[30:81])
    defparam mux_12_i3_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1677_4_lut (.I0(n206[2]), .I1(ADV_VSYNC_c), .I2(n174[2]), 
            .I3(n3853), .O(n26));   // ../tx.v(68[12] 91[8])
    defparam i1677_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 mux_12_i4_3_lut (.I0(ADDR_Y_COMPONENT[3]), .I1(TX_ADDR[3]), 
            .I2(Y_DELTA_PATTERN[0]), .I3(GND_net), .O(n174[3]));   // ../tx.v(79[30:81])
    defparam mux_12_i4_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1678_4_lut (.I0(n206[3]), .I1(ADV_VSYNC_c), .I2(n174[3]), 
            .I3(n3853), .O(n25));   // ../tx.v(68[12] 91[8])
    defparam i1678_4_lut.LUT_INIT = 16'h3022;
    SB_LUT4 mux_12_i5_3_lut (.I0(ADDR_Y_COMPONENT[4]), .I1(TX_ADDR[4]), 
            .I2(Y_DELTA_PATTERN[0]), .I3(GND_net), .O(n174[4]));   // ../tx.v(79[30:81])
    defparam mux_12_i5_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1679_4_lut (.I0(n206[4]), .I1(ADV_VSYNC_c), .I2(n174[4]), 
            .I3(n3853), .O(n24));   // ../tx.v(68[12] 91[8])
    defparam i1679_4_lut.LUT_INIT = 16'h3022;
    SB_DFFSR BRAM_ADDR__i13 (.Q(DEBUG_c_2), .C(ADV_CLK_c), .D(n2775), 
            .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESR ADDR_Y_COMPONENT__i12 (.Q(ADDR_Y_COMPONENT[12]), .C(ADV_CLK_c), 
            .E(n2321), .D(\TX_ADDR[12] ), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESR ADDR_Y_COMPONENT__i11 (.Q(ADDR_Y_COMPONENT[11]), .C(ADV_CLK_c), 
            .E(n2321), .D(\TX_ADDR[11] ), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESR ADDR_Y_COMPONENT__i10 (.Q(ADDR_Y_COMPONENT[10]), .C(ADV_CLK_c), 
            .E(n2321), .D(TX_ADDR[10]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESR ADDR_Y_COMPONENT__i9 (.Q(ADDR_Y_COMPONENT[9]), .C(ADV_CLK_c), 
            .E(n2321), .D(TX_ADDR[9]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESR ADDR_Y_COMPONENT__i8 (.Q(ADDR_Y_COMPONENT[8]), .C(ADV_CLK_c), 
            .E(n2321), .D(TX_ADDR[8]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESR ADDR_Y_COMPONENT__i7 (.Q(ADDR_Y_COMPONENT[7]), .C(ADV_CLK_c), 
            .E(n2321), .D(TX_ADDR[7]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESR ADDR_Y_COMPONENT__i6 (.Q(ADDR_Y_COMPONENT[6]), .C(ADV_CLK_c), 
            .E(n2321), .D(TX_ADDR[6]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESR ADDR_Y_COMPONENT__i5 (.Q(ADDR_Y_COMPONENT[5]), .C(ADV_CLK_c), 
            .E(n2321), .D(TX_ADDR[5]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESR ADDR_Y_COMPONENT__i1 (.Q(ADDR_Y_COMPONENT[1]), .C(ADV_CLK_c), 
            .E(n2321), .D(TX_ADDR[1]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESR ADDR_Y_COMPONENT__i4 (.Q(ADDR_Y_COMPONENT[4]), .C(ADV_CLK_c), 
            .E(n2321), .D(TX_ADDR[4]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    SB_DFFESR ADDR_Y_COMPONENT__i2 (.Q(ADDR_Y_COMPONENT[2]), .C(ADV_CLK_c), 
            .E(n2321), .D(TX_ADDR[2]), .R(ADV_VSYNC_c));   // ../tx.v(68[12] 91[8])
    VGA_CONTROL video_signal_controller (.ADV_CLK_c(ADV_CLK_c), .GND_net(GND_net), 
            .VCC_net(VCC_net), .ADV_HSYNC_c(ADV_HSYNC_c), .ADV_VSYNC_c(ADV_VSYNC_c), 
            .DEBUG_c_6(DEBUG_c_6), .n3855(n3855), .n3549(n3549), .n190({n190}), 
            .\TX_ADDR[6] (TX_ADDR[6]), .n214(n206[6]), .\TX_ADDR[5] (TX_ADDR[5]), 
            .n215(n206[5]), .n3859(n3859), .\ADDR_Y_COMPONENT[12] (ADDR_Y_COMPONENT[12]), 
            .\BRAM_ADDR_13__N_256[12] (BRAM_ADDR_13__N_256[12]), .\Y_DELTA_PATTERN[0] (Y_DELTA_PATTERN[0]), 
            .n2321(n2321), .old_VGA_HS(old_VGA_HS), .n2125(n2125), .n3853(n3853), 
            .\ADDR_Y_COMPONENT[11] (ADDR_Y_COMPONENT[11]), .\BRAM_ADDR_13__N_256[11] (BRAM_ADDR_13__N_256[11]), 
            .\ADDR_Y_COMPONENT[13] (ADDR_Y_COMPONENT[13]), .\BRAM_ADDR_13__N_256[13] (BRAM_ADDR_13__N_256[13]), 
            .\TX_ADDR[0] (TX_ADDR[0]), .n220(n206[0]), .\TX_ADDR[1] (TX_ADDR[1]), 
            .n219(n206[1]), .\TX_ADDR[2] (TX_ADDR[2]), .n218(n206[2]), 
            .\TX_ADDR[3] (TX_ADDR[3]), .n217(n206[3]), .\TX_ADDR[10] (TX_ADDR[10]), 
            .n210(n206[10]), .n2404(n2404), .n3852(n3852), .\TX_ADDR[8] (TX_ADDR[8]), 
            .n212(n206[8]), .\TX_ADDR[9] (TX_ADDR[9]), .n211(n206[9]), 
            .\TX_ADDR[7] (TX_ADDR[7]), .n213(n206[7]), .n3865(n3865), 
            .n3864(n3864), .\TX_ADDR[4] (TX_ADDR[4]), .n216(n206[4])) /* synthesis syn_module_defined=1 */ ;   // ../tx.v(42[17] 56[67])
    
endmodule
//
// Verilog Description of module VGA_CONTROL
//

module VGA_CONTROL (ADV_CLK_c, GND_net, VCC_net, ADV_HSYNC_c, ADV_VSYNC_c, 
            DEBUG_c_6, n3855, n3549, n190, \TX_ADDR[6] , n214, \TX_ADDR[5] , 
            n215, n3859, \ADDR_Y_COMPONENT[12] , \BRAM_ADDR_13__N_256[12] , 
            \Y_DELTA_PATTERN[0] , n2321, old_VGA_HS, n2125, n3853, 
            \ADDR_Y_COMPONENT[11] , \BRAM_ADDR_13__N_256[11] , \ADDR_Y_COMPONENT[13] , 
            \BRAM_ADDR_13__N_256[13] , \TX_ADDR[0] , n220, \TX_ADDR[1] , 
            n219, \TX_ADDR[2] , n218, \TX_ADDR[3] , n217, \TX_ADDR[10] , 
            n210, n2404, n3852, \TX_ADDR[8] , n212, \TX_ADDR[9] , 
            n211, \TX_ADDR[7] , n213, n3865, n3864, \TX_ADDR[4] , 
            n216) /* synthesis syn_module_defined=1 */ ;
    input ADV_CLK_c;
    input GND_net;
    input VCC_net;
    output ADV_HSYNC_c;
    output ADV_VSYNC_c;
    input DEBUG_c_6;
    output n3855;
    output n3549;
    input [13:0]n190;
    input \TX_ADDR[6] ;
    output n214;
    input \TX_ADDR[5] ;
    output n215;
    output n3859;
    input \ADDR_Y_COMPONENT[12] ;
    output \BRAM_ADDR_13__N_256[12] ;
    input \Y_DELTA_PATTERN[0] ;
    output n2321;
    input old_VGA_HS;
    output n2125;
    output n3853;
    input \ADDR_Y_COMPONENT[11] ;
    output \BRAM_ADDR_13__N_256[11] ;
    input \ADDR_Y_COMPONENT[13] ;
    output \BRAM_ADDR_13__N_256[13] ;
    input \TX_ADDR[0] ;
    output n220;
    input \TX_ADDR[1] ;
    output n219;
    input \TX_ADDR[2] ;
    output n218;
    input \TX_ADDR[3] ;
    output n217;
    input \TX_ADDR[10] ;
    output n210;
    output n2404;
    output n3852;
    input \TX_ADDR[8] ;
    output n212;
    input \TX_ADDR[9] ;
    output n211;
    input \TX_ADDR[7] ;
    output n213;
    output n3865;
    output n3864;
    input \TX_ADDR[4] ;
    output n216;
    
    wire ADV_CLK_c /* synthesis SET_AS_NETWORK=ADV_CLK_c, is_clock=1 */ ;   // ../main.v(13[14:21])
    wire [11:0]n1;
    
    wire n2030;
    wire [11:0]VGA_Y;   // ../vga_control.v(54[23:28])
    
    wire n2551;
    wire [10:0]n49;
    wire [11:0]VGA_X;   // ../vga_control.v(54[16:21])
    
    wire n3379, n3380, n3378, n3377, n3376, SYNC_BUFF1, SYNC_BUFF2, 
        n3381, n3375, n3385, VGA_HS_N_543, VGA_VS_N_546, n3386, 
        n3374, n3373, n3372, n3371, n3370, n3575, n6, n2015, 
        n3369, n3368, n3367, n3384, n3023, n3383, n8, n3382, 
        n3366, n3577, n3858, n6_adj_568, n3697, n21, n3603, n4, 
        n23, n8_adj_569, n3857, n3029, n3856;
    
    SB_DFFESR VGA_Y_265__i10 (.Q(VGA_Y[10]), .C(ADV_CLK_c), .E(n2030), 
            .D(n1[10]), .R(n2551));   // ../vga_control.v(91[30:39])
    SB_DFFESR VGA_Y_265__i9 (.Q(VGA_Y[9]), .C(ADV_CLK_c), .E(n2030), .D(n1[9]), 
            .R(n2551));   // ../vga_control.v(91[30:39])
    SB_LUT4 VGA_X_266_267_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(VGA_X[3]), 
            .I3(n3379), .O(n49[3])) /* synthesis syn_instantiated=1 */ ;
    defparam VGA_X_266_267_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR VGA_Y_265__i8 (.Q(VGA_Y[8]), .C(ADV_CLK_c), .E(n2030), .D(n1[8]), 
            .R(n2551));   // ../vga_control.v(91[30:39])
    SB_DFFESR VGA_Y_265__i7 (.Q(VGA_Y[7]), .C(ADV_CLK_c), .E(n2030), .D(n1[7]), 
            .R(n2551));   // ../vga_control.v(91[30:39])
    SB_DFFESR VGA_Y_265__i6 (.Q(VGA_Y[6]), .C(ADV_CLK_c), .E(n2030), .D(n1[6]), 
            .R(n2551));   // ../vga_control.v(91[30:39])
    SB_DFFESR VGA_Y_265__i5 (.Q(VGA_Y[5]), .C(ADV_CLK_c), .E(n2030), .D(n1[5]), 
            .R(n2551));   // ../vga_control.v(91[30:39])
    SB_DFFESR VGA_Y_265__i4 (.Q(VGA_Y[4]), .C(ADV_CLK_c), .E(n2030), .D(n1[4]), 
            .R(n2551));   // ../vga_control.v(91[30:39])
    SB_DFFESR VGA_Y_265__i3 (.Q(VGA_Y[3]), .C(ADV_CLK_c), .E(n2030), .D(n1[3]), 
            .R(n2551));   // ../vga_control.v(91[30:39])
    SB_DFFSR VGA_X_266_267__i1 (.Q(VGA_X[0]), .C(ADV_CLK_c), .D(n49[0]), 
            .R(n2030));   // ../vga_control.v(85[26:35])
    SB_DFFESR VGA_Y_265__i2 (.Q(VGA_Y[2]), .C(ADV_CLK_c), .E(n2030), .D(n1[2]), 
            .R(n2551));   // ../vga_control.v(91[30:39])
    SB_CARRY VGA_X_266_267_add_4_5 (.CI(n3379), .I0(GND_net), .I1(VGA_X[3]), 
            .CO(n3380));
    SB_DFFESR VGA_Y_265__i1 (.Q(VGA_Y[1]), .C(ADV_CLK_c), .E(n2030), .D(n1[1]), 
            .R(n2551));   // ../vga_control.v(91[30:39])
    SB_LUT4 VGA_X_266_267_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(VGA_X[2]), 
            .I3(n3378), .O(n49[2])) /* synthesis syn_instantiated=1 */ ;
    defparam VGA_X_266_267_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY VGA_X_266_267_add_4_4 (.CI(n3378), .I0(GND_net), .I1(VGA_X[2]), 
            .CO(n3379));
    SB_LUT4 VGA_X_266_267_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(VGA_X[1]), 
            .I3(n3377), .O(n49[1])) /* synthesis syn_instantiated=1 */ ;
    defparam VGA_X_266_267_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY VGA_X_266_267_add_4_3 (.CI(n3377), .I0(GND_net), .I1(VGA_X[1]), 
            .CO(n3378));
    SB_LUT4 VGA_X_266_267_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(VGA_X[0]), 
            .I3(VCC_net), .O(n49[0])) /* synthesis syn_instantiated=1 */ ;
    defparam VGA_X_266_267_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY VGA_X_266_267_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(VGA_X[0]), 
            .CO(n3377));
    SB_LUT4 VGA_Y_265_add_4_13_lut (.I0(GND_net), .I1(GND_net), .I2(VGA_Y[11]), 
            .I3(n3376), .O(n1[11])) /* synthesis syn_instantiated=1 */ ;
    defparam VGA_Y_265_add_4_13_lut.LUT_INIT = 16'hC33C;
    SB_DFF SYNC_BUFF2_52 (.Q(SYNC_BUFF2), .C(ADV_CLK_c), .D(SYNC_BUFF1));   // ../vga_control.v(73[12] 100[8])
    SB_CARRY VGA_X_266_267_add_4_6 (.CI(n3380), .I0(GND_net), .I1(VGA_X[4]), 
            .CO(n3381));
    SB_LUT4 VGA_Y_265_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(VGA_Y[10]), 
            .I3(n3375), .O(n1[10])) /* synthesis syn_instantiated=1 */ ;
    defparam VGA_Y_265_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_CARRY VGA_Y_265_add_4_12 (.CI(n3375), .I0(GND_net), .I1(VGA_Y[10]), 
            .CO(n3376));
    SB_LUT4 VGA_X_266_267_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(VGA_X[9]), 
            .I3(n3385), .O(n49[9])) /* synthesis syn_instantiated=1 */ ;
    defparam VGA_X_266_267_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_DFF VGA_HS_54 (.Q(ADV_HSYNC_c), .C(ADV_CLK_c), .D(VGA_HS_N_543));   // ../vga_control.v(73[12] 100[8])
    SB_DFF VGA_VS_55 (.Q(ADV_VSYNC_c), .C(ADV_CLK_c), .D(VGA_VS_N_546));   // ../vga_control.v(73[12] 100[8])
    SB_DFF SYNC_BUFF1_51 (.Q(SYNC_BUFF1), .C(ADV_CLK_c), .D(DEBUG_c_6));   // ../vga_control.v(73[12] 100[8])
    SB_LUT4 VGA_X_266_267_add_4_12_lut (.I0(GND_net), .I1(GND_net), .I2(VGA_X[10]), 
            .I3(n3386), .O(n49[10])) /* synthesis syn_instantiated=1 */ ;
    defparam VGA_X_266_267_add_4_12_lut.LUT_INIT = 16'hC33C;
    SB_DFFESR VGA_Y_265__i11 (.Q(VGA_Y[11]), .C(ADV_CLK_c), .E(n2030), 
            .D(n1[11]), .R(n2551));   // ../vga_control.v(91[30:39])
    SB_LUT4 VGA_Y_265_add_4_11_lut (.I0(GND_net), .I1(GND_net), .I2(VGA_Y[9]), 
            .I3(n3374), .O(n1[9])) /* synthesis syn_instantiated=1 */ ;
    defparam VGA_Y_265_add_4_11_lut.LUT_INIT = 16'hC33C;
    SB_CARRY VGA_Y_265_add_4_11 (.CI(n3374), .I0(GND_net), .I1(VGA_Y[9]), 
            .CO(n3375));
    SB_LUT4 VGA_Y_265_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(VGA_Y[8]), 
            .I3(n3373), .O(n1[8])) /* synthesis syn_instantiated=1 */ ;
    defparam VGA_Y_265_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 mux_15_i7_3_lut_4_lut (.I0(n3855), .I1(n3549), .I2(n190[6]), 
            .I3(\TX_ADDR[6] ), .O(n214));   // ../vga_control.v(57[28:124])
    defparam mux_15_i7_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_CARRY VGA_Y_265_add_4_10 (.CI(n3373), .I0(GND_net), .I1(VGA_Y[8]), 
            .CO(n3374));
    SB_LUT4 VGA_Y_265_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(VGA_Y[7]), 
            .I3(n3372), .O(n1[7])) /* synthesis syn_instantiated=1 */ ;
    defparam VGA_Y_265_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY VGA_Y_265_add_4_9 (.CI(n3372), .I0(GND_net), .I1(VGA_Y[7]), 
            .CO(n3373));
    SB_LUT4 VGA_Y_265_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(VGA_Y[6]), 
            .I3(n3371), .O(n1[6])) /* synthesis syn_instantiated=1 */ ;
    defparam VGA_Y_265_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY VGA_Y_265_add_4_8 (.CI(n3371), .I0(GND_net), .I1(VGA_Y[6]), 
            .CO(n3372));
    SB_LUT4 VGA_Y_265_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(VGA_Y[5]), 
            .I3(n3370), .O(n1[5])) /* synthesis syn_instantiated=1 */ ;
    defparam VGA_Y_265_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 i4_4_lut (.I0(VGA_Y[5]), .I1(VGA_Y[9]), .I2(n3575), .I3(n6), 
            .O(n2015));
    defparam i4_4_lut.LUT_INIT = 16'hfffe;
    SB_CARRY VGA_Y_265_add_4_7 (.CI(n3370), .I0(GND_net), .I1(VGA_Y[5]), 
            .CO(n3371));
    SB_LUT4 VGA_Y_265_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(VGA_Y[4]), 
            .I3(n3369), .O(n1[4])) /* synthesis syn_instantiated=1 */ ;
    defparam VGA_Y_265_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_CARRY VGA_Y_265_add_4_6 (.CI(n3369), .I0(GND_net), .I1(VGA_Y[4]), 
            .CO(n3370));
    SB_LUT4 VGA_Y_265_add_4_5_lut (.I0(GND_net), .I1(GND_net), .I2(VGA_Y[3]), 
            .I3(n3368), .O(n1[3])) /* synthesis syn_instantiated=1 */ ;
    defparam VGA_Y_265_add_4_5_lut.LUT_INIT = 16'hC33C;
    SB_CARRY VGA_Y_265_add_4_5 (.CI(n3368), .I0(GND_net), .I1(VGA_Y[3]), 
            .CO(n3369));
    SB_LUT4 VGA_Y_265_add_4_4_lut (.I0(GND_net), .I1(GND_net), .I2(VGA_Y[2]), 
            .I3(n3367), .O(n1[2])) /* synthesis syn_instantiated=1 */ ;
    defparam VGA_Y_265_add_4_4_lut.LUT_INIT = 16'hC33C;
    SB_CARRY VGA_Y_265_add_4_4 (.CI(n3367), .I0(GND_net), .I1(VGA_Y[2]), 
            .CO(n3368));
    SB_CARRY VGA_X_266_267_add_4_11 (.CI(n3385), .I0(GND_net), .I1(VGA_X[9]), 
            .CO(n3386));
    SB_LUT4 VGA_X_266_267_add_4_10_lut (.I0(GND_net), .I1(GND_net), .I2(VGA_X[8]), 
            .I3(n3384), .O(n49[8])) /* synthesis syn_instantiated=1 */ ;
    defparam VGA_X_266_267_add_4_10_lut.LUT_INIT = 16'hC33C;
    SB_CARRY VGA_X_266_267_add_4_10 (.CI(n3384), .I0(GND_net), .I1(VGA_X[8]), 
            .CO(n3385));
    SB_LUT4 i1_2_lut (.I0(VGA_Y[7]), .I1(VGA_Y[8]), .I2(GND_net), .I3(GND_net), 
            .O(n3575));
    defparam i1_2_lut.LUT_INIT = 16'heeee;
    SB_LUT4 i1753_4_lut (.I0(VGA_Y[2]), .I1(VGA_Y[4]), .I2(VGA_Y[3]), 
            .I3(VGA_Y[1]), .O(n3023));
    defparam i1753_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 VGA_X_266_267_add_4_9_lut (.I0(GND_net), .I1(GND_net), .I2(VGA_X[7]), 
            .I3(n3383), .O(n49[7])) /* synthesis syn_instantiated=1 */ ;
    defparam VGA_X_266_267_add_4_9_lut.LUT_INIT = 16'hC33C;
    SB_CARRY VGA_X_266_267_add_4_9 (.CI(n3383), .I0(GND_net), .I1(VGA_X[7]), 
            .CO(n3384));
    SB_LUT4 i487_3_lut (.I0(VGA_Y[1]), .I1(VGA_Y[3]), .I2(VGA_Y[2]), .I3(GND_net), 
            .O(n8));
    defparam i487_3_lut.LUT_INIT = 16'hecec;
    SB_LUT4 VGA_X_266_267_add_4_8_lut (.I0(GND_net), .I1(GND_net), .I2(VGA_X[6]), 
            .I3(n3382), .O(n49[6])) /* synthesis syn_instantiated=1 */ ;
    defparam VGA_X_266_267_add_4_8_lut.LUT_INIT = 16'hC33C;
    SB_CARRY VGA_X_266_267_add_4_8 (.CI(n3382), .I0(GND_net), .I1(VGA_X[6]), 
            .CO(n3383));
    SB_LUT4 VGA_X_266_267_add_4_7_lut (.I0(GND_net), .I1(GND_net), .I2(VGA_X[5]), 
            .I3(n3381), .O(n49[5])) /* synthesis syn_instantiated=1 */ ;
    defparam VGA_X_266_267_add_4_7_lut.LUT_INIT = 16'hC33C;
    SB_CARRY VGA_X_266_267_add_4_7 (.CI(n3381), .I0(GND_net), .I1(VGA_X[5]), 
            .CO(n3382));
    SB_LUT4 VGA_X_266_267_add_4_6_lut (.I0(GND_net), .I1(GND_net), .I2(VGA_X[4]), 
            .I3(n3380), .O(n49[4])) /* synthesis syn_instantiated=1 */ ;
    defparam VGA_X_266_267_add_4_6_lut.LUT_INIT = 16'hC33C;
    SB_LUT4 VGA_Y_265_add_4_3_lut (.I0(GND_net), .I1(GND_net), .I2(VGA_Y[1]), 
            .I3(n3366), .O(n1[1])) /* synthesis syn_instantiated=1 */ ;
    defparam VGA_Y_265_add_4_3_lut.LUT_INIT = 16'hC33C;
    SB_CARRY VGA_Y_265_add_4_3 (.CI(n3366), .I0(GND_net), .I1(VGA_Y[1]), 
            .CO(n3367));
    SB_LUT4 VGA_Y_265_add_4_2_lut (.I0(GND_net), .I1(GND_net), .I2(VGA_Y[0]), 
            .I3(VCC_net), .O(n1[0])) /* synthesis syn_instantiated=1 */ ;
    defparam VGA_Y_265_add_4_2_lut.LUT_INIT = 16'hC33C;
    SB_CARRY VGA_Y_265_add_4_2 (.CI(VCC_net), .I0(GND_net), .I1(VGA_Y[0]), 
            .CO(n3366));
    SB_LUT4 i1_4_lut (.I0(VGA_Y[5]), .I1(n3575), .I2(VGA_Y[6]), .I3(n3023), 
            .O(n3577));
    defparam i1_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i2_4_lut (.I0(n8), .I1(n3858), .I2(n2015), .I3(VGA_Y[4]), 
            .O(n6_adj_568));
    defparam i2_4_lut.LUT_INIT = 16'h3230;
    SB_LUT4 i2335_3_lut (.I0(VGA_Y[4]), .I1(n2015), .I2(VGA_Y[3]), .I3(GND_net), 
            .O(n3697));
    defparam i2335_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i4_4_lut_adj_13 (.I0(VGA_Y[0]), .I1(n3697), .I2(VGA_Y[2]), 
            .I3(VGA_Y[1]), .O(VGA_VS_N_546));
    defparam i4_4_lut_adj_13.LUT_INIT = 16'h0302;
    SB_LUT4 i1_3_lut (.I0(VGA_X[5]), .I1(VGA_X[3]), .I2(VGA_X[4]), .I3(GND_net), 
            .O(n21));
    defparam i1_3_lut.LUT_INIT = 16'ha8a8;
    SB_LUT4 i3_4_lut (.I0(n3603), .I1(n6_adj_568), .I2(n3577), .I3(VGA_Y[9]), 
            .O(n3549));
    defparam i3_4_lut.LUT_INIT = 16'h0444;
    SB_LUT4 i1_2_lut_adj_14 (.I0(VGA_X[4]), .I1(VGA_X[5]), .I2(GND_net), 
            .I3(GND_net), .O(n4));
    defparam i1_2_lut_adj_14.LUT_INIT = 16'heeee;
    SB_LUT4 i37_4_lut (.I0(VGA_X[6]), .I1(n4), .I2(VGA_X[7]), .I3(n21), 
            .O(n23));
    defparam i37_4_lut.LUT_INIT = 16'h1f1a;
    SB_DFFSR VGA_X_266_267__i2 (.Q(VGA_X[1]), .C(ADV_CLK_c), .D(n49[1]), 
            .R(n2030));   // ../vga_control.v(85[26:35])
    SB_DFFSR VGA_X_266_267__i3 (.Q(VGA_X[2]), .C(ADV_CLK_c), .D(n49[2]), 
            .R(n2030));   // ../vga_control.v(85[26:35])
    SB_DFFSR VGA_X_266_267__i4 (.Q(VGA_X[3]), .C(ADV_CLK_c), .D(n49[3]), 
            .R(n2030));   // ../vga_control.v(85[26:35])
    SB_DFFSR VGA_X_266_267__i5 (.Q(VGA_X[4]), .C(ADV_CLK_c), .D(n49[4]), 
            .R(n2030));   // ../vga_control.v(85[26:35])
    SB_DFFSR VGA_X_266_267__i6 (.Q(VGA_X[5]), .C(ADV_CLK_c), .D(n49[5]), 
            .R(n2030));   // ../vga_control.v(85[26:35])
    SB_DFFSR VGA_X_266_267__i7 (.Q(VGA_X[6]), .C(ADV_CLK_c), .D(n49[6]), 
            .R(n2030));   // ../vga_control.v(85[26:35])
    SB_DFFSR VGA_X_266_267__i8 (.Q(VGA_X[7]), .C(ADV_CLK_c), .D(n49[7]), 
            .R(n2030));   // ../vga_control.v(85[26:35])
    SB_DFFSR VGA_X_266_267__i9 (.Q(VGA_X[8]), .C(ADV_CLK_c), .D(n49[8]), 
            .R(n2030));   // ../vga_control.v(85[26:35])
    SB_DFFSR VGA_X_266_267__i10 (.Q(VGA_X[9]), .C(ADV_CLK_c), .D(n49[9]), 
            .R(n2030));   // ../vga_control.v(85[26:35])
    SB_DFFSR VGA_X_266_267__i11 (.Q(VGA_X[10]), .C(ADV_CLK_c), .D(n49[10]), 
            .R(n2030));   // ../vga_control.v(85[26:35])
    SB_LUT4 mux_15_i6_3_lut_4_lut (.I0(n3855), .I1(n3549), .I2(n190[5]), 
            .I3(\TX_ADDR[5] ), .O(n215));   // ../vga_control.v(57[28:124])
    defparam mux_15_i6_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1078_3_lut_4_lut (.I0(n3549), .I1(n3859), .I2(\ADDR_Y_COMPONENT[12] ), 
            .I3(n190[12]), .O(\BRAM_ADDR_13__N_256[12] ));   // ../vga_control.v(57[28:124])
    defparam i1078_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_3_lut_4_lut (.I0(n3549), .I1(n3859), .I2(\Y_DELTA_PATTERN[0] ), 
            .I3(ADV_VSYNC_c), .O(n2321));   // ../vga_control.v(57[28:124])
    defparam i1_3_lut_4_lut.LUT_INIT = 16'hff80;
    SB_DFFESR VGA_Y_265__i0 (.Q(VGA_Y[0]), .C(ADV_CLK_c), .E(n2030), .D(n1[0]), 
            .R(n2551));   // ../vga_control.v(91[30:39])
    SB_LUT4 i271_2_lut_3_lut_4_lut (.I0(ADV_HSYNC_c), .I1(old_VGA_HS), .I2(ADV_VSYNC_c), 
            .I3(n3549), .O(n2125));   // ../vga_control.v(57[28:124])
    defparam i271_2_lut_3_lut_4_lut.LUT_INIT = 16'hf4f0;
    SB_LUT4 i1_2_lut_rep_17_3_lut (.I0(ADV_HSYNC_c), .I1(old_VGA_HS), .I2(n3549), 
            .I3(GND_net), .O(n3853));   // ../vga_control.v(57[28:124])
    defparam i1_2_lut_rep_17_3_lut.LUT_INIT = 16'h4040;
    SB_LUT4 i1289_2_lut (.I0(n2030), .I1(SYNC_BUFF2), .I2(GND_net), .I3(GND_net), 
            .O(n2551));   // ../vga_control.v(91[30:39])
    defparam i1289_2_lut.LUT_INIT = 16'h8888;
    SB_LUT4 i3_3_lut (.I0(VGA_X[1]), .I1(VGA_X[3]), .I2(VGA_X[2]), .I3(GND_net), 
            .O(n8_adj_569));
    defparam i3_3_lut.LUT_INIT = 16'h8080;
    SB_LUT4 i1_2_lut_rep_23 (.I0(ADV_HSYNC_c), .I1(old_VGA_HS), .I2(GND_net), 
            .I3(GND_net), .O(n3859));   // ../vga_control.v(57[28:124])
    defparam i1_2_lut_rep_23.LUT_INIT = 16'h4444;
    SB_LUT4 i1759_4_lut (.I0(VGA_X[0]), .I1(n3857), .I2(n8_adj_569), .I3(VGA_X[4]), 
            .O(n3029));
    defparam i1759_4_lut.LUT_INIT = 16'heccc;
    SB_LUT4 i1_2_lut_3_lut (.I0(VGA_Y[10]), .I1(VGA_Y[11]), .I2(VGA_Y[6]), 
            .I3(GND_net), .O(n6));
    defparam i1_2_lut_3_lut.LUT_INIT = 16'hfefe;
    SB_LUT4 i1080_3_lut_4_lut (.I0(n3549), .I1(n3859), .I2(\ADDR_Y_COMPONENT[11] ), 
            .I3(n190[11]), .O(\BRAM_ADDR_13__N_256[11] ));   // ../vga_control.v(57[28:124])
    defparam i1080_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1076_3_lut_4_lut (.I0(n3549), .I1(n3859), .I2(\ADDR_Y_COMPONENT[13] ), 
            .I3(n190[13]), .O(\BRAM_ADDR_13__N_256[13] ));   // ../vga_control.v(57[28:124])
    defparam i1076_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1_2_lut_rep_22 (.I0(VGA_Y[10]), .I1(VGA_Y[11]), .I2(GND_net), 
            .I3(GND_net), .O(n3858));
    defparam i1_2_lut_rep_22.LUT_INIT = 16'heeee;
    SB_LUT4 mux_15_i1_3_lut_4_lut (.I0(n3855), .I1(n3549), .I2(n190[0]), 
            .I3(\TX_ADDR[0] ), .O(n220));   // ../vga_control.v(57[28:124])
    defparam mux_15_i1_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 mux_15_i2_3_lut_4_lut (.I0(n3855), .I1(n3549), .I2(n190[1]), 
            .I3(\TX_ADDR[1] ), .O(n219));   // ../vga_control.v(57[28:124])
    defparam mux_15_i2_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 mux_15_i3_3_lut_4_lut (.I0(n3855), .I1(n3549), .I2(n190[2]), 
            .I3(\TX_ADDR[2] ), .O(n218));   // ../vga_control.v(57[28:124])
    defparam mux_15_i3_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 mux_15_i4_3_lut_4_lut (.I0(n3855), .I1(n3549), .I2(n190[3]), 
            .I3(\TX_ADDR[3] ), .O(n217));   // ../vga_control.v(57[28:124])
    defparam mux_15_i4_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i2_3_lut_rep_21 (.I0(VGA_X[6]), .I1(VGA_X[5]), .I2(VGA_X[7]), 
            .I3(GND_net), .O(n3857));
    defparam i2_3_lut_rep_21.LUT_INIT = 16'hfefe;
    SB_LUT4 i2387_3_lut_4_lut (.I0(VGA_X[9]), .I1(VGA_X[10]), .I2(VGA_X[8]), 
            .I3(n23), .O(VGA_HS_N_543));
    defparam i2387_3_lut_4_lut.LUT_INIT = 16'hfeff;
    SB_LUT4 i1_2_lut_rep_19_3_lut_4_lut (.I0(VGA_X[9]), .I1(VGA_X[10]), 
            .I2(VGA_X[8]), .I3(n3857), .O(n3855));
    defparam i1_2_lut_rep_19_3_lut_4_lut.LUT_INIT = 16'hfeee;
    SB_LUT4 i1_2_lut_rep_20 (.I0(VGA_X[9]), .I1(VGA_X[10]), .I2(GND_net), 
            .I3(GND_net), .O(n3856));
    defparam i1_2_lut_rep_20.LUT_INIT = 16'heeee;
    SB_LUT4 mux_15_i11_3_lut_4_lut (.I0(n3855), .I1(n3549), .I2(n190[10]), 
            .I3(\TX_ADDR[10] ), .O(n210));   // ../vga_control.v(57[28:124])
    defparam mux_15_i11_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1133_1_lut_2_lut_3_lut_4_lut (.I0(n3857), .I1(VGA_X[8]), .I2(n3549), 
            .I3(n3856), .O(n2404));
    defparam i1133_1_lut_2_lut_3_lut_4_lut.LUT_INIT = 16'h0f7f;
    SB_LUT4 i1_2_lut_rep_16_3_lut_4_lut (.I0(n3857), .I1(VGA_X[8]), .I2(n3549), 
            .I3(n3856), .O(n3852));
    defparam i1_2_lut_rep_16_3_lut_4_lut.LUT_INIT = 16'hf080;
    SB_LUT4 i2242_3_lut_4_lut (.I0(n3857), .I1(VGA_X[8]), .I2(VGA_X[9]), 
            .I3(VGA_X[10]), .O(n3603));
    defparam i2242_3_lut_4_lut.LUT_INIT = 16'hf800;
    SB_LUT4 mux_15_i9_3_lut_4_lut (.I0(n3855), .I1(n3549), .I2(n190[8]), 
            .I3(\TX_ADDR[8] ), .O(n212));   // ../vga_control.v(57[28:124])
    defparam mux_15_i9_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 mux_15_i10_3_lut_4_lut (.I0(n3855), .I1(n3549), .I2(n190[9]), 
            .I3(\TX_ADDR[9] ), .O(n211));   // ../vga_control.v(57[28:124])
    defparam mux_15_i10_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i1777_4_lut (.I0(n3029), .I1(VGA_X[10]), .I2(VGA_X[9]), .I3(VGA_X[8]), 
            .O(n2030));
    defparam i1777_4_lut.LUT_INIT = 16'hc8c0;
    SB_LUT4 mux_15_i8_3_lut_4_lut (.I0(n3855), .I1(n3549), .I2(n190[7]), 
            .I3(\TX_ADDR[7] ), .O(n213));   // ../vga_control.v(57[28:124])
    defparam mux_15_i8_3_lut_4_lut.LUT_INIT = 16'hf780;
    SB_LUT4 i271_2_lut_3_lut_4_lut_rep_29 (.I0(ADV_HSYNC_c), .I1(old_VGA_HS), 
            .I2(ADV_VSYNC_c), .I3(n3549), .O(n3865));   // ../vga_control.v(57[28:124])
    defparam i271_2_lut_3_lut_4_lut_rep_29.LUT_INIT = 16'hf4f0;
    SB_LUT4 i271_2_lut_3_lut_4_lut_rep_28 (.I0(ADV_HSYNC_c), .I1(old_VGA_HS), 
            .I2(ADV_VSYNC_c), .I3(n3549), .O(n3864));   // ../vga_control.v(57[28:124])
    defparam i271_2_lut_3_lut_4_lut_rep_28.LUT_INIT = 16'hf4f0;
    SB_LUT4 mux_15_i5_3_lut_4_lut (.I0(n3855), .I1(n3549), .I2(n190[4]), 
            .I3(\TX_ADDR[4] ), .O(n216));   // ../vga_control.v(57[28:124])
    defparam mux_15_i5_3_lut_4_lut.LUT_INIT = 16'hf780;
    
endmodule
//
// Verilog Description of module TX_PLL
//

module TX_PLL (TVP_CLK_c, VCC_net, GND_net, ADV_CLK_c) /* synthesis syn_module_defined=1 */ ;
    input TVP_CLK_c;
    input VCC_net;
    input GND_net;
    output ADV_CLK_c;
    
    wire TVP_CLK_c /* synthesis SET_AS_NETWORK=TVP_CLK_c, is_clock=1 */ ;   // ../main.v(3[13:20])
    wire ADV_CLK_c /* synthesis SET_AS_NETWORK=ADV_CLK_c, is_clock=1 */ ;   // ../main.v(13[14:21])
    
    SB_PLL40_CORE TX_PLL_inst (.REFERENCECLK(TVP_CLK_c), .PLLOUTCORE(ADV_CLK_c), 
            .BYPASS(GND_net), .RESETB(VCC_net)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=14, LSE_LCOL=9, LSE_RCOL=27, LSE_LLINE=20, LSE_RLINE=24 */ ;   // ../main.v(20[9] 24[27])
    defparam TX_PLL_inst.FEEDBACK_PATH = "SIMPLE";
    defparam TX_PLL_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
    defparam TX_PLL_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
    defparam TX_PLL_inst.SHIFTREG_DIV_MODE = 2'b00;
    defparam TX_PLL_inst.FDA_FEEDBACK = 4'b0000;
    defparam TX_PLL_inst.FDA_RELATIVE = 4'b0000;
    defparam TX_PLL_inst.PLLOUT_SELECT = "GENCLK";
    defparam TX_PLL_inst.DIVR = 4'b0000;
    defparam TX_PLL_inst.DIVF = 7'b0100110;
    defparam TX_PLL_inst.DIVQ = 3'b100;
    defparam TX_PLL_inst.FILTER_RANGE = 3'b010;
    defparam TX_PLL_inst.ENABLE_ICEGATE = 1'b0;
    defparam TX_PLL_inst.TEST_MODE = 1'b0;
    defparam TX_PLL_inst.EXTERNAL_DIVIDE_FACTOR = 1;
    
endmodule
//
// Verilog Description of module RAM
//

module RAM (\TX_ADDR[11] , \TX_ADDR[12] , TX_DATA, ADV_CLK_c, DEBUG_c_2, 
            \RX_ADDR[0] , \RX_ADDR[1] , \RX_ADDR[2] , \RX_ADDR[3] , 
            \RX_ADDR[4] , \RX_ADDR[5] , \RX_ADDR[6] , \RX_ADDR[7] , 
            \RX_ADDR[8] , \RX_ADDR[9] , \RX_ADDR[10] , n28, n27, n26, 
            n25, n24, n23, n22, n21, n20, n19, n18, TVP_VIDEO_c_8, 
            TVP_VIDEO_c_9, TVP_CLK_c, VCC_net, TVP_VIDEO_c_6, TVP_VIDEO_c_7, 
            TVP_VIDEO_c_4, TVP_VIDEO_c_5, TVP_VIDEO_c_2, TVP_VIDEO_c_3, 
            \RX_ADDR[11] , \RX_ADDR[12] , DEBUG_c_3, DEBUG_c_5, GND_net) /* synthesis syn_module_defined=1 */ ;
    input \TX_ADDR[11] ;
    input \TX_ADDR[12] ;
    output [7:0]TX_DATA;
    input ADV_CLK_c;
    input DEBUG_c_2;
    input \RX_ADDR[0] ;
    input \RX_ADDR[1] ;
    input \RX_ADDR[2] ;
    input \RX_ADDR[3] ;
    input \RX_ADDR[4] ;
    input \RX_ADDR[5] ;
    input \RX_ADDR[6] ;
    input \RX_ADDR[7] ;
    input \RX_ADDR[8] ;
    input \RX_ADDR[9] ;
    input \RX_ADDR[10] ;
    input n28;
    input n27;
    input n26;
    input n25;
    input n24;
    input n23;
    input n22;
    input n21;
    input n20;
    input n19;
    input n18;
    input TVP_VIDEO_c_8;
    input TVP_VIDEO_c_9;
    input TVP_CLK_c;
    input VCC_net;
    input TVP_VIDEO_c_6;
    input TVP_VIDEO_c_7;
    input TVP_VIDEO_c_4;
    input TVP_VIDEO_c_5;
    input TVP_VIDEO_c_2;
    input TVP_VIDEO_c_3;
    input \RX_ADDR[11] ;
    input \RX_ADDR[12] ;
    input DEBUG_c_3;
    input DEBUG_c_5;
    input GND_net;
    
    wire ADV_CLK_c /* synthesis SET_AS_NETWORK=ADV_CLK_c, is_clock=1 */ ;   // ../main.v(13[14:21])
    wire TVP_CLK_c /* synthesis SET_AS_NETWORK=TVP_CLK_c, is_clock=1 */ ;   // ../main.v(3[13:20])
    
    wire n626, n634, n3779;
    wire [7:0]dout_7__N_553;
    
    wire n570, n562, n3782, n3705, n3706, n3773, n566, n567, 
        n577, n499, n500, n512, n497, n498, n495, n496, n564, 
        n565, n598, n599, n609, n563, n560, n561, n596, n597, 
        n509, n510, n513, n594, n595, n592, n593, n507, n508, 
        n630, n631, n641, n505, n506, n503, n504, n628, n629, 
        n574, n575, n578, n627, n624, n625, n572, n573, n606, 
        n607, n610, n571, n568, n569, n604, n605, n638, n639, 
        n642, n602, n603, n3833, n600, n601, n3836, n636, n637, 
        n501, n502, n635, n632, n633, n3827, n3830, n3821, n3824, 
        n3815, n3818, n3809, n3812, n3803, n3806, n3699, n3700, 
        n3797, n3721, n3720, n3702, n3703, n3791, n3718, n3717, 
        n3785, n3788, n3761, n3764, n3714, n3715, n3770, n3767;
    
    SB_LUT4 TX_ADDR_11__bdd_4_lut_2420 (.I0(\TX_ADDR[11] ), .I1(n626), .I2(n634), 
            .I3(\TX_ADDR[12] ), .O(n3779));
    defparam TX_ADDR_11__bdd_4_lut_2420.LUT_INIT = 16'he4aa;
    SB_DFF dout_i0 (.Q(TX_DATA[0]), .C(ADV_CLK_c), .D(dout_7__N_553[0]));   // ../ram.v(14[9] 16[5])
    SB_LUT4 n3779_bdd_4_lut (.I0(n3779), .I1(n570), .I2(n562), .I3(\TX_ADDR[12] ), 
            .O(n3782));
    defparam n3779_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 TX_ADDR_12__bdd_4_lut_2425 (.I0(\TX_ADDR[12] ), .I1(n3705), 
            .I2(n3706), .I3(DEBUG_c_2), .O(n3773));
    defparam TX_ADDR_12__bdd_4_lut_2425.LUT_INIT = 16'he4aa;
    SB_RAM2048x2 mem0 (.RDATA({n567, n566}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n577), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_9, TVP_VIDEO_c_8}));
    defparam mem0.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem0.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem8 (.RDATA({n500, n499}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n512), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_7, TVP_VIDEO_c_6}));
    defparam mem8.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem8.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem9 (.RDATA({n498, n497}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n512), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_5, TVP_VIDEO_c_4}));
    defparam mem9.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem9.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem10 (.RDATA({n496, n495}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n512), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_3, TVP_VIDEO_c_2}));
    defparam mem10.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem10.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem11 (.RDATA({n565, n564}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n577), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_7, TVP_VIDEO_c_6}));
    defparam mem11.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem11.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem1 (.RDATA({n599, n598}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n609), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_9, TVP_VIDEO_c_8}));
    defparam mem1.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem1.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem1.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem1.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem1.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem1.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem1.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem1.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem1.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem1.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem1.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem1.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem1.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem1.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem1.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem1.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_LUT4 i1_2_lut_3_lut_4_lut (.I0(\RX_ADDR[11] ), .I1(\RX_ADDR[12] ), 
            .I2(DEBUG_c_3), .I3(DEBUG_c_5), .O(n577));
    defparam i1_2_lut_3_lut_4_lut.LUT_INIT = 16'h1000;
    SB_RAM2048x2 mem12 (.RDATA({n563, n562}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n577), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_5, TVP_VIDEO_c_4}));
    defparam mem12.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem12.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem13 (.RDATA({n561, n560}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n577), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_3, TVP_VIDEO_c_2}));
    defparam mem13.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem13.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem14 (.RDATA({n597, n596}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n609), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_7, TVP_VIDEO_c_6}));
    defparam mem14.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem14.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem14.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem14.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem14.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem14.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem14.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem14.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem14.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem14.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem14.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem14.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem14.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem14.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem14.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem14.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem2 (.RDATA({n510, n509}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n513), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_9, TVP_VIDEO_c_8}));
    defparam mem2.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem2.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem15 (.RDATA({n595, n594}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n609), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_5, TVP_VIDEO_c_4}));
    defparam mem15.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem15.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem15.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem15.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem15.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem15.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem15.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem15.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem15.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem15.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem15.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem15.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem15.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem15.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem15.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem15.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem16 (.RDATA({n593, n592}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n609), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_3, TVP_VIDEO_c_2}));
    defparam mem16.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem16.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem16.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem16.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem16.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem16.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem16.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem16.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem16.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem16.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem16.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem16.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem16.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem16.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem16.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem16.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem17 (.RDATA({n508, n507}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n513), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_7, TVP_VIDEO_c_6}));
    defparam mem17.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem17.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem3 (.RDATA({n631, n630}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n641), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_9, TVP_VIDEO_c_8}));
    defparam mem3.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem3.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_LUT4 i2390_2_lut_3_lut_4_lut (.I0(\RX_ADDR[11] ), .I1(\RX_ADDR[12] ), 
            .I2(DEBUG_c_3), .I3(DEBUG_c_5), .O(n512));
    defparam i2390_2_lut_3_lut_4_lut.LUT_INIT = 16'h0100;
    SB_RAM2048x2 mem18 (.RDATA({n506, n505}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n513), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_5, TVP_VIDEO_c_4}));
    defparam mem18.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem18.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem19 (.RDATA({n504, n503}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n513), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_3, TVP_VIDEO_c_2}));
    defparam mem19.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem19.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem20 (.RDATA({n629, n628}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n641), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_7, TVP_VIDEO_c_6}));
    defparam mem20.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem20.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem4 (.RDATA({n575, n574}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n578), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_9, TVP_VIDEO_c_8}));
    defparam mem4.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem4.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem21 (.RDATA({n627, n626}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n641), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_5, TVP_VIDEO_c_4}));
    defparam mem21.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem21.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem22 (.RDATA({n625, n624}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n641), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_3, TVP_VIDEO_c_2}));
    defparam mem22.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem22.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem23 (.RDATA({n573, n572}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n578), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_7, TVP_VIDEO_c_6}));
    defparam mem23.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem23.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem5 (.RDATA({n607, n606}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n610), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_9, TVP_VIDEO_c_8}));
    defparam mem5.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem5.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem5.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem5.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem5.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem5.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem5.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem5.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem5.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem5.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem5.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem5.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem5.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem5.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem5.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem5.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem24 (.RDATA({n571, n570}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n578), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_5, TVP_VIDEO_c_4}));
    defparam mem24.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem24.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem25 (.RDATA({n569, n568}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n578), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_3, TVP_VIDEO_c_2}));
    defparam mem25.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem25.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem26 (.RDATA({n605, n604}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n610), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_7, TVP_VIDEO_c_6}));
    defparam mem26.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem26.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem26.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem26.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem26.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem26.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem26.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem26.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem26.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem26.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem26.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem26.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem26.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem26.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem26.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem26.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem6 (.RDATA({n639, n638}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n642), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_9, TVP_VIDEO_c_8}));
    defparam mem6.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem6.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem6.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem6.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem6.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem6.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem6.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem6.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem6.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem6.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem6.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem6.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem6.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem6.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem6.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem6.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem27 (.RDATA({n603, n602}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n610), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_5, TVP_VIDEO_c_4}));
    defparam mem27.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem27.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem27.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem27.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem27.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem27.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem27.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem27.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem27.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem27.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem27.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem27.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem27.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem27.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem27.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem27.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_LUT4 TX_ADDR_11__bdd_4_lut (.I0(\TX_ADDR[11] ), .I1(n597), .I2(n605), 
            .I3(\TX_ADDR[12] ), .O(n3833));
    defparam TX_ADDR_11__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_RAM2048x2 mem28 (.RDATA({n601, n600}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n610), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_3, TVP_VIDEO_c_2}));
    defparam mem28.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem28.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem28.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem28.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem28.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem28.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem28.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem28.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem28.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem28.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem28.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem28.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem28.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem28.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem28.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem28.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_LUT4 n3833_bdd_4_lut (.I0(n3833), .I1(n508), .I2(n500), .I3(\TX_ADDR[12] ), 
            .O(n3836));
    defparam n3833_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_RAM2048x2 mem29 (.RDATA({n637, n636}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n642), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_7, TVP_VIDEO_c_6}));
    defparam mem29.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem29.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem29.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem29.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem29.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem29.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem29.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem29.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem29.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem29.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem29.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem29.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem29.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem29.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem29.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem29.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem7 (.RDATA({n502, n501}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n512), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_9, TVP_VIDEO_c_8}));
    defparam mem7.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem7.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem30 (.RDATA({n635, n634}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n642), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_5, TVP_VIDEO_c_4}));
    defparam mem30.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem30.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem30.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem30.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem30.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem30.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem30.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem30.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem30.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem30.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem30.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem30.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem30.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem30.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem30.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem30.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM2048x2 mem31 (.RDATA({n633, n632}), .RCLK(ADV_CLK_c), .RCLKE(VCC_net), 
            .RE(VCC_net), .RADDR({n18, n19, n20, n21, n22, n23, 
            n24, n25, n26, n27, n28}), .WCLK(TVP_CLK_c), .WCLKE(VCC_net), 
            .WE(n642), .WADDR({\RX_ADDR[10] , \RX_ADDR[9] , \RX_ADDR[8] , 
            \RX_ADDR[7] , \RX_ADDR[6] , \RX_ADDR[5] , \RX_ADDR[4] , 
            \RX_ADDR[3] , \RX_ADDR[2] , \RX_ADDR[1] , \RX_ADDR[0] }), 
            .WDATA({TVP_VIDEO_c_3, TVP_VIDEO_c_2}));
    defparam mem31.INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem31.INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem31.INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem31.INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem31.INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem31.INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem31.INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem31.INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem31.INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem31.INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem31.INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem31.INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem31.INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem31.INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem31.INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam mem31.INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    SB_LUT4 TX_ADDR_11__bdd_4_lut_2460 (.I0(\TX_ADDR[11] ), .I1(n625), .I2(n633), 
            .I3(\TX_ADDR[12] ), .O(n3827));
    defparam TX_ADDR_11__bdd_4_lut_2460.LUT_INIT = 16'he4aa;
    SB_LUT4 n3827_bdd_4_lut (.I0(n3827), .I1(n569), .I2(n561), .I3(\TX_ADDR[12] ), 
            .O(n3830));
    defparam n3827_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 TX_ADDR_11__bdd_4_lut_2455 (.I0(\TX_ADDR[11] ), .I1(n624), .I2(n632), 
            .I3(\TX_ADDR[12] ), .O(n3821));
    defparam TX_ADDR_11__bdd_4_lut_2455.LUT_INIT = 16'he4aa;
    SB_DFF dout_i1 (.Q(TX_DATA[1]), .C(ADV_CLK_c), .D(dout_7__N_553[1]));   // ../ram.v(14[9] 16[5])
    SB_LUT4 n3821_bdd_4_lut (.I0(n3821), .I1(n568), .I2(n560), .I3(\TX_ADDR[12] ), 
            .O(n3824));
    defparam n3821_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 TX_ADDR_11__bdd_4_lut_2450 (.I0(\TX_ADDR[11] ), .I1(n592), .I2(n600), 
            .I3(\TX_ADDR[12] ), .O(n3815));
    defparam TX_ADDR_11__bdd_4_lut_2450.LUT_INIT = 16'he4aa;
    SB_LUT4 n3815_bdd_4_lut (.I0(n3815), .I1(n503), .I2(n495), .I3(\TX_ADDR[12] ), 
            .O(n3818));
    defparam n3815_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 TX_ADDR_11__bdd_4_lut_2445 (.I0(\TX_ADDR[11] ), .I1(n593), .I2(n601), 
            .I3(\TX_ADDR[12] ), .O(n3809));
    defparam TX_ADDR_11__bdd_4_lut_2445.LUT_INIT = 16'he4aa;
    SB_LUT4 n3809_bdd_4_lut (.I0(n3809), .I1(n504), .I2(n496), .I3(\TX_ADDR[12] ), 
            .O(n3812));
    defparam n3809_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 TX_ADDR_11__bdd_4_lut_2440 (.I0(\TX_ADDR[11] ), .I1(n594), .I2(n602), 
            .I3(\TX_ADDR[12] ), .O(n3803));
    defparam TX_ADDR_11__bdd_4_lut_2440.LUT_INIT = 16'he4aa;
    SB_LUT4 n3803_bdd_4_lut (.I0(n3803), .I1(n505), .I2(n497), .I3(\TX_ADDR[12] ), 
            .O(n3806));
    defparam n3803_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 TX_ADDR_12__bdd_4_lut (.I0(\TX_ADDR[12] ), .I1(n3699), .I2(n3700), 
            .I3(DEBUG_c_2), .O(n3797));
    defparam TX_ADDR_12__bdd_4_lut.LUT_INIT = 16'he4aa;
    SB_LUT4 n3797_bdd_4_lut (.I0(n3797), .I1(n3721), .I2(n3720), .I3(DEBUG_c_2), 
            .O(dout_7__N_553[4]));
    defparam n3797_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 TX_ADDR_12__bdd_4_lut_2430 (.I0(\TX_ADDR[12] ), .I1(n3702), 
            .I2(n3703), .I3(DEBUG_c_2), .O(n3791));
    defparam TX_ADDR_12__bdd_4_lut_2430.LUT_INIT = 16'he4aa;
    SB_LUT4 n3791_bdd_4_lut (.I0(n3791), .I1(n3718), .I2(n3717), .I3(DEBUG_c_2), 
            .O(dout_7__N_553[7]));
    defparam n3791_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 TX_ADDR_11__bdd_4_lut_2435 (.I0(\TX_ADDR[11] ), .I1(n630), .I2(n638), 
            .I3(\TX_ADDR[12] ), .O(n3785));
    defparam TX_ADDR_11__bdd_4_lut_2435.LUT_INIT = 16'he4aa;
    SB_LUT4 n3785_bdd_4_lut (.I0(n3785), .I1(n574), .I2(n566), .I3(\TX_ADDR[12] ), 
            .O(n3788));
    defparam n3785_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_7 (.I0(\RX_ADDR[12] ), .I1(\RX_ADDR[11] ), 
            .I2(DEBUG_c_3), .I3(DEBUG_c_5), .O(n641));
    defparam i1_2_lut_3_lut_4_lut_adj_7.LUT_INIT = 16'h2000;
    SB_LUT4 n3761_bdd_4_lut (.I0(n3761), .I1(n573), .I2(n565), .I3(\TX_ADDR[12] ), 
            .O(n3764));
    defparam n3761_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_8 (.I0(\RX_ADDR[12] ), .I1(\RX_ADDR[11] ), 
            .I2(DEBUG_c_3), .I3(DEBUG_c_5), .O(n609));
    defparam i1_2_lut_3_lut_4_lut_adj_8.LUT_INIT = 16'h0200;
    SB_LUT4 i2352_3_lut (.I0(n498), .I1(n506), .I2(\TX_ADDR[11] ), .I3(GND_net), 
            .O(n3714));
    defparam i2352_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2353_3_lut (.I0(n595), .I1(n603), .I2(\TX_ADDR[11] ), .I3(GND_net), 
            .O(n3715));
    defparam i2353_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i182929_i1_3_lut (.I0(n3770), .I1(n3788), .I2(DEBUG_c_2), 
            .I3(GND_net), .O(dout_7__N_553[6]));
    defparam i182929_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i182326_i1_3_lut (.I0(n3836), .I1(n3764), .I2(DEBUG_c_2), 
            .I3(GND_net), .O(dout_7__N_553[5]));
    defparam i182326_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_DFF dout_i2 (.Q(TX_DATA[2]), .C(ADV_CLK_c), .D(dout_7__N_553[2]));   // ../ram.v(14[9] 16[5])
    SB_DFF dout_i3 (.Q(TX_DATA[3]), .C(ADV_CLK_c), .D(dout_7__N_553[3]));   // ../ram.v(14[9] 16[5])
    SB_DFF dout_i4 (.Q(TX_DATA[4]), .C(ADV_CLK_c), .D(dout_7__N_553[4]));   // ../ram.v(14[9] 16[5])
    SB_DFF dout_i5 (.Q(TX_DATA[5]), .C(ADV_CLK_c), .D(dout_7__N_553[5]));   // ../ram.v(14[9] 16[5])
    SB_DFF dout_i6 (.Q(TX_DATA[6]), .C(ADV_CLK_c), .D(dout_7__N_553[6]));   // ../ram.v(14[9] 16[5])
    SB_DFF dout_i7 (.Q(TX_DATA[7]), .C(ADV_CLK_c), .D(dout_7__N_553[7]));   // ../ram.v(14[9] 16[5])
    SB_LUT4 i180517_i1_3_lut (.I0(n3806), .I1(n3782), .I2(DEBUG_c_2), 
            .I3(GND_net), .O(dout_7__N_553[2]));
    defparam i180517_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 n3773_bdd_4_lut (.I0(n3773), .I1(n3715), .I2(n3714), .I3(DEBUG_c_2), 
            .O(dout_7__N_553[3]));
    defparam n3773_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 i2355_3_lut (.I0(n502), .I1(n510), .I2(\TX_ADDR[11] ), .I3(GND_net), 
            .O(n3717));
    defparam i2355_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2356_3_lut (.I0(n599), .I1(n607), .I2(\TX_ADDR[11] ), .I3(GND_net), 
            .O(n3718));
    defparam i2356_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2341_3_lut (.I0(n631), .I1(n639), .I2(\TX_ADDR[11] ), .I3(GND_net), 
            .O(n3703));
    defparam i2341_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2340_3_lut (.I0(n567), .I1(n575), .I2(\TX_ADDR[11] ), .I3(GND_net), 
            .O(n3702));
    defparam i2340_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2358_3_lut (.I0(n499), .I1(n507), .I2(\TX_ADDR[11] ), .I3(GND_net), 
            .O(n3720));
    defparam i2358_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2359_3_lut (.I0(n596), .I1(n604), .I2(\TX_ADDR[11] ), .I3(GND_net), 
            .O(n3721));
    defparam i2359_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2338_3_lut (.I0(n628), .I1(n636), .I2(\TX_ADDR[11] ), .I3(GND_net), 
            .O(n3700));
    defparam i2338_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2337_3_lut (.I0(n564), .I1(n572), .I2(\TX_ADDR[11] ), .I3(GND_net), 
            .O(n3699));
    defparam i2337_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i179914_i1_3_lut (.I0(n3812), .I1(n3830), .I2(DEBUG_c_2), 
            .I3(GND_net), .O(dout_7__N_553[1]));
    defparam i179914_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_9 (.I0(\RX_ADDR[11] ), .I1(\RX_ADDR[12] ), 
            .I2(DEBUG_c_3), .I3(DEBUG_c_5), .O(n578));
    defparam i1_2_lut_3_lut_4_lut_adj_9.LUT_INIT = 16'h2000;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_10 (.I0(\RX_ADDR[11] ), .I1(\RX_ADDR[12] ), 
            .I2(DEBUG_c_3), .I3(DEBUG_c_5), .O(n513));
    defparam i1_2_lut_3_lut_4_lut_adj_10.LUT_INIT = 16'h0200;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_11 (.I0(\RX_ADDR[12] ), .I1(\RX_ADDR[11] ), 
            .I2(DEBUG_c_3), .I3(DEBUG_c_5), .O(n642));
    defparam i1_2_lut_3_lut_4_lut_adj_11.LUT_INIT = 16'h8000;
    SB_LUT4 i1_2_lut_3_lut_4_lut_adj_12 (.I0(\RX_ADDR[12] ), .I1(\RX_ADDR[11] ), 
            .I2(DEBUG_c_3), .I3(DEBUG_c_5), .O(n610));
    defparam i1_2_lut_3_lut_4_lut_adj_12.LUT_INIT = 16'h0800;
    SB_LUT4 i179311_i1_3_lut (.I0(n3818), .I1(n3824), .I2(DEBUG_c_2), 
            .I3(GND_net), .O(dout_7__N_553[0]));
    defparam i179311_i1_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2344_3_lut (.I0(n627), .I1(n635), .I2(\TX_ADDR[11] ), .I3(GND_net), 
            .O(n3706));
    defparam i2344_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 i2343_3_lut (.I0(n563), .I1(n571), .I2(\TX_ADDR[11] ), .I3(GND_net), 
            .O(n3705));
    defparam i2343_3_lut.LUT_INIT = 16'hcaca;
    SB_LUT4 TX_ADDR_11__bdd_4_lut_2415 (.I0(\TX_ADDR[11] ), .I1(n598), .I2(n606), 
            .I3(\TX_ADDR[12] ), .O(n3767));
    defparam TX_ADDR_11__bdd_4_lut_2415.LUT_INIT = 16'he4aa;
    SB_LUT4 n3767_bdd_4_lut (.I0(n3767), .I1(n509), .I2(n501), .I3(\TX_ADDR[12] ), 
            .O(n3770));
    defparam n3767_bdd_4_lut.LUT_INIT = 16'haad8;
    SB_LUT4 TX_ADDR_11__bdd_4_lut_2406 (.I0(\TX_ADDR[11] ), .I1(n629), .I2(n637), 
            .I3(\TX_ADDR[12] ), .O(n3761));
    defparam TX_ADDR_11__bdd_4_lut_2406.LUT_INIT = 16'he4aa;
    
endmodule
