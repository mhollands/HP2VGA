-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     Sep 23 2018 23:07:33

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "main" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of main
entity main is
port (
    TVP_VIDEO : in std_logic_vector(9 downto 0);
    ADV_B : out std_logic_vector(7 downto 0);
    ADV_G : out std_logic_vector(7 downto 0);
    ADV_R : out std_logic_vector(7 downto 0);
    DEBUG : inout std_logic_vector(7 downto 0);
    TVP_CLK : in std_logic;
    ADV_CLK : out std_logic;
    TVP_HSYNC : in std_logic;
    ADV_HSYNC : out std_logic;
    TVP_VSYNC : in std_logic;
    ADV_VSYNC : out std_logic;
    ADV_BLANK_N : out std_logic;
    LED : out std_logic;
    ADV_SYNC_N : out std_logic);
end main;

-- Architecture of main
-- View name is \INTERFACE\
architecture \INTERFACE\ of main is

signal \N__24376\ : std_logic;
signal \N__24375\ : std_logic;
signal \N__24374\ : std_logic;
signal \N__24365\ : std_logic;
signal \N__24364\ : std_logic;
signal \N__24363\ : std_logic;
signal \N__24356\ : std_logic;
signal \N__24355\ : std_logic;
signal \N__24354\ : std_logic;
signal \N__24347\ : std_logic;
signal \N__24346\ : std_logic;
signal \N__24345\ : std_logic;
signal \N__24338\ : std_logic;
signal \N__24337\ : std_logic;
signal \N__24336\ : std_logic;
signal \N__24329\ : std_logic;
signal \N__24328\ : std_logic;
signal \N__24327\ : std_logic;
signal \N__24320\ : std_logic;
signal \N__24319\ : std_logic;
signal \N__24318\ : std_logic;
signal \N__24311\ : std_logic;
signal \N__24310\ : std_logic;
signal \N__24309\ : std_logic;
signal \N__24302\ : std_logic;
signal \N__24301\ : std_logic;
signal \N__24300\ : std_logic;
signal \N__24293\ : std_logic;
signal \N__24292\ : std_logic;
signal \N__24291\ : std_logic;
signal \N__24284\ : std_logic;
signal \N__24283\ : std_logic;
signal \N__24282\ : std_logic;
signal \N__24275\ : std_logic;
signal \N__24274\ : std_logic;
signal \N__24273\ : std_logic;
signal \N__24266\ : std_logic;
signal \N__24265\ : std_logic;
signal \N__24264\ : std_logic;
signal \N__24257\ : std_logic;
signal \N__24256\ : std_logic;
signal \N__24255\ : std_logic;
signal \N__24248\ : std_logic;
signal \N__24247\ : std_logic;
signal \N__24246\ : std_logic;
signal \N__24239\ : std_logic;
signal \N__24238\ : std_logic;
signal \N__24237\ : std_logic;
signal \N__24230\ : std_logic;
signal \N__24229\ : std_logic;
signal \N__24228\ : std_logic;
signal \N__24221\ : std_logic;
signal \N__24220\ : std_logic;
signal \N__24219\ : std_logic;
signal \N__24212\ : std_logic;
signal \N__24211\ : std_logic;
signal \N__24210\ : std_logic;
signal \N__24203\ : std_logic;
signal \N__24202\ : std_logic;
signal \N__24201\ : std_logic;
signal \N__24194\ : std_logic;
signal \N__24193\ : std_logic;
signal \N__24192\ : std_logic;
signal \N__24185\ : std_logic;
signal \N__24184\ : std_logic;
signal \N__24183\ : std_logic;
signal \N__24176\ : std_logic;
signal \N__24175\ : std_logic;
signal \N__24174\ : std_logic;
signal \N__24167\ : std_logic;
signal \N__24166\ : std_logic;
signal \N__24165\ : std_logic;
signal \N__24158\ : std_logic;
signal \N__24157\ : std_logic;
signal \N__24156\ : std_logic;
signal \N__24149\ : std_logic;
signal \N__24148\ : std_logic;
signal \N__24147\ : std_logic;
signal \N__24140\ : std_logic;
signal \N__24139\ : std_logic;
signal \N__24138\ : std_logic;
signal \N__24131\ : std_logic;
signal \N__24130\ : std_logic;
signal \N__24129\ : std_logic;
signal \N__24122\ : std_logic;
signal \N__24121\ : std_logic;
signal \N__24120\ : std_logic;
signal \N__24113\ : std_logic;
signal \N__24112\ : std_logic;
signal \N__24111\ : std_logic;
signal \N__24104\ : std_logic;
signal \N__24103\ : std_logic;
signal \N__24102\ : std_logic;
signal \N__24095\ : std_logic;
signal \N__24094\ : std_logic;
signal \N__24093\ : std_logic;
signal \N__24086\ : std_logic;
signal \N__24085\ : std_logic;
signal \N__24084\ : std_logic;
signal \N__24077\ : std_logic;
signal \N__24076\ : std_logic;
signal \N__24075\ : std_logic;
signal \N__24068\ : std_logic;
signal \N__24067\ : std_logic;
signal \N__24066\ : std_logic;
signal \N__24059\ : std_logic;
signal \N__24058\ : std_logic;
signal \N__24057\ : std_logic;
signal \N__24050\ : std_logic;
signal \N__24049\ : std_logic;
signal \N__24048\ : std_logic;
signal \N__24041\ : std_logic;
signal \N__24040\ : std_logic;
signal \N__24039\ : std_logic;
signal \N__24032\ : std_logic;
signal \N__24031\ : std_logic;
signal \N__24030\ : std_logic;
signal \N__24023\ : std_logic;
signal \N__24022\ : std_logic;
signal \N__24021\ : std_logic;
signal \N__24014\ : std_logic;
signal \N__24013\ : std_logic;
signal \N__24012\ : std_logic;
signal \N__24005\ : std_logic;
signal \N__24004\ : std_logic;
signal \N__24003\ : std_logic;
signal \N__23996\ : std_logic;
signal \N__23995\ : std_logic;
signal \N__23994\ : std_logic;
signal \N__23987\ : std_logic;
signal \N__23986\ : std_logic;
signal \N__23985\ : std_logic;
signal \N__23978\ : std_logic;
signal \N__23977\ : std_logic;
signal \N__23976\ : std_logic;
signal \N__23969\ : std_logic;
signal \N__23968\ : std_logic;
signal \N__23967\ : std_logic;
signal \N__23960\ : std_logic;
signal \N__23959\ : std_logic;
signal \N__23958\ : std_logic;
signal \N__23951\ : std_logic;
signal \N__23950\ : std_logic;
signal \N__23949\ : std_logic;
signal \N__23942\ : std_logic;
signal \N__23941\ : std_logic;
signal \N__23940\ : std_logic;
signal \N__23923\ : std_logic;
signal \N__23920\ : std_logic;
signal \N__23917\ : std_logic;
signal \N__23914\ : std_logic;
signal \N__23911\ : std_logic;
signal \N__23908\ : std_logic;
signal \N__23905\ : std_logic;
signal \N__23902\ : std_logic;
signal \N__23899\ : std_logic;
signal \N__23896\ : std_logic;
signal \N__23893\ : std_logic;
signal \N__23890\ : std_logic;
signal \N__23887\ : std_logic;
signal \N__23884\ : std_logic;
signal \N__23881\ : std_logic;
signal \N__23878\ : std_logic;
signal \N__23875\ : std_logic;
signal \N__23872\ : std_logic;
signal \N__23869\ : std_logic;
signal \N__23866\ : std_logic;
signal \N__23863\ : std_logic;
signal \N__23860\ : std_logic;
signal \N__23859\ : std_logic;
signal \N__23856\ : std_logic;
signal \N__23855\ : std_logic;
signal \N__23852\ : std_logic;
signal \N__23851\ : std_logic;
signal \N__23850\ : std_logic;
signal \N__23849\ : std_logic;
signal \N__23848\ : std_logic;
signal \N__23847\ : std_logic;
signal \N__23846\ : std_logic;
signal \N__23845\ : std_logic;
signal \N__23844\ : std_logic;
signal \N__23843\ : std_logic;
signal \N__23842\ : std_logic;
signal \N__23841\ : std_logic;
signal \N__23840\ : std_logic;
signal \N__23839\ : std_logic;
signal \N__23838\ : std_logic;
signal \N__23837\ : std_logic;
signal \N__23836\ : std_logic;
signal \N__23833\ : std_logic;
signal \N__23830\ : std_logic;
signal \N__23829\ : std_logic;
signal \N__23828\ : std_logic;
signal \N__23825\ : std_logic;
signal \N__23822\ : std_logic;
signal \N__23819\ : std_logic;
signal \N__23818\ : std_logic;
signal \N__23813\ : std_logic;
signal \N__23808\ : std_logic;
signal \N__23807\ : std_logic;
signal \N__23806\ : std_logic;
signal \N__23803\ : std_logic;
signal \N__23800\ : std_logic;
signal \N__23795\ : std_logic;
signal \N__23790\ : std_logic;
signal \N__23783\ : std_logic;
signal \N__23780\ : std_logic;
signal \N__23775\ : std_logic;
signal \N__23772\ : std_logic;
signal \N__23769\ : std_logic;
signal \N__23762\ : std_logic;
signal \N__23759\ : std_logic;
signal \N__23756\ : std_logic;
signal \N__23753\ : std_logic;
signal \N__23750\ : std_logic;
signal \N__23747\ : std_logic;
signal \N__23742\ : std_logic;
signal \N__23741\ : std_logic;
signal \N__23736\ : std_logic;
signal \N__23731\ : std_logic;
signal \N__23720\ : std_logic;
signal \N__23715\ : std_logic;
signal \N__23712\ : std_logic;
signal \N__23709\ : std_logic;
signal \N__23706\ : std_logic;
signal \N__23703\ : std_logic;
signal \N__23700\ : std_logic;
signal \N__23697\ : std_logic;
signal \N__23694\ : std_logic;
signal \N__23685\ : std_logic;
signal \N__23674\ : std_logic;
signal \N__23671\ : std_logic;
signal \N__23668\ : std_logic;
signal \N__23665\ : std_logic;
signal \N__23662\ : std_logic;
signal \N__23659\ : std_logic;
signal \N__23656\ : std_logic;
signal \N__23653\ : std_logic;
signal \N__23650\ : std_logic;
signal \N__23647\ : std_logic;
signal \N__23644\ : std_logic;
signal \N__23641\ : std_logic;
signal \N__23638\ : std_logic;
signal \N__23635\ : std_logic;
signal \N__23632\ : std_logic;
signal \N__23629\ : std_logic;
signal \N__23626\ : std_logic;
signal \N__23623\ : std_logic;
signal \N__23620\ : std_logic;
signal \N__23617\ : std_logic;
signal \N__23614\ : std_logic;
signal \N__23613\ : std_logic;
signal \N__23612\ : std_logic;
signal \N__23611\ : std_logic;
signal \N__23608\ : std_logic;
signal \N__23605\ : std_logic;
signal \N__23604\ : std_logic;
signal \N__23603\ : std_logic;
signal \N__23602\ : std_logic;
signal \N__23601\ : std_logic;
signal \N__23600\ : std_logic;
signal \N__23599\ : std_logic;
signal \N__23598\ : std_logic;
signal \N__23595\ : std_logic;
signal \N__23592\ : std_logic;
signal \N__23591\ : std_logic;
signal \N__23590\ : std_logic;
signal \N__23587\ : std_logic;
signal \N__23586\ : std_logic;
signal \N__23583\ : std_logic;
signal \N__23578\ : std_logic;
signal \N__23577\ : std_logic;
signal \N__23576\ : std_logic;
signal \N__23573\ : std_logic;
signal \N__23570\ : std_logic;
signal \N__23563\ : std_logic;
signal \N__23560\ : std_logic;
signal \N__23557\ : std_logic;
signal \N__23554\ : std_logic;
signal \N__23553\ : std_logic;
signal \N__23550\ : std_logic;
signal \N__23547\ : std_logic;
signal \N__23544\ : std_logic;
signal \N__23543\ : std_logic;
signal \N__23540\ : std_logic;
signal \N__23537\ : std_logic;
signal \N__23536\ : std_logic;
signal \N__23535\ : std_logic;
signal \N__23532\ : std_logic;
signal \N__23529\ : std_logic;
signal \N__23522\ : std_logic;
signal \N__23519\ : std_logic;
signal \N__23518\ : std_logic;
signal \N__23513\ : std_logic;
signal \N__23510\ : std_logic;
signal \N__23503\ : std_logic;
signal \N__23500\ : std_logic;
signal \N__23497\ : std_logic;
signal \N__23494\ : std_logic;
signal \N__23493\ : std_logic;
signal \N__23492\ : std_logic;
signal \N__23489\ : std_logic;
signal \N__23486\ : std_logic;
signal \N__23485\ : std_logic;
signal \N__23482\ : std_logic;
signal \N__23479\ : std_logic;
signal \N__23474\ : std_logic;
signal \N__23471\ : std_logic;
signal \N__23468\ : std_logic;
signal \N__23465\ : std_logic;
signal \N__23462\ : std_logic;
signal \N__23459\ : std_logic;
signal \N__23454\ : std_logic;
signal \N__23449\ : std_logic;
signal \N__23444\ : std_logic;
signal \N__23441\ : std_logic;
signal \N__23438\ : std_logic;
signal \N__23431\ : std_logic;
signal \N__23422\ : std_logic;
signal \N__23419\ : std_logic;
signal \N__23414\ : std_logic;
signal \N__23401\ : std_logic;
signal \N__23398\ : std_logic;
signal \N__23395\ : std_logic;
signal \N__23394\ : std_logic;
signal \N__23391\ : std_logic;
signal \N__23388\ : std_logic;
signal \N__23387\ : std_logic;
signal \N__23386\ : std_logic;
signal \N__23385\ : std_logic;
signal \N__23380\ : std_logic;
signal \N__23377\ : std_logic;
signal \N__23374\ : std_logic;
signal \N__23373\ : std_logic;
signal \N__23372\ : std_logic;
signal \N__23371\ : std_logic;
signal \N__23370\ : std_logic;
signal \N__23367\ : std_logic;
signal \N__23360\ : std_logic;
signal \N__23357\ : std_logic;
signal \N__23354\ : std_logic;
signal \N__23353\ : std_logic;
signal \N__23352\ : std_logic;
signal \N__23349\ : std_logic;
signal \N__23346\ : std_logic;
signal \N__23345\ : std_logic;
signal \N__23344\ : std_logic;
signal \N__23343\ : std_logic;
signal \N__23340\ : std_logic;
signal \N__23333\ : std_logic;
signal \N__23330\ : std_logic;
signal \N__23327\ : std_logic;
signal \N__23326\ : std_logic;
signal \N__23325\ : std_logic;
signal \N__23324\ : std_logic;
signal \N__23323\ : std_logic;
signal \N__23318\ : std_logic;
signal \N__23315\ : std_logic;
signal \N__23312\ : std_logic;
signal \N__23311\ : std_logic;
signal \N__23310\ : std_logic;
signal \N__23309\ : std_logic;
signal \N__23308\ : std_logic;
signal \N__23307\ : std_logic;
signal \N__23306\ : std_logic;
signal \N__23305\ : std_logic;
signal \N__23304\ : std_logic;
signal \N__23303\ : std_logic;
signal \N__23300\ : std_logic;
signal \N__23299\ : std_logic;
signal \N__23296\ : std_logic;
signal \N__23289\ : std_logic;
signal \N__23286\ : std_logic;
signal \N__23283\ : std_logic;
signal \N__23282\ : std_logic;
signal \N__23281\ : std_logic;
signal \N__23278\ : std_logic;
signal \N__23275\ : std_logic;
signal \N__23268\ : std_logic;
signal \N__23265\ : std_logic;
signal \N__23262\ : std_logic;
signal \N__23261\ : std_logic;
signal \N__23260\ : std_logic;
signal \N__23257\ : std_logic;
signal \N__23256\ : std_logic;
signal \N__23253\ : std_logic;
signal \N__23252\ : std_logic;
signal \N__23249\ : std_logic;
signal \N__23246\ : std_logic;
signal \N__23245\ : std_logic;
signal \N__23242\ : std_logic;
signal \N__23239\ : std_logic;
signal \N__23238\ : std_logic;
signal \N__23235\ : std_logic;
signal \N__23232\ : std_logic;
signal \N__23229\ : std_logic;
signal \N__23228\ : std_logic;
signal \N__23227\ : std_logic;
signal \N__23224\ : std_logic;
signal \N__23217\ : std_logic;
signal \N__23214\ : std_logic;
signal \N__23211\ : std_logic;
signal \N__23206\ : std_logic;
signal \N__23199\ : std_logic;
signal \N__23196\ : std_logic;
signal \N__23193\ : std_logic;
signal \N__23192\ : std_logic;
signal \N__23191\ : std_logic;
signal \N__23190\ : std_logic;
signal \N__23189\ : std_logic;
signal \N__23178\ : std_logic;
signal \N__23175\ : std_logic;
signal \N__23164\ : std_logic;
signal \N__23161\ : std_logic;
signal \N__23158\ : std_logic;
signal \N__23155\ : std_logic;
signal \N__23152\ : std_logic;
signal \N__23143\ : std_logic;
signal \N__23140\ : std_logic;
signal \N__23139\ : std_logic;
signal \N__23138\ : std_logic;
signal \N__23131\ : std_logic;
signal \N__23128\ : std_logic;
signal \N__23125\ : std_logic;
signal \N__23124\ : std_logic;
signal \N__23121\ : std_logic;
signal \N__23118\ : std_logic;
signal \N__23117\ : std_logic;
signal \N__23112\ : std_logic;
signal \N__23109\ : std_logic;
signal \N__23098\ : std_logic;
signal \N__23095\ : std_logic;
signal \N__23092\ : std_logic;
signal \N__23089\ : std_logic;
signal \N__23082\ : std_logic;
signal \N__23079\ : std_logic;
signal \N__23074\ : std_logic;
signal \N__23071\ : std_logic;
signal \N__23068\ : std_logic;
signal \N__23065\ : std_logic;
signal \N__23062\ : std_logic;
signal \N__23055\ : std_logic;
signal \N__23046\ : std_logic;
signal \N__23043\ : std_logic;
signal \N__23040\ : std_logic;
signal \N__23037\ : std_logic;
signal \N__23032\ : std_logic;
signal \N__23029\ : std_logic;
signal \N__23026\ : std_logic;
signal \N__23023\ : std_logic;
signal \N__23020\ : std_logic;
signal \N__23011\ : std_logic;
signal \N__23008\ : std_logic;
signal \N__23005\ : std_logic;
signal \N__23002\ : std_logic;
signal \N__22999\ : std_logic;
signal \N__22996\ : std_logic;
signal \N__22993\ : std_logic;
signal \N__22990\ : std_logic;
signal \N__22987\ : std_logic;
signal \N__22984\ : std_logic;
signal \N__22981\ : std_logic;
signal \N__22978\ : std_logic;
signal \N__22975\ : std_logic;
signal \N__22972\ : std_logic;
signal \N__22969\ : std_logic;
signal \N__22966\ : std_logic;
signal \N__22963\ : std_logic;
signal \N__22960\ : std_logic;
signal \N__22957\ : std_logic;
signal \N__22954\ : std_logic;
signal \N__22951\ : std_logic;
signal \N__22948\ : std_logic;
signal \N__22945\ : std_logic;
signal \N__22942\ : std_logic;
signal \N__22939\ : std_logic;
signal \N__22936\ : std_logic;
signal \N__22933\ : std_logic;
signal \N__22930\ : std_logic;
signal \N__22927\ : std_logic;
signal \N__22924\ : std_logic;
signal \N__22921\ : std_logic;
signal \N__22918\ : std_logic;
signal \N__22915\ : std_logic;
signal \N__22912\ : std_logic;
signal \N__22909\ : std_logic;
signal \N__22906\ : std_logic;
signal \N__22903\ : std_logic;
signal \N__22900\ : std_logic;
signal \N__22897\ : std_logic;
signal \N__22894\ : std_logic;
signal \N__22891\ : std_logic;
signal \N__22888\ : std_logic;
signal \N__22885\ : std_logic;
signal \N__22882\ : std_logic;
signal \N__22879\ : std_logic;
signal \N__22876\ : std_logic;
signal \N__22873\ : std_logic;
signal \N__22870\ : std_logic;
signal \N__22869\ : std_logic;
signal \N__22866\ : std_logic;
signal \N__22865\ : std_logic;
signal \N__22862\ : std_logic;
signal \N__22859\ : std_logic;
signal \N__22858\ : std_logic;
signal \N__22857\ : std_logic;
signal \N__22856\ : std_logic;
signal \N__22853\ : std_logic;
signal \N__22850\ : std_logic;
signal \N__22847\ : std_logic;
signal \N__22846\ : std_logic;
signal \N__22843\ : std_logic;
signal \N__22842\ : std_logic;
signal \N__22839\ : std_logic;
signal \N__22836\ : std_logic;
signal \N__22835\ : std_logic;
signal \N__22830\ : std_logic;
signal \N__22829\ : std_logic;
signal \N__22826\ : std_logic;
signal \N__22823\ : std_logic;
signal \N__22820\ : std_logic;
signal \N__22819\ : std_logic;
signal \N__22818\ : std_logic;
signal \N__22815\ : std_logic;
signal \N__22812\ : std_logic;
signal \N__22809\ : std_logic;
signal \N__22806\ : std_logic;
signal \N__22803\ : std_logic;
signal \N__22802\ : std_logic;
signal \N__22799\ : std_logic;
signal \N__22794\ : std_logic;
signal \N__22793\ : std_logic;
signal \N__22790\ : std_logic;
signal \N__22787\ : std_logic;
signal \N__22784\ : std_logic;
signal \N__22779\ : std_logic;
signal \N__22776\ : std_logic;
signal \N__22771\ : std_logic;
signal \N__22768\ : std_logic;
signal \N__22765\ : std_logic;
signal \N__22764\ : std_logic;
signal \N__22761\ : std_logic;
signal \N__22758\ : std_logic;
signal \N__22755\ : std_logic;
signal \N__22748\ : std_logic;
signal \N__22741\ : std_logic;
signal \N__22738\ : std_logic;
signal \N__22735\ : std_logic;
signal \N__22726\ : std_logic;
signal \N__22723\ : std_logic;
signal \N__22714\ : std_logic;
signal \N__22711\ : std_logic;
signal \N__22708\ : std_logic;
signal \N__22705\ : std_logic;
signal \N__22702\ : std_logic;
signal \N__22699\ : std_logic;
signal \N__22696\ : std_logic;
signal \N__22693\ : std_logic;
signal \N__22690\ : std_logic;
signal \N__22689\ : std_logic;
signal \N__22688\ : std_logic;
signal \N__22685\ : std_logic;
signal \N__22684\ : std_logic;
signal \N__22681\ : std_logic;
signal \N__22678\ : std_logic;
signal \N__22677\ : std_logic;
signal \N__22676\ : std_logic;
signal \N__22675\ : std_logic;
signal \N__22672\ : std_logic;
signal \N__22669\ : std_logic;
signal \N__22668\ : std_logic;
signal \N__22665\ : std_logic;
signal \N__22662\ : std_logic;
signal \N__22659\ : std_logic;
signal \N__22656\ : std_logic;
signal \N__22655\ : std_logic;
signal \N__22654\ : std_logic;
signal \N__22651\ : std_logic;
signal \N__22650\ : std_logic;
signal \N__22649\ : std_logic;
signal \N__22644\ : std_logic;
signal \N__22641\ : std_logic;
signal \N__22640\ : std_logic;
signal \N__22633\ : std_logic;
signal \N__22630\ : std_logic;
signal \N__22627\ : std_logic;
signal \N__22624\ : std_logic;
signal \N__22623\ : std_logic;
signal \N__22622\ : std_logic;
signal \N__22621\ : std_logic;
signal \N__22620\ : std_logic;
signal \N__22619\ : std_logic;
signal \N__22616\ : std_logic;
signal \N__22613\ : std_logic;
signal \N__22610\ : std_logic;
signal \N__22609\ : std_logic;
signal \N__22604\ : std_logic;
signal \N__22601\ : std_logic;
signal \N__22600\ : std_logic;
signal \N__22593\ : std_logic;
signal \N__22590\ : std_logic;
signal \N__22587\ : std_logic;
signal \N__22584\ : std_logic;
signal \N__22583\ : std_logic;
signal \N__22582\ : std_logic;
signal \N__22581\ : std_logic;
signal \N__22580\ : std_logic;
signal \N__22579\ : std_logic;
signal \N__22578\ : std_logic;
signal \N__22575\ : std_logic;
signal \N__22574\ : std_logic;
signal \N__22573\ : std_logic;
signal \N__22572\ : std_logic;
signal \N__22569\ : std_logic;
signal \N__22566\ : std_logic;
signal \N__22565\ : std_logic;
signal \N__22564\ : std_logic;
signal \N__22563\ : std_logic;
signal \N__22562\ : std_logic;
signal \N__22561\ : std_logic;
signal \N__22560\ : std_logic;
signal \N__22555\ : std_logic;
signal \N__22552\ : std_logic;
signal \N__22549\ : std_logic;
signal \N__22548\ : std_logic;
signal \N__22547\ : std_logic;
signal \N__22542\ : std_logic;
signal \N__22539\ : std_logic;
signal \N__22538\ : std_logic;
signal \N__22537\ : std_logic;
signal \N__22536\ : std_logic;
signal \N__22535\ : std_logic;
signal \N__22534\ : std_logic;
signal \N__22533\ : std_logic;
signal \N__22526\ : std_logic;
signal \N__22523\ : std_logic;
signal \N__22520\ : std_logic;
signal \N__22517\ : std_logic;
signal \N__22516\ : std_logic;
signal \N__22515\ : std_logic;
signal \N__22514\ : std_logic;
signal \N__22513\ : std_logic;
signal \N__22512\ : std_logic;
signal \N__22509\ : std_logic;
signal \N__22506\ : std_logic;
signal \N__22503\ : std_logic;
signal \N__22500\ : std_logic;
signal \N__22499\ : std_logic;
signal \N__22498\ : std_logic;
signal \N__22495\ : std_logic;
signal \N__22492\ : std_logic;
signal \N__22489\ : std_logic;
signal \N__22488\ : std_logic;
signal \N__22487\ : std_logic;
signal \N__22486\ : std_logic;
signal \N__22483\ : std_logic;
signal \N__22478\ : std_logic;
signal \N__22475\ : std_logic;
signal \N__22474\ : std_logic;
signal \N__22471\ : std_logic;
signal \N__22470\ : std_logic;
signal \N__22467\ : std_logic;
signal \N__22466\ : std_logic;
signal \N__22465\ : std_logic;
signal \N__22462\ : std_logic;
signal \N__22459\ : std_logic;
signal \N__22456\ : std_logic;
signal \N__22449\ : std_logic;
signal \N__22446\ : std_logic;
signal \N__22445\ : std_logic;
signal \N__22444\ : std_logic;
signal \N__22441\ : std_logic;
signal \N__22440\ : std_logic;
signal \N__22439\ : std_logic;
signal \N__22438\ : std_logic;
signal \N__22437\ : std_logic;
signal \N__22436\ : std_logic;
signal \N__22435\ : std_logic;
signal \N__22434\ : std_logic;
signal \N__22429\ : std_logic;
signal \N__22426\ : std_logic;
signal \N__22423\ : std_logic;
signal \N__22422\ : std_logic;
signal \N__22421\ : std_logic;
signal \N__22420\ : std_logic;
signal \N__22419\ : std_logic;
signal \N__22416\ : std_logic;
signal \N__22413\ : std_logic;
signal \N__22410\ : std_logic;
signal \N__22409\ : std_logic;
signal \N__22408\ : std_logic;
signal \N__22407\ : std_logic;
signal \N__22404\ : std_logic;
signal \N__22397\ : std_logic;
signal \N__22394\ : std_logic;
signal \N__22391\ : std_logic;
signal \N__22388\ : std_logic;
signal \N__22387\ : std_logic;
signal \N__22386\ : std_logic;
signal \N__22383\ : std_logic;
signal \N__22380\ : std_logic;
signal \N__22377\ : std_logic;
signal \N__22374\ : std_logic;
signal \N__22371\ : std_logic;
signal \N__22366\ : std_logic;
signal \N__22363\ : std_logic;
signal \N__22360\ : std_logic;
signal \N__22353\ : std_logic;
signal \N__22352\ : std_logic;
signal \N__22349\ : std_logic;
signal \N__22348\ : std_logic;
signal \N__22347\ : std_logic;
signal \N__22344\ : std_logic;
signal \N__22341\ : std_logic;
signal \N__22340\ : std_logic;
signal \N__22337\ : std_logic;
signal \N__22332\ : std_logic;
signal \N__22329\ : std_logic;
signal \N__22326\ : std_logic;
signal \N__22323\ : std_logic;
signal \N__22322\ : std_logic;
signal \N__22319\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22315\ : std_logic;
signal \N__22314\ : std_logic;
signal \N__22311\ : std_logic;
signal \N__22308\ : std_logic;
signal \N__22303\ : std_logic;
signal \N__22298\ : std_logic;
signal \N__22295\ : std_logic;
signal \N__22292\ : std_logic;
signal \N__22289\ : std_logic;
signal \N__22286\ : std_logic;
signal \N__22283\ : std_logic;
signal \N__22282\ : std_logic;
signal \N__22279\ : std_logic;
signal \N__22276\ : std_logic;
signal \N__22273\ : std_logic;
signal \N__22270\ : std_logic;
signal \N__22267\ : std_logic;
signal \N__22266\ : std_logic;
signal \N__22263\ : std_logic;
signal \N__22258\ : std_logic;
signal \N__22255\ : std_logic;
signal \N__22252\ : std_logic;
signal \N__22249\ : std_logic;
signal \N__22248\ : std_logic;
signal \N__22247\ : std_logic;
signal \N__22244\ : std_logic;
signal \N__22243\ : std_logic;
signal \N__22240\ : std_logic;
signal \N__22239\ : std_logic;
signal \N__22234\ : std_logic;
signal \N__22231\ : std_logic;
signal \N__22230\ : std_logic;
signal \N__22229\ : std_logic;
signal \N__22226\ : std_logic;
signal \N__22225\ : std_logic;
signal \N__22222\ : std_logic;
signal \N__22219\ : std_logic;
signal \N__22212\ : std_logic;
signal \N__22209\ : std_logic;
signal \N__22206\ : std_logic;
signal \N__22205\ : std_logic;
signal \N__22202\ : std_logic;
signal \N__22199\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22193\ : std_logic;
signal \N__22180\ : std_logic;
signal \N__22177\ : std_logic;
signal \N__22174\ : std_logic;
signal \N__22171\ : std_logic;
signal \N__22168\ : std_logic;
signal \N__22165\ : std_logic;
signal \N__22162\ : std_logic;
signal \N__22159\ : std_logic;
signal \N__22154\ : std_logic;
signal \N__22151\ : std_logic;
signal \N__22146\ : std_logic;
signal \N__22143\ : std_logic;
signal \N__22140\ : std_logic;
signal \N__22137\ : std_logic;
signal \N__22134\ : std_logic;
signal \N__22131\ : std_logic;
signal \N__22128\ : std_logic;
signal \N__22117\ : std_logic;
signal \N__22112\ : std_logic;
signal \N__22109\ : std_logic;
signal \N__22106\ : std_logic;
signal \N__22101\ : std_logic;
signal \N__22096\ : std_logic;
signal \N__22093\ : std_logic;
signal \N__22090\ : std_logic;
signal \N__22083\ : std_logic;
signal \N__22080\ : std_logic;
signal \N__22077\ : std_logic;
signal \N__22074\ : std_logic;
signal \N__22071\ : std_logic;
signal \N__22070\ : std_logic;
signal \N__22069\ : std_logic;
signal \N__22066\ : std_logic;
signal \N__22063\ : std_logic;
signal \N__22062\ : std_logic;
signal \N__22061\ : std_logic;
signal \N__22058\ : std_logic;
signal \N__22055\ : std_logic;
signal \N__22050\ : std_logic;
signal \N__22047\ : std_logic;
signal \N__22044\ : std_logic;
signal \N__22041\ : std_logic;
signal \N__22038\ : std_logic;
signal \N__22037\ : std_logic;
signal \N__22034\ : std_logic;
signal \N__22031\ : std_logic;
signal \N__22024\ : std_logic;
signal \N__22021\ : std_logic;
signal \N__22020\ : std_logic;
signal \N__22017\ : std_logic;
signal \N__22006\ : std_logic;
signal \N__21999\ : std_logic;
signal \N__21992\ : std_logic;
signal \N__21985\ : std_logic;
signal \N__21982\ : std_logic;
signal \N__21977\ : std_logic;
signal \N__21972\ : std_logic;
signal \N__21965\ : std_logic;
signal \N__21960\ : std_logic;
signal \N__21959\ : std_logic;
signal \N__21958\ : std_logic;
signal \N__21949\ : std_logic;
signal \N__21938\ : std_logic;
signal \N__21935\ : std_logic;
signal \N__21932\ : std_logic;
signal \N__21927\ : std_logic;
signal \N__21924\ : std_logic;
signal \N__21921\ : std_logic;
signal \N__21918\ : std_logic;
signal \N__21915\ : std_logic;
signal \N__21908\ : std_logic;
signal \N__21903\ : std_logic;
signal \N__21900\ : std_logic;
signal \N__21897\ : std_logic;
signal \N__21894\ : std_logic;
signal \N__21891\ : std_logic;
signal \N__21888\ : std_logic;
signal \N__21885\ : std_logic;
signal \N__21882\ : std_logic;
signal \N__21875\ : std_logic;
signal \N__21870\ : std_logic;
signal \N__21865\ : std_logic;
signal \N__21860\ : std_logic;
signal \N__21857\ : std_logic;
signal \N__21854\ : std_logic;
signal \N__21845\ : std_logic;
signal \N__21838\ : std_logic;
signal \N__21833\ : std_logic;
signal \N__21830\ : std_logic;
signal \N__21825\ : std_logic;
signal \N__21820\ : std_logic;
signal \N__21815\ : std_logic;
signal \N__21812\ : std_logic;
signal \N__21809\ : std_logic;
signal \N__21806\ : std_logic;
signal \N__21801\ : std_logic;
signal \N__21798\ : std_logic;
signal \N__21793\ : std_logic;
signal \N__21788\ : std_logic;
signal \N__21785\ : std_logic;
signal \N__21780\ : std_logic;
signal \N__21773\ : std_logic;
signal \N__21768\ : std_logic;
signal \N__21765\ : std_logic;
signal \N__21762\ : std_logic;
signal \N__21757\ : std_logic;
signal \N__21752\ : std_logic;
signal \N__21739\ : std_logic;
signal \N__21736\ : std_logic;
signal \N__21733\ : std_logic;
signal \N__21730\ : std_logic;
signal \N__21727\ : std_logic;
signal \N__21724\ : std_logic;
signal \N__21721\ : std_logic;
signal \N__21718\ : std_logic;
signal \N__21715\ : std_logic;
signal \N__21712\ : std_logic;
signal \N__21709\ : std_logic;
signal \N__21706\ : std_logic;
signal \N__21703\ : std_logic;
signal \N__21700\ : std_logic;
signal \N__21697\ : std_logic;
signal \N__21694\ : std_logic;
signal \N__21691\ : std_logic;
signal \N__21688\ : std_logic;
signal \N__21685\ : std_logic;
signal \N__21682\ : std_logic;
signal \N__21679\ : std_logic;
signal \N__21676\ : std_logic;
signal \N__21673\ : std_logic;
signal \N__21670\ : std_logic;
signal \N__21667\ : std_logic;
signal \N__21664\ : std_logic;
signal \N__21661\ : std_logic;
signal \N__21658\ : std_logic;
signal \N__21655\ : std_logic;
signal \N__21652\ : std_logic;
signal \N__21649\ : std_logic;
signal \N__21646\ : std_logic;
signal \N__21643\ : std_logic;
signal \N__21640\ : std_logic;
signal \N__21637\ : std_logic;
signal \N__21634\ : std_logic;
signal \N__21631\ : std_logic;
signal \N__21628\ : std_logic;
signal \N__21625\ : std_logic;
signal \N__21622\ : std_logic;
signal \N__21619\ : std_logic;
signal \N__21616\ : std_logic;
signal \N__21613\ : std_logic;
signal \N__21610\ : std_logic;
signal \N__21607\ : std_logic;
signal \N__21604\ : std_logic;
signal \N__21601\ : std_logic;
signal \N__21598\ : std_logic;
signal \N__21595\ : std_logic;
signal \N__21592\ : std_logic;
signal \N__21589\ : std_logic;
signal \N__21586\ : std_logic;
signal \N__21583\ : std_logic;
signal \N__21580\ : std_logic;
signal \N__21577\ : std_logic;
signal \N__21574\ : std_logic;
signal \N__21571\ : std_logic;
signal \N__21568\ : std_logic;
signal \N__21565\ : std_logic;
signal \N__21562\ : std_logic;
signal \N__21559\ : std_logic;
signal \N__21556\ : std_logic;
signal \N__21553\ : std_logic;
signal \N__21550\ : std_logic;
signal \N__21547\ : std_logic;
signal \N__21544\ : std_logic;
signal \N__21541\ : std_logic;
signal \N__21538\ : std_logic;
signal \N__21535\ : std_logic;
signal \N__21532\ : std_logic;
signal \N__21529\ : std_logic;
signal \N__21526\ : std_logic;
signal \N__21523\ : std_logic;
signal \N__21520\ : std_logic;
signal \N__21517\ : std_logic;
signal \N__21514\ : std_logic;
signal \N__21511\ : std_logic;
signal \N__21508\ : std_logic;
signal \N__21505\ : std_logic;
signal \N__21502\ : std_logic;
signal \N__21499\ : std_logic;
signal \N__21496\ : std_logic;
signal \N__21493\ : std_logic;
signal \N__21490\ : std_logic;
signal \N__21489\ : std_logic;
signal \N__21488\ : std_logic;
signal \N__21487\ : std_logic;
signal \N__21484\ : std_logic;
signal \N__21481\ : std_logic;
signal \N__21480\ : std_logic;
signal \N__21477\ : std_logic;
signal \N__21474\ : std_logic;
signal \N__21473\ : std_logic;
signal \N__21468\ : std_logic;
signal \N__21465\ : std_logic;
signal \N__21464\ : std_logic;
signal \N__21463\ : std_logic;
signal \N__21460\ : std_logic;
signal \N__21459\ : std_logic;
signal \N__21458\ : std_logic;
signal \N__21457\ : std_logic;
signal \N__21456\ : std_logic;
signal \N__21453\ : std_logic;
signal \N__21450\ : std_logic;
signal \N__21447\ : std_logic;
signal \N__21444\ : std_logic;
signal \N__21441\ : std_logic;
signal \N__21438\ : std_logic;
signal \N__21437\ : std_logic;
signal \N__21436\ : std_logic;
signal \N__21433\ : std_logic;
signal \N__21430\ : std_logic;
signal \N__21427\ : std_logic;
signal \N__21424\ : std_logic;
signal \N__21421\ : std_logic;
signal \N__21416\ : std_logic;
signal \N__21409\ : std_logic;
signal \N__21406\ : std_logic;
signal \N__21403\ : std_logic;
signal \N__21400\ : std_logic;
signal \N__21395\ : std_logic;
signal \N__21392\ : std_logic;
signal \N__21389\ : std_logic;
signal \N__21386\ : std_logic;
signal \N__21379\ : std_logic;
signal \N__21374\ : std_logic;
signal \N__21371\ : std_logic;
signal \N__21368\ : std_logic;
signal \N__21365\ : std_logic;
signal \N__21360\ : std_logic;
signal \N__21357\ : std_logic;
signal \N__21346\ : std_logic;
signal \N__21345\ : std_logic;
signal \N__21344\ : std_logic;
signal \N__21343\ : std_logic;
signal \N__21342\ : std_logic;
signal \N__21341\ : std_logic;
signal \N__21340\ : std_logic;
signal \N__21339\ : std_logic;
signal \N__21338\ : std_logic;
signal \N__21337\ : std_logic;
signal \N__21336\ : std_logic;
signal \N__21335\ : std_logic;
signal \N__21332\ : std_logic;
signal \N__21329\ : std_logic;
signal \N__21326\ : std_logic;
signal \N__21325\ : std_logic;
signal \N__21324\ : std_logic;
signal \N__21323\ : std_logic;
signal \N__21322\ : std_logic;
signal \N__21321\ : std_logic;
signal \N__21318\ : std_logic;
signal \N__21317\ : std_logic;
signal \N__21314\ : std_logic;
signal \N__21311\ : std_logic;
signal \N__21308\ : std_logic;
signal \N__21307\ : std_logic;
signal \N__21306\ : std_logic;
signal \N__21303\ : std_logic;
signal \N__21300\ : std_logic;
signal \N__21297\ : std_logic;
signal \N__21296\ : std_logic;
signal \N__21295\ : std_logic;
signal \N__21294\ : std_logic;
signal \N__21293\ : std_logic;
signal \N__21292\ : std_logic;
signal \N__21289\ : std_logic;
signal \N__21288\ : std_logic;
signal \N__21285\ : std_logic;
signal \N__21282\ : std_logic;
signal \N__21281\ : std_logic;
signal \N__21280\ : std_logic;
signal \N__21279\ : std_logic;
signal \N__21278\ : std_logic;
signal \N__21273\ : std_logic;
signal \N__21270\ : std_logic;
signal \N__21269\ : std_logic;
signal \N__21268\ : std_logic;
signal \N__21267\ : std_logic;
signal \N__21266\ : std_logic;
signal \N__21263\ : std_logic;
signal \N__21262\ : std_logic;
signal \N__21261\ : std_logic;
signal \N__21260\ : std_logic;
signal \N__21259\ : std_logic;
signal \N__21256\ : std_logic;
signal \N__21253\ : std_logic;
signal \N__21252\ : std_logic;
signal \N__21251\ : std_logic;
signal \N__21248\ : std_logic;
signal \N__21245\ : std_logic;
signal \N__21242\ : std_logic;
signal \N__21237\ : std_logic;
signal \N__21234\ : std_logic;
signal \N__21231\ : std_logic;
signal \N__21228\ : std_logic;
signal \N__21225\ : std_logic;
signal \N__21220\ : std_logic;
signal \N__21219\ : std_logic;
signal \N__21218\ : std_logic;
signal \N__21217\ : std_logic;
signal \N__21214\ : std_logic;
signal \N__21211\ : std_logic;
signal \N__21210\ : std_logic;
signal \N__21209\ : std_logic;
signal \N__21206\ : std_logic;
signal \N__21203\ : std_logic;
signal \N__21200\ : std_logic;
signal \N__21199\ : std_logic;
signal \N__21198\ : std_logic;
signal \N__21197\ : std_logic;
signal \N__21196\ : std_logic;
signal \N__21195\ : std_logic;
signal \N__21194\ : std_logic;
signal \N__21191\ : std_logic;
signal \N__21188\ : std_logic;
signal \N__21185\ : std_logic;
signal \N__21182\ : std_logic;
signal \N__21181\ : std_logic;
signal \N__21180\ : std_logic;
signal \N__21179\ : std_logic;
signal \N__21176\ : std_logic;
signal \N__21173\ : std_logic;
signal \N__21172\ : std_logic;
signal \N__21171\ : std_logic;
signal \N__21168\ : std_logic;
signal \N__21167\ : std_logic;
signal \N__21166\ : std_logic;
signal \N__21163\ : std_logic;
signal \N__21158\ : std_logic;
signal \N__21155\ : std_logic;
signal \N__21152\ : std_logic;
signal \N__21151\ : std_logic;
signal \N__21148\ : std_logic;
signal \N__21147\ : std_logic;
signal \N__21144\ : std_logic;
signal \N__21141\ : std_logic;
signal \N__21138\ : std_logic;
signal \N__21135\ : std_logic;
signal \N__21132\ : std_logic;
signal \N__21129\ : std_logic;
signal \N__21124\ : std_logic;
signal \N__21121\ : std_logic;
signal \N__21118\ : std_logic;
signal \N__21115\ : std_logic;
signal \N__21108\ : std_logic;
signal \N__21097\ : std_logic;
signal \N__21094\ : std_logic;
signal \N__21093\ : std_logic;
signal \N__21092\ : std_logic;
signal \N__21087\ : std_logic;
signal \N__21084\ : std_logic;
signal \N__21081\ : std_logic;
signal \N__21078\ : std_logic;
signal \N__21063\ : std_logic;
signal \N__21060\ : std_logic;
signal \N__21057\ : std_logic;
signal \N__21056\ : std_logic;
signal \N__21055\ : std_logic;
signal \N__21052\ : std_logic;
signal \N__21049\ : std_logic;
signal \N__21046\ : std_logic;
signal \N__21041\ : std_logic;
signal \N__21038\ : std_logic;
signal \N__21037\ : std_logic;
signal \N__21036\ : std_logic;
signal \N__21035\ : std_logic;
signal \N__21034\ : std_logic;
signal \N__21033\ : std_logic;
signal \N__21030\ : std_logic;
signal \N__21027\ : std_logic;
signal \N__21024\ : std_logic;
signal \N__21019\ : std_logic;
signal \N__21016\ : std_logic;
signal \N__21013\ : std_logic;
signal \N__21010\ : std_logic;
signal \N__21007\ : std_logic;
signal \N__21000\ : std_logic;
signal \N__20997\ : std_logic;
signal \N__20994\ : std_logic;
signal \N__20991\ : std_logic;
signal \N__20988\ : std_logic;
signal \N__20985\ : std_logic;
signal \N__20976\ : std_logic;
signal \N__20973\ : std_logic;
signal \N__20970\ : std_logic;
signal \N__20959\ : std_logic;
signal \N__20956\ : std_logic;
signal \N__20955\ : std_logic;
signal \N__20952\ : std_logic;
signal \N__20949\ : std_logic;
signal \N__20946\ : std_logic;
signal \N__20937\ : std_logic;
signal \N__20932\ : std_logic;
signal \N__20929\ : std_logic;
signal \N__20926\ : std_logic;
signal \N__20923\ : std_logic;
signal \N__20920\ : std_logic;
signal \N__20915\ : std_logic;
signal \N__20912\ : std_logic;
signal \N__20909\ : std_logic;
signal \N__20906\ : std_logic;
signal \N__20903\ : std_logic;
signal \N__20896\ : std_logic;
signal \N__20889\ : std_logic;
signal \N__20886\ : std_logic;
signal \N__20881\ : std_logic;
signal \N__20874\ : std_logic;
signal \N__20871\ : std_logic;
signal \N__20862\ : std_logic;
signal \N__20853\ : std_logic;
signal \N__20850\ : std_logic;
signal \N__20845\ : std_logic;
signal \N__20838\ : std_logic;
signal \N__20835\ : std_logic;
signal \N__20832\ : std_logic;
signal \N__20829\ : std_logic;
signal \N__20824\ : std_logic;
signal \N__20811\ : std_logic;
signal \N__20808\ : std_logic;
signal \N__20805\ : std_logic;
signal \N__20802\ : std_logic;
signal \N__20797\ : std_logic;
signal \N__20794\ : std_logic;
signal \N__20787\ : std_logic;
signal \N__20776\ : std_logic;
signal \N__20761\ : std_logic;
signal \N__20758\ : std_logic;
signal \N__20755\ : std_logic;
signal \N__20752\ : std_logic;
signal \N__20749\ : std_logic;
signal \N__20746\ : std_logic;
signal \N__20743\ : std_logic;
signal \N__20740\ : std_logic;
signal \N__20737\ : std_logic;
signal \N__20734\ : std_logic;
signal \N__20731\ : std_logic;
signal \N__20728\ : std_logic;
signal \N__20725\ : std_logic;
signal \N__20722\ : std_logic;
signal \N__20719\ : std_logic;
signal \N__20716\ : std_logic;
signal \N__20713\ : std_logic;
signal \N__20710\ : std_logic;
signal \N__20707\ : std_logic;
signal \N__20704\ : std_logic;
signal \N__20701\ : std_logic;
signal \N__20698\ : std_logic;
signal \N__20695\ : std_logic;
signal \N__20692\ : std_logic;
signal \N__20689\ : std_logic;
signal \N__20686\ : std_logic;
signal \N__20683\ : std_logic;
signal \N__20680\ : std_logic;
signal \N__20677\ : std_logic;
signal \N__20674\ : std_logic;
signal \N__20671\ : std_logic;
signal \N__20668\ : std_logic;
signal \N__20665\ : std_logic;
signal \N__20662\ : std_logic;
signal \N__20659\ : std_logic;
signal \N__20656\ : std_logic;
signal \N__20653\ : std_logic;
signal \N__20650\ : std_logic;
signal \N__20647\ : std_logic;
signal \N__20644\ : std_logic;
signal \N__20641\ : std_logic;
signal \N__20638\ : std_logic;
signal \N__20635\ : std_logic;
signal \N__20632\ : std_logic;
signal \N__20629\ : std_logic;
signal \N__20626\ : std_logic;
signal \N__20623\ : std_logic;
signal \N__20622\ : std_logic;
signal \N__20619\ : std_logic;
signal \N__20618\ : std_logic;
signal \N__20615\ : std_logic;
signal \N__20614\ : std_logic;
signal \N__20611\ : std_logic;
signal \N__20608\ : std_logic;
signal \N__20607\ : std_logic;
signal \N__20606\ : std_logic;
signal \N__20603\ : std_logic;
signal \N__20600\ : std_logic;
signal \N__20599\ : std_logic;
signal \N__20598\ : std_logic;
signal \N__20597\ : std_logic;
signal \N__20596\ : std_logic;
signal \N__20591\ : std_logic;
signal \N__20588\ : std_logic;
signal \N__20587\ : std_logic;
signal \N__20584\ : std_logic;
signal \N__20583\ : std_logic;
signal \N__20578\ : std_logic;
signal \N__20575\ : std_logic;
signal \N__20572\ : std_logic;
signal \N__20569\ : std_logic;
signal \N__20566\ : std_logic;
signal \N__20565\ : std_logic;
signal \N__20560\ : std_logic;
signal \N__20557\ : std_logic;
signal \N__20554\ : std_logic;
signal \N__20551\ : std_logic;
signal \N__20550\ : std_logic;
signal \N__20547\ : std_logic;
signal \N__20542\ : std_logic;
signal \N__20539\ : std_logic;
signal \N__20536\ : std_logic;
signal \N__20533\ : std_logic;
signal \N__20530\ : std_logic;
signal \N__20527\ : std_logic;
signal \N__20522\ : std_logic;
signal \N__20519\ : std_logic;
signal \N__20514\ : std_logic;
signal \N__20511\ : std_logic;
signal \N__20508\ : std_logic;
signal \N__20505\ : std_logic;
signal \N__20496\ : std_logic;
signal \N__20485\ : std_logic;
signal \N__20482\ : std_logic;
signal \N__20479\ : std_logic;
signal \N__20476\ : std_logic;
signal \N__20473\ : std_logic;
signal \N__20470\ : std_logic;
signal \N__20467\ : std_logic;
signal \N__20464\ : std_logic;
signal \N__20461\ : std_logic;
signal \N__20458\ : std_logic;
signal \N__20455\ : std_logic;
signal \N__20452\ : std_logic;
signal \N__20449\ : std_logic;
signal \N__20446\ : std_logic;
signal \N__20443\ : std_logic;
signal \N__20440\ : std_logic;
signal \N__20437\ : std_logic;
signal \N__20434\ : std_logic;
signal \N__20431\ : std_logic;
signal \N__20428\ : std_logic;
signal \N__20425\ : std_logic;
signal \N__20422\ : std_logic;
signal \N__20419\ : std_logic;
signal \N__20416\ : std_logic;
signal \N__20413\ : std_logic;
signal \N__20410\ : std_logic;
signal \N__20407\ : std_logic;
signal \N__20404\ : std_logic;
signal \N__20401\ : std_logic;
signal \N__20398\ : std_logic;
signal \N__20395\ : std_logic;
signal \N__20392\ : std_logic;
signal \N__20389\ : std_logic;
signal \N__20386\ : std_logic;
signal \N__20383\ : std_logic;
signal \N__20380\ : std_logic;
signal \N__20377\ : std_logic;
signal \N__20374\ : std_logic;
signal \N__20371\ : std_logic;
signal \N__20368\ : std_logic;
signal \N__20365\ : std_logic;
signal \N__20362\ : std_logic;
signal \N__20359\ : std_logic;
signal \N__20356\ : std_logic;
signal \N__20353\ : std_logic;
signal \N__20350\ : std_logic;
signal \N__20347\ : std_logic;
signal \N__20344\ : std_logic;
signal \N__20341\ : std_logic;
signal \N__20338\ : std_logic;
signal \N__20335\ : std_logic;
signal \N__20332\ : std_logic;
signal \N__20329\ : std_logic;
signal \N__20326\ : std_logic;
signal \N__20323\ : std_logic;
signal \N__20320\ : std_logic;
signal \N__20317\ : std_logic;
signal \N__20314\ : std_logic;
signal \N__20311\ : std_logic;
signal \N__20308\ : std_logic;
signal \N__20305\ : std_logic;
signal \N__20302\ : std_logic;
signal \N__20299\ : std_logic;
signal \N__20296\ : std_logic;
signal \N__20293\ : std_logic;
signal \N__20290\ : std_logic;
signal \N__20287\ : std_logic;
signal \N__20284\ : std_logic;
signal \N__20281\ : std_logic;
signal \N__20278\ : std_logic;
signal \N__20275\ : std_logic;
signal \N__20274\ : std_logic;
signal \N__20271\ : std_logic;
signal \N__20268\ : std_logic;
signal \N__20265\ : std_logic;
signal \N__20260\ : std_logic;
signal \N__20259\ : std_logic;
signal \N__20256\ : std_logic;
signal \N__20253\ : std_logic;
signal \N__20250\ : std_logic;
signal \N__20245\ : std_logic;
signal \N__20242\ : std_logic;
signal \N__20241\ : std_logic;
signal \N__20240\ : std_logic;
signal \N__20239\ : std_logic;
signal \N__20236\ : std_logic;
signal \N__20233\ : std_logic;
signal \N__20230\ : std_logic;
signal \N__20229\ : std_logic;
signal \N__20228\ : std_logic;
signal \N__20225\ : std_logic;
signal \N__20220\ : std_logic;
signal \N__20217\ : std_logic;
signal \N__20216\ : std_logic;
signal \N__20215\ : std_logic;
signal \N__20210\ : std_logic;
signal \N__20209\ : std_logic;
signal \N__20202\ : std_logic;
signal \N__20199\ : std_logic;
signal \N__20198\ : std_logic;
signal \N__20197\ : std_logic;
signal \N__20196\ : std_logic;
signal \N__20195\ : std_logic;
signal \N__20194\ : std_logic;
signal \N__20193\ : std_logic;
signal \N__20192\ : std_logic;
signal \N__20191\ : std_logic;
signal \N__20188\ : std_logic;
signal \N__20185\ : std_logic;
signal \N__20182\ : std_logic;
signal \N__20179\ : std_logic;
signal \N__20176\ : std_logic;
signal \N__20171\ : std_logic;
signal \N__20170\ : std_logic;
signal \N__20169\ : std_logic;
signal \N__20168\ : std_logic;
signal \N__20167\ : std_logic;
signal \N__20166\ : std_logic;
signal \N__20153\ : std_logic;
signal \N__20150\ : std_logic;
signal \N__20139\ : std_logic;
signal \N__20132\ : std_logic;
signal \N__20127\ : std_logic;
signal \N__20116\ : std_logic;
signal \N__20115\ : std_logic;
signal \N__20112\ : std_logic;
signal \N__20109\ : std_logic;
signal \N__20106\ : std_logic;
signal \N__20103\ : std_logic;
signal \N__20100\ : std_logic;
signal \N__20097\ : std_logic;
signal \N__20094\ : std_logic;
signal \N__20091\ : std_logic;
signal \N__20088\ : std_logic;
signal \N__20085\ : std_logic;
signal \N__20082\ : std_logic;
signal \N__20079\ : std_logic;
signal \N__20076\ : std_logic;
signal \N__20073\ : std_logic;
signal \N__20070\ : std_logic;
signal \N__20067\ : std_logic;
signal \N__20064\ : std_logic;
signal \N__20061\ : std_logic;
signal \N__20058\ : std_logic;
signal \N__20055\ : std_logic;
signal \N__20052\ : std_logic;
signal \N__20049\ : std_logic;
signal \N__20046\ : std_logic;
signal \N__20043\ : std_logic;
signal \N__20040\ : std_logic;
signal \N__20037\ : std_logic;
signal \N__20034\ : std_logic;
signal \N__20031\ : std_logic;
signal \N__20028\ : std_logic;
signal \N__20025\ : std_logic;
signal \N__20022\ : std_logic;
signal \N__20019\ : std_logic;
signal \N__20016\ : std_logic;
signal \N__20013\ : std_logic;
signal \N__20010\ : std_logic;
signal \N__20007\ : std_logic;
signal \N__20004\ : std_logic;
signal \N__20001\ : std_logic;
signal \N__19998\ : std_logic;
signal \N__19995\ : std_logic;
signal \N__19992\ : std_logic;
signal \N__19989\ : std_logic;
signal \N__19986\ : std_logic;
signal \N__19983\ : std_logic;
signal \N__19980\ : std_logic;
signal \N__19977\ : std_logic;
signal \N__19974\ : std_logic;
signal \N__19971\ : std_logic;
signal \N__19968\ : std_logic;
signal \N__19965\ : std_logic;
signal \N__19962\ : std_logic;
signal \N__19959\ : std_logic;
signal \N__19956\ : std_logic;
signal \N__19953\ : std_logic;
signal \N__19950\ : std_logic;
signal \N__19947\ : std_logic;
signal \N__19944\ : std_logic;
signal \N__19941\ : std_logic;
signal \N__19938\ : std_logic;
signal \N__19935\ : std_logic;
signal \N__19932\ : std_logic;
signal \N__19929\ : std_logic;
signal \N__19926\ : std_logic;
signal \N__19923\ : std_logic;
signal \N__19920\ : std_logic;
signal \N__19917\ : std_logic;
signal \N__19912\ : std_logic;
signal \N__19909\ : std_logic;
signal \N__19906\ : std_logic;
signal \N__19903\ : std_logic;
signal \N__19900\ : std_logic;
signal \N__19897\ : std_logic;
signal \N__19894\ : std_logic;
signal \N__19891\ : std_logic;
signal \N__19888\ : std_logic;
signal \N__19885\ : std_logic;
signal \N__19882\ : std_logic;
signal \N__19881\ : std_logic;
signal \N__19878\ : std_logic;
signal \N__19877\ : std_logic;
signal \N__19876\ : std_logic;
signal \N__19875\ : std_logic;
signal \N__19874\ : std_logic;
signal \N__19871\ : std_logic;
signal \N__19870\ : std_logic;
signal \N__19869\ : std_logic;
signal \N__19866\ : std_logic;
signal \N__19863\ : std_logic;
signal \N__19860\ : std_logic;
signal \N__19857\ : std_logic;
signal \N__19854\ : std_logic;
signal \N__19853\ : std_logic;
signal \N__19850\ : std_logic;
signal \N__19847\ : std_logic;
signal \N__19844\ : std_logic;
signal \N__19841\ : std_logic;
signal \N__19836\ : std_logic;
signal \N__19831\ : std_logic;
signal \N__19828\ : std_logic;
signal \N__19825\ : std_logic;
signal \N__19822\ : std_logic;
signal \N__19819\ : std_logic;
signal \N__19814\ : std_logic;
signal \N__19809\ : std_logic;
signal \N__19804\ : std_logic;
signal \N__19799\ : std_logic;
signal \N__19796\ : std_logic;
signal \N__19789\ : std_logic;
signal \N__19786\ : std_logic;
signal \N__19783\ : std_logic;
signal \N__19780\ : std_logic;
signal \N__19777\ : std_logic;
signal \N__19774\ : std_logic;
signal \N__19771\ : std_logic;
signal \N__19768\ : std_logic;
signal \N__19765\ : std_logic;
signal \N__19762\ : std_logic;
signal \N__19759\ : std_logic;
signal \N__19756\ : std_logic;
signal \N__19753\ : std_logic;
signal \N__19750\ : std_logic;
signal \N__19747\ : std_logic;
signal \N__19744\ : std_logic;
signal \N__19741\ : std_logic;
signal \N__19738\ : std_logic;
signal \N__19735\ : std_logic;
signal \N__19732\ : std_logic;
signal \N__19729\ : std_logic;
signal \N__19726\ : std_logic;
signal \N__19723\ : std_logic;
signal \N__19720\ : std_logic;
signal \N__19717\ : std_logic;
signal \N__19716\ : std_logic;
signal \N__19715\ : std_logic;
signal \N__19714\ : std_logic;
signal \N__19713\ : std_logic;
signal \N__19710\ : std_logic;
signal \N__19707\ : std_logic;
signal \N__19702\ : std_logic;
signal \N__19701\ : std_logic;
signal \N__19698\ : std_logic;
signal \N__19697\ : std_logic;
signal \N__19694\ : std_logic;
signal \N__19693\ : std_logic;
signal \N__19692\ : std_logic;
signal \N__19691\ : std_logic;
signal \N__19686\ : std_logic;
signal \N__19683\ : std_logic;
signal \N__19680\ : std_logic;
signal \N__19677\ : std_logic;
signal \N__19674\ : std_logic;
signal \N__19671\ : std_logic;
signal \N__19670\ : std_logic;
signal \N__19667\ : std_logic;
signal \N__19664\ : std_logic;
signal \N__19663\ : std_logic;
signal \N__19662\ : std_logic;
signal \N__19661\ : std_logic;
signal \N__19658\ : std_logic;
signal \N__19651\ : std_logic;
signal \N__19646\ : std_logic;
signal \N__19643\ : std_logic;
signal \N__19638\ : std_logic;
signal \N__19635\ : std_logic;
signal \N__19632\ : std_logic;
signal \N__19629\ : std_logic;
signal \N__19626\ : std_logic;
signal \N__19623\ : std_logic;
signal \N__19612\ : std_logic;
signal \N__19603\ : std_logic;
signal \N__19600\ : std_logic;
signal \N__19597\ : std_logic;
signal \N__19594\ : std_logic;
signal \N__19591\ : std_logic;
signal \N__19588\ : std_logic;
signal \N__19587\ : std_logic;
signal \N__19584\ : std_logic;
signal \N__19583\ : std_logic;
signal \N__19582\ : std_logic;
signal \N__19579\ : std_logic;
signal \N__19576\ : std_logic;
signal \N__19573\ : std_logic;
signal \N__19572\ : std_logic;
signal \N__19569\ : std_logic;
signal \N__19566\ : std_logic;
signal \N__19563\ : std_logic;
signal \N__19560\ : std_logic;
signal \N__19557\ : std_logic;
signal \N__19552\ : std_logic;
signal \N__19543\ : std_logic;
signal \N__19540\ : std_logic;
signal \N__19537\ : std_logic;
signal \N__19534\ : std_logic;
signal \N__19533\ : std_logic;
signal \N__19532\ : std_logic;
signal \N__19529\ : std_logic;
signal \N__19526\ : std_logic;
signal \N__19525\ : std_logic;
signal \N__19522\ : std_logic;
signal \N__19521\ : std_logic;
signal \N__19520\ : std_logic;
signal \N__19517\ : std_logic;
signal \N__19514\ : std_logic;
signal \N__19513\ : std_logic;
signal \N__19512\ : std_logic;
signal \N__19511\ : std_logic;
signal \N__19508\ : std_logic;
signal \N__19505\ : std_logic;
signal \N__19502\ : std_logic;
signal \N__19501\ : std_logic;
signal \N__19500\ : std_logic;
signal \N__19497\ : std_logic;
signal \N__19496\ : std_logic;
signal \N__19495\ : std_logic;
signal \N__19494\ : std_logic;
signal \N__19493\ : std_logic;
signal \N__19492\ : std_logic;
signal \N__19487\ : std_logic;
signal \N__19480\ : std_logic;
signal \N__19477\ : std_logic;
signal \N__19472\ : std_logic;
signal \N__19471\ : std_logic;
signal \N__19470\ : std_logic;
signal \N__19469\ : std_logic;
signal \N__19468\ : std_logic;
signal \N__19467\ : std_logic;
signal \N__19462\ : std_logic;
signal \N__19459\ : std_logic;
signal \N__19448\ : std_logic;
signal \N__19443\ : std_logic;
signal \N__19438\ : std_logic;
signal \N__19433\ : std_logic;
signal \N__19426\ : std_logic;
signal \N__19411\ : std_logic;
signal \N__19410\ : std_logic;
signal \N__19407\ : std_logic;
signal \N__19404\ : std_logic;
signal \N__19401\ : std_logic;
signal \N__19398\ : std_logic;
signal \N__19397\ : std_logic;
signal \N__19394\ : std_logic;
signal \N__19391\ : std_logic;
signal \N__19388\ : std_logic;
signal \N__19381\ : std_logic;
signal \N__19378\ : std_logic;
signal \N__19375\ : std_logic;
signal \N__19372\ : std_logic;
signal \N__19369\ : std_logic;
signal \N__19368\ : std_logic;
signal \N__19367\ : std_logic;
signal \N__19366\ : std_logic;
signal \N__19365\ : std_logic;
signal \N__19364\ : std_logic;
signal \N__19363\ : std_logic;
signal \N__19362\ : std_logic;
signal \N__19361\ : std_logic;
signal \N__19360\ : std_logic;
signal \N__19359\ : std_logic;
signal \N__19356\ : std_logic;
signal \N__19355\ : std_logic;
signal \N__19354\ : std_logic;
signal \N__19353\ : std_logic;
signal \N__19352\ : std_logic;
signal \N__19351\ : std_logic;
signal \N__19350\ : std_logic;
signal \N__19349\ : std_logic;
signal \N__19348\ : std_logic;
signal \N__19347\ : std_logic;
signal \N__19346\ : std_logic;
signal \N__19345\ : std_logic;
signal \N__19344\ : std_logic;
signal \N__19343\ : std_logic;
signal \N__19342\ : std_logic;
signal \N__19341\ : std_logic;
signal \N__19340\ : std_logic;
signal \N__19339\ : std_logic;
signal \N__19338\ : std_logic;
signal \N__19337\ : std_logic;
signal \N__19336\ : std_logic;
signal \N__19335\ : std_logic;
signal \N__19334\ : std_logic;
signal \N__19333\ : std_logic;
signal \N__19332\ : std_logic;
signal \N__19331\ : std_logic;
signal \N__19330\ : std_logic;
signal \N__19329\ : std_logic;
signal \N__19328\ : std_logic;
signal \N__19327\ : std_logic;
signal \N__19326\ : std_logic;
signal \N__19325\ : std_logic;
signal \N__19324\ : std_logic;
signal \N__19323\ : std_logic;
signal \N__19322\ : std_logic;
signal \N__19321\ : std_logic;
signal \N__19228\ : std_logic;
signal \N__19225\ : std_logic;
signal \N__19222\ : std_logic;
signal \N__19219\ : std_logic;
signal \N__19216\ : std_logic;
signal \N__19215\ : std_logic;
signal \N__19212\ : std_logic;
signal \N__19209\ : std_logic;
signal \N__19206\ : std_logic;
signal \N__19203\ : std_logic;
signal \N__19200\ : std_logic;
signal \N__19197\ : std_logic;
signal \N__19192\ : std_logic;
signal \N__19189\ : std_logic;
signal \N__19186\ : std_logic;
signal \N__19183\ : std_logic;
signal \N__19180\ : std_logic;
signal \N__19177\ : std_logic;
signal \N__19174\ : std_logic;
signal \N__19171\ : std_logic;
signal \N__19168\ : std_logic;
signal \N__19165\ : std_logic;
signal \N__19162\ : std_logic;
signal \N__19159\ : std_logic;
signal \N__19156\ : std_logic;
signal \N__19153\ : std_logic;
signal \N__19150\ : std_logic;
signal \N__19147\ : std_logic;
signal \N__19144\ : std_logic;
signal \N__19141\ : std_logic;
signal \N__19138\ : std_logic;
signal \N__19135\ : std_logic;
signal \N__19132\ : std_logic;
signal \N__19129\ : std_logic;
signal \N__19128\ : std_logic;
signal \N__19127\ : std_logic;
signal \N__19126\ : std_logic;
signal \N__19123\ : std_logic;
signal \N__19122\ : std_logic;
signal \N__19121\ : std_logic;
signal \N__19120\ : std_logic;
signal \N__19117\ : std_logic;
signal \N__19114\ : std_logic;
signal \N__19111\ : std_logic;
signal \N__19108\ : std_logic;
signal \N__19105\ : std_logic;
signal \N__19104\ : std_logic;
signal \N__19103\ : std_logic;
signal \N__19102\ : std_logic;
signal \N__19101\ : std_logic;
signal \N__19100\ : std_logic;
signal \N__19099\ : std_logic;
signal \N__19096\ : std_logic;
signal \N__19095\ : std_logic;
signal \N__19092\ : std_logic;
signal \N__19089\ : std_logic;
signal \N__19084\ : std_logic;
signal \N__19079\ : std_logic;
signal \N__19076\ : std_logic;
signal \N__19071\ : std_logic;
signal \N__19068\ : std_logic;
signal \N__19065\ : std_logic;
signal \N__19058\ : std_logic;
signal \N__19053\ : std_logic;
signal \N__19042\ : std_logic;
signal \N__19037\ : std_logic;
signal \N__19030\ : std_logic;
signal \N__19027\ : std_logic;
signal \N__19026\ : std_logic;
signal \N__19023\ : std_logic;
signal \N__19022\ : std_logic;
signal \N__19021\ : std_logic;
signal \N__19018\ : std_logic;
signal \N__19013\ : std_logic;
signal \N__19010\ : std_logic;
signal \N__19003\ : std_logic;
signal \N__19000\ : std_logic;
signal \N__18997\ : std_logic;
signal \N__18994\ : std_logic;
signal \N__18991\ : std_logic;
signal \N__18988\ : std_logic;
signal \N__18987\ : std_logic;
signal \N__18984\ : std_logic;
signal \N__18983\ : std_logic;
signal \N__18982\ : std_logic;
signal \N__18979\ : std_logic;
signal \N__18976\ : std_logic;
signal \N__18971\ : std_logic;
signal \N__18968\ : std_logic;
signal \N__18961\ : std_logic;
signal \N__18960\ : std_logic;
signal \N__18957\ : std_logic;
signal \N__18954\ : std_logic;
signal \N__18949\ : std_logic;
signal \N__18946\ : std_logic;
signal \N__18943\ : std_logic;
signal \N__18942\ : std_logic;
signal \N__18939\ : std_logic;
signal \N__18936\ : std_logic;
signal \N__18933\ : std_logic;
signal \N__18930\ : std_logic;
signal \N__18927\ : std_logic;
signal \N__18924\ : std_logic;
signal \N__18921\ : std_logic;
signal \N__18918\ : std_logic;
signal \N__18915\ : std_logic;
signal \N__18912\ : std_logic;
signal \N__18909\ : std_logic;
signal \N__18906\ : std_logic;
signal \N__18903\ : std_logic;
signal \N__18900\ : std_logic;
signal \N__18897\ : std_logic;
signal \N__18894\ : std_logic;
signal \N__18891\ : std_logic;
signal \N__18888\ : std_logic;
signal \N__18885\ : std_logic;
signal \N__18882\ : std_logic;
signal \N__18879\ : std_logic;
signal \N__18876\ : std_logic;
signal \N__18873\ : std_logic;
signal \N__18870\ : std_logic;
signal \N__18867\ : std_logic;
signal \N__18864\ : std_logic;
signal \N__18861\ : std_logic;
signal \N__18858\ : std_logic;
signal \N__18855\ : std_logic;
signal \N__18852\ : std_logic;
signal \N__18849\ : std_logic;
signal \N__18846\ : std_logic;
signal \N__18843\ : std_logic;
signal \N__18840\ : std_logic;
signal \N__18837\ : std_logic;
signal \N__18834\ : std_logic;
signal \N__18831\ : std_logic;
signal \N__18828\ : std_logic;
signal \N__18825\ : std_logic;
signal \N__18822\ : std_logic;
signal \N__18819\ : std_logic;
signal \N__18816\ : std_logic;
signal \N__18813\ : std_logic;
signal \N__18810\ : std_logic;
signal \N__18807\ : std_logic;
signal \N__18804\ : std_logic;
signal \N__18801\ : std_logic;
signal \N__18798\ : std_logic;
signal \N__18795\ : std_logic;
signal \N__18792\ : std_logic;
signal \N__18789\ : std_logic;
signal \N__18786\ : std_logic;
signal \N__18783\ : std_logic;
signal \N__18780\ : std_logic;
signal \N__18777\ : std_logic;
signal \N__18774\ : std_logic;
signal \N__18771\ : std_logic;
signal \N__18768\ : std_logic;
signal \N__18765\ : std_logic;
signal \N__18762\ : std_logic;
signal \N__18759\ : std_logic;
signal \N__18756\ : std_logic;
signal \N__18753\ : std_logic;
signal \N__18750\ : std_logic;
signal \N__18747\ : std_logic;
signal \N__18744\ : std_logic;
signal \N__18739\ : std_logic;
signal \N__18736\ : std_logic;
signal \N__18733\ : std_logic;
signal \N__18732\ : std_logic;
signal \N__18729\ : std_logic;
signal \N__18726\ : std_logic;
signal \N__18723\ : std_logic;
signal \N__18718\ : std_logic;
signal \N__18715\ : std_logic;
signal \N__18712\ : std_logic;
signal \N__18711\ : std_logic;
signal \N__18708\ : std_logic;
signal \N__18705\ : std_logic;
signal \N__18702\ : std_logic;
signal \N__18699\ : std_logic;
signal \N__18696\ : std_logic;
signal \N__18693\ : std_logic;
signal \N__18690\ : std_logic;
signal \N__18687\ : std_logic;
signal \N__18684\ : std_logic;
signal \N__18681\ : std_logic;
signal \N__18678\ : std_logic;
signal \N__18675\ : std_logic;
signal \N__18672\ : std_logic;
signal \N__18669\ : std_logic;
signal \N__18666\ : std_logic;
signal \N__18663\ : std_logic;
signal \N__18660\ : std_logic;
signal \N__18657\ : std_logic;
signal \N__18654\ : std_logic;
signal \N__18651\ : std_logic;
signal \N__18648\ : std_logic;
signal \N__18645\ : std_logic;
signal \N__18642\ : std_logic;
signal \N__18639\ : std_logic;
signal \N__18636\ : std_logic;
signal \N__18633\ : std_logic;
signal \N__18630\ : std_logic;
signal \N__18627\ : std_logic;
signal \N__18624\ : std_logic;
signal \N__18621\ : std_logic;
signal \N__18618\ : std_logic;
signal \N__18615\ : std_logic;
signal \N__18612\ : std_logic;
signal \N__18609\ : std_logic;
signal \N__18606\ : std_logic;
signal \N__18603\ : std_logic;
signal \N__18600\ : std_logic;
signal \N__18597\ : std_logic;
signal \N__18594\ : std_logic;
signal \N__18591\ : std_logic;
signal \N__18588\ : std_logic;
signal \N__18585\ : std_logic;
signal \N__18582\ : std_logic;
signal \N__18579\ : std_logic;
signal \N__18576\ : std_logic;
signal \N__18573\ : std_logic;
signal \N__18570\ : std_logic;
signal \N__18567\ : std_logic;
signal \N__18564\ : std_logic;
signal \N__18561\ : std_logic;
signal \N__18558\ : std_logic;
signal \N__18555\ : std_logic;
signal \N__18552\ : std_logic;
signal \N__18549\ : std_logic;
signal \N__18546\ : std_logic;
signal \N__18543\ : std_logic;
signal \N__18540\ : std_logic;
signal \N__18537\ : std_logic;
signal \N__18534\ : std_logic;
signal \N__18531\ : std_logic;
signal \N__18528\ : std_logic;
signal \N__18525\ : std_logic;
signal \N__18522\ : std_logic;
signal \N__18519\ : std_logic;
signal \N__18516\ : std_logic;
signal \N__18513\ : std_logic;
signal \N__18510\ : std_logic;
signal \N__18507\ : std_logic;
signal \N__18504\ : std_logic;
signal \N__18499\ : std_logic;
signal \N__18496\ : std_logic;
signal \N__18493\ : std_logic;
signal \N__18490\ : std_logic;
signal \N__18487\ : std_logic;
signal \N__18484\ : std_logic;
signal \N__18481\ : std_logic;
signal \N__18478\ : std_logic;
signal \N__18475\ : std_logic;
signal \N__18472\ : std_logic;
signal \N__18469\ : std_logic;
signal \N__18466\ : std_logic;
signal \N__18465\ : std_logic;
signal \N__18464\ : std_logic;
signal \N__18461\ : std_logic;
signal \N__18458\ : std_logic;
signal \N__18457\ : std_logic;
signal \N__18454\ : std_logic;
signal \N__18451\ : std_logic;
signal \N__18448\ : std_logic;
signal \N__18445\ : std_logic;
signal \N__18442\ : std_logic;
signal \N__18433\ : std_logic;
signal \N__18430\ : std_logic;
signal \N__18427\ : std_logic;
signal \N__18424\ : std_logic;
signal \N__18421\ : std_logic;
signal \N__18420\ : std_logic;
signal \N__18417\ : std_logic;
signal \N__18414\ : std_logic;
signal \N__18411\ : std_logic;
signal \N__18408\ : std_logic;
signal \N__18407\ : std_logic;
signal \N__18406\ : std_logic;
signal \N__18403\ : std_logic;
signal \N__18400\ : std_logic;
signal \N__18397\ : std_logic;
signal \N__18394\ : std_logic;
signal \N__18385\ : std_logic;
signal \N__18382\ : std_logic;
signal \N__18379\ : std_logic;
signal \N__18376\ : std_logic;
signal \N__18375\ : std_logic;
signal \N__18374\ : std_logic;
signal \N__18373\ : std_logic;
signal \N__18370\ : std_logic;
signal \N__18367\ : std_logic;
signal \N__18364\ : std_logic;
signal \N__18361\ : std_logic;
signal \N__18352\ : std_logic;
signal \N__18349\ : std_logic;
signal \N__18346\ : std_logic;
signal \N__18343\ : std_logic;
signal \N__18340\ : std_logic;
signal \N__18337\ : std_logic;
signal \N__18334\ : std_logic;
signal \N__18331\ : std_logic;
signal \N__18328\ : std_logic;
signal \N__18325\ : std_logic;
signal \N__18322\ : std_logic;
signal \N__18321\ : std_logic;
signal \N__18320\ : std_logic;
signal \N__18319\ : std_logic;
signal \N__18316\ : std_logic;
signal \N__18313\ : std_logic;
signal \N__18310\ : std_logic;
signal \N__18307\ : std_logic;
signal \N__18302\ : std_logic;
signal \N__18299\ : std_logic;
signal \N__18292\ : std_logic;
signal \N__18291\ : std_logic;
signal \N__18288\ : std_logic;
signal \N__18285\ : std_logic;
signal \N__18282\ : std_logic;
signal \N__18279\ : std_logic;
signal \N__18274\ : std_logic;
signal \N__18271\ : std_logic;
signal \N__18268\ : std_logic;
signal \N__18265\ : std_logic;
signal \N__18262\ : std_logic;
signal \N__18261\ : std_logic;
signal \N__18258\ : std_logic;
signal \N__18255\ : std_logic;
signal \N__18252\ : std_logic;
signal \N__18249\ : std_logic;
signal \N__18246\ : std_logic;
signal \N__18243\ : std_logic;
signal \N__18240\ : std_logic;
signal \N__18237\ : std_logic;
signal \N__18234\ : std_logic;
signal \N__18231\ : std_logic;
signal \N__18228\ : std_logic;
signal \N__18225\ : std_logic;
signal \N__18222\ : std_logic;
signal \N__18219\ : std_logic;
signal \N__18216\ : std_logic;
signal \N__18213\ : std_logic;
signal \N__18210\ : std_logic;
signal \N__18207\ : std_logic;
signal \N__18204\ : std_logic;
signal \N__18201\ : std_logic;
signal \N__18198\ : std_logic;
signal \N__18195\ : std_logic;
signal \N__18192\ : std_logic;
signal \N__18189\ : std_logic;
signal \N__18186\ : std_logic;
signal \N__18183\ : std_logic;
signal \N__18180\ : std_logic;
signal \N__18177\ : std_logic;
signal \N__18174\ : std_logic;
signal \N__18171\ : std_logic;
signal \N__18168\ : std_logic;
signal \N__18165\ : std_logic;
signal \N__18162\ : std_logic;
signal \N__18159\ : std_logic;
signal \N__18156\ : std_logic;
signal \N__18153\ : std_logic;
signal \N__18150\ : std_logic;
signal \N__18147\ : std_logic;
signal \N__18144\ : std_logic;
signal \N__18141\ : std_logic;
signal \N__18138\ : std_logic;
signal \N__18135\ : std_logic;
signal \N__18132\ : std_logic;
signal \N__18129\ : std_logic;
signal \N__18126\ : std_logic;
signal \N__18123\ : std_logic;
signal \N__18120\ : std_logic;
signal \N__18117\ : std_logic;
signal \N__18114\ : std_logic;
signal \N__18111\ : std_logic;
signal \N__18108\ : std_logic;
signal \N__18105\ : std_logic;
signal \N__18102\ : std_logic;
signal \N__18099\ : std_logic;
signal \N__18096\ : std_logic;
signal \N__18093\ : std_logic;
signal \N__18090\ : std_logic;
signal \N__18087\ : std_logic;
signal \N__18084\ : std_logic;
signal \N__18081\ : std_logic;
signal \N__18078\ : std_logic;
signal \N__18075\ : std_logic;
signal \N__18072\ : std_logic;
signal \N__18069\ : std_logic;
signal \N__18066\ : std_logic;
signal \N__18063\ : std_logic;
signal \N__18060\ : std_logic;
signal \N__18057\ : std_logic;
signal \N__18052\ : std_logic;
signal \N__18049\ : std_logic;
signal \N__18046\ : std_logic;
signal \N__18043\ : std_logic;
signal \N__18040\ : std_logic;
signal \N__18037\ : std_logic;
signal \N__18034\ : std_logic;
signal \N__18031\ : std_logic;
signal \N__18028\ : std_logic;
signal \N__18025\ : std_logic;
signal \N__18022\ : std_logic;
signal \N__18019\ : std_logic;
signal \N__18016\ : std_logic;
signal \N__18013\ : std_logic;
signal \N__18010\ : std_logic;
signal \N__18007\ : std_logic;
signal \N__18004\ : std_logic;
signal \N__18001\ : std_logic;
signal \N__17998\ : std_logic;
signal \N__17995\ : std_logic;
signal \N__17992\ : std_logic;
signal \N__17989\ : std_logic;
signal \N__17986\ : std_logic;
signal \N__17983\ : std_logic;
signal \N__17980\ : std_logic;
signal \N__17977\ : std_logic;
signal \N__17974\ : std_logic;
signal \N__17971\ : std_logic;
signal \N__17968\ : std_logic;
signal \N__17965\ : std_logic;
signal \N__17962\ : std_logic;
signal \N__17959\ : std_logic;
signal \N__17956\ : std_logic;
signal \N__17955\ : std_logic;
signal \N__17952\ : std_logic;
signal \N__17951\ : std_logic;
signal \N__17948\ : std_logic;
signal \N__17945\ : std_logic;
signal \N__17944\ : std_logic;
signal \N__17941\ : std_logic;
signal \N__17938\ : std_logic;
signal \N__17935\ : std_logic;
signal \N__17932\ : std_logic;
signal \N__17925\ : std_logic;
signal \N__17920\ : std_logic;
signal \N__17917\ : std_logic;
signal \N__17914\ : std_logic;
signal \N__17911\ : std_logic;
signal \N__17908\ : std_logic;
signal \N__17905\ : std_logic;
signal \N__17902\ : std_logic;
signal \N__17899\ : std_logic;
signal \N__17896\ : std_logic;
signal \N__17893\ : std_logic;
signal \N__17890\ : std_logic;
signal \N__17887\ : std_logic;
signal \N__17886\ : std_logic;
signal \N__17885\ : std_logic;
signal \N__17884\ : std_logic;
signal \N__17881\ : std_logic;
signal \N__17878\ : std_logic;
signal \N__17873\ : std_logic;
signal \N__17866\ : std_logic;
signal \N__17863\ : std_logic;
signal \N__17860\ : std_logic;
signal \N__17857\ : std_logic;
signal \N__17854\ : std_logic;
signal \N__17851\ : std_logic;
signal \N__17848\ : std_logic;
signal \N__17845\ : std_logic;
signal \N__17842\ : std_logic;
signal \N__17839\ : std_logic;
signal \N__17838\ : std_logic;
signal \N__17835\ : std_logic;
signal \N__17832\ : std_logic;
signal \N__17829\ : std_logic;
signal \N__17824\ : std_logic;
signal \N__17823\ : std_logic;
signal \N__17822\ : std_logic;
signal \N__17821\ : std_logic;
signal \N__17818\ : std_logic;
signal \N__17815\ : std_logic;
signal \N__17812\ : std_logic;
signal \N__17809\ : std_logic;
signal \N__17804\ : std_logic;
signal \N__17797\ : std_logic;
signal \N__17794\ : std_logic;
signal \N__17791\ : std_logic;
signal \N__17788\ : std_logic;
signal \N__17785\ : std_logic;
signal \N__17782\ : std_logic;
signal \N__17779\ : std_logic;
signal \N__17776\ : std_logic;
signal \N__17773\ : std_logic;
signal \N__17770\ : std_logic;
signal \N__17767\ : std_logic;
signal \N__17764\ : std_logic;
signal \N__17761\ : std_logic;
signal \N__17758\ : std_logic;
signal \N__17757\ : std_logic;
signal \N__17756\ : std_logic;
signal \N__17753\ : std_logic;
signal \N__17750\ : std_logic;
signal \N__17747\ : std_logic;
signal \N__17742\ : std_logic;
signal \N__17741\ : std_logic;
signal \N__17738\ : std_logic;
signal \N__17735\ : std_logic;
signal \N__17732\ : std_logic;
signal \N__17725\ : std_logic;
signal \N__17722\ : std_logic;
signal \N__17719\ : std_logic;
signal \N__17716\ : std_logic;
signal \N__17713\ : std_logic;
signal \N__17712\ : std_logic;
signal \N__17709\ : std_logic;
signal \N__17708\ : std_logic;
signal \N__17705\ : std_logic;
signal \N__17704\ : std_logic;
signal \N__17701\ : std_logic;
signal \N__17698\ : std_logic;
signal \N__17695\ : std_logic;
signal \N__17692\ : std_logic;
signal \N__17683\ : std_logic;
signal \N__17680\ : std_logic;
signal \N__17677\ : std_logic;
signal \N__17674\ : std_logic;
signal \N__17671\ : std_logic;
signal \N__17668\ : std_logic;
signal \N__17665\ : std_logic;
signal \N__17662\ : std_logic;
signal \N__17659\ : std_logic;
signal \N__17656\ : std_logic;
signal \N__17653\ : std_logic;
signal \N__17650\ : std_logic;
signal \N__17647\ : std_logic;
signal \N__17644\ : std_logic;
signal \N__17641\ : std_logic;
signal \N__17638\ : std_logic;
signal \N__17635\ : std_logic;
signal \N__17632\ : std_logic;
signal \N__17629\ : std_logic;
signal \N__17626\ : std_logic;
signal \N__17623\ : std_logic;
signal \N__17620\ : std_logic;
signal \N__17617\ : std_logic;
signal \N__17614\ : std_logic;
signal \N__17611\ : std_logic;
signal \N__17608\ : std_logic;
signal \N__17605\ : std_logic;
signal \N__17602\ : std_logic;
signal \N__17599\ : std_logic;
signal \N__17596\ : std_logic;
signal \N__17593\ : std_logic;
signal \N__17590\ : std_logic;
signal \N__17587\ : std_logic;
signal \N__17584\ : std_logic;
signal \N__17583\ : std_logic;
signal \N__17582\ : std_logic;
signal \N__17579\ : std_logic;
signal \N__17578\ : std_logic;
signal \N__17575\ : std_logic;
signal \N__17572\ : std_logic;
signal \N__17571\ : std_logic;
signal \N__17568\ : std_logic;
signal \N__17565\ : std_logic;
signal \N__17562\ : std_logic;
signal \N__17559\ : std_logic;
signal \N__17556\ : std_logic;
signal \N__17551\ : std_logic;
signal \N__17548\ : std_logic;
signal \N__17541\ : std_logic;
signal \N__17536\ : std_logic;
signal \N__17535\ : std_logic;
signal \N__17532\ : std_logic;
signal \N__17529\ : std_logic;
signal \N__17526\ : std_logic;
signal \N__17521\ : std_logic;
signal \N__17518\ : std_logic;
signal \N__17515\ : std_logic;
signal \N__17512\ : std_logic;
signal \N__17509\ : std_logic;
signal \N__17506\ : std_logic;
signal \N__17503\ : std_logic;
signal \N__17502\ : std_logic;
signal \N__17499\ : std_logic;
signal \N__17498\ : std_logic;
signal \N__17497\ : std_logic;
signal \N__17494\ : std_logic;
signal \N__17491\ : std_logic;
signal \N__17488\ : std_logic;
signal \N__17485\ : std_logic;
signal \N__17476\ : std_logic;
signal \N__17475\ : std_logic;
signal \N__17472\ : std_logic;
signal \N__17471\ : std_logic;
signal \N__17470\ : std_logic;
signal \N__17467\ : std_logic;
signal \N__17464\ : std_logic;
signal \N__17461\ : std_logic;
signal \N__17458\ : std_logic;
signal \N__17449\ : std_logic;
signal \N__17446\ : std_logic;
signal \N__17443\ : std_logic;
signal \N__17442\ : std_logic;
signal \N__17441\ : std_logic;
signal \N__17438\ : std_logic;
signal \N__17437\ : std_logic;
signal \N__17434\ : std_logic;
signal \N__17431\ : std_logic;
signal \N__17426\ : std_logic;
signal \N__17419\ : std_logic;
signal \N__17416\ : std_logic;
signal \N__17413\ : std_logic;
signal \N__17412\ : std_logic;
signal \N__17409\ : std_logic;
signal \N__17408\ : std_logic;
signal \N__17407\ : std_logic;
signal \N__17404\ : std_logic;
signal \N__17401\ : std_logic;
signal \N__17398\ : std_logic;
signal \N__17395\ : std_logic;
signal \N__17386\ : std_logic;
signal \N__17383\ : std_logic;
signal \N__17380\ : std_logic;
signal \N__17377\ : std_logic;
signal \N__17374\ : std_logic;
signal \N__17371\ : std_logic;
signal \N__17370\ : std_logic;
signal \N__17367\ : std_logic;
signal \N__17364\ : std_logic;
signal \N__17359\ : std_logic;
signal \N__17356\ : std_logic;
signal \N__17353\ : std_logic;
signal \N__17350\ : std_logic;
signal \N__17347\ : std_logic;
signal \N__17344\ : std_logic;
signal \N__17343\ : std_logic;
signal \N__17340\ : std_logic;
signal \N__17337\ : std_logic;
signal \N__17332\ : std_logic;
signal \N__17331\ : std_logic;
signal \N__17328\ : std_logic;
signal \N__17325\ : std_logic;
signal \N__17320\ : std_logic;
signal \N__17317\ : std_logic;
signal \N__17314\ : std_logic;
signal \N__17311\ : std_logic;
signal \N__17308\ : std_logic;
signal \N__17305\ : std_logic;
signal \N__17302\ : std_logic;
signal \N__17299\ : std_logic;
signal \N__17296\ : std_logic;
signal \N__17293\ : std_logic;
signal \N__17290\ : std_logic;
signal \N__17287\ : std_logic;
signal \N__17284\ : std_logic;
signal \N__17281\ : std_logic;
signal \N__17278\ : std_logic;
signal \N__17275\ : std_logic;
signal \N__17272\ : std_logic;
signal \N__17269\ : std_logic;
signal \N__17266\ : std_logic;
signal \N__17263\ : std_logic;
signal \N__17260\ : std_logic;
signal \N__17257\ : std_logic;
signal \N__17254\ : std_logic;
signal \N__17251\ : std_logic;
signal \N__17248\ : std_logic;
signal \N__17245\ : std_logic;
signal \N__17242\ : std_logic;
signal \N__17239\ : std_logic;
signal \N__17236\ : std_logic;
signal \N__17233\ : std_logic;
signal \N__17230\ : std_logic;
signal \N__17227\ : std_logic;
signal \N__17224\ : std_logic;
signal \N__17221\ : std_logic;
signal \N__17218\ : std_logic;
signal \N__17215\ : std_logic;
signal \N__17212\ : std_logic;
signal \N__17209\ : std_logic;
signal \N__17206\ : std_logic;
signal \N__17203\ : std_logic;
signal \N__17200\ : std_logic;
signal \N__17197\ : std_logic;
signal \N__17194\ : std_logic;
signal \N__17191\ : std_logic;
signal \N__17188\ : std_logic;
signal \N__17187\ : std_logic;
signal \N__17184\ : std_logic;
signal \N__17181\ : std_logic;
signal \N__17176\ : std_logic;
signal \N__17173\ : std_logic;
signal \N__17172\ : std_logic;
signal \N__17169\ : std_logic;
signal \N__17166\ : std_logic;
signal \N__17161\ : std_logic;
signal \N__17158\ : std_logic;
signal \N__17157\ : std_logic;
signal \N__17154\ : std_logic;
signal \N__17151\ : std_logic;
signal \N__17146\ : std_logic;
signal \N__17143\ : std_logic;
signal \N__17140\ : std_logic;
signal \N__17139\ : std_logic;
signal \N__17136\ : std_logic;
signal \N__17133\ : std_logic;
signal \N__17128\ : std_logic;
signal \N__17125\ : std_logic;
signal \N__17122\ : std_logic;
signal \N__17119\ : std_logic;
signal \N__17118\ : std_logic;
signal \N__17113\ : std_logic;
signal \N__17110\ : std_logic;
signal \N__17107\ : std_logic;
signal \N__17106\ : std_logic;
signal \N__17103\ : std_logic;
signal \N__17100\ : std_logic;
signal \N__17099\ : std_logic;
signal \N__17098\ : std_logic;
signal \N__17097\ : std_logic;
signal \N__17094\ : std_logic;
signal \N__17091\ : std_logic;
signal \N__17084\ : std_logic;
signal \N__17077\ : std_logic;
signal \N__17074\ : std_logic;
signal \N__17073\ : std_logic;
signal \N__17072\ : std_logic;
signal \N__17071\ : std_logic;
signal \N__17068\ : std_logic;
signal \N__17065\ : std_logic;
signal \N__17062\ : std_logic;
signal \N__17057\ : std_logic;
signal \N__17050\ : std_logic;
signal \N__17049\ : std_logic;
signal \N__17048\ : std_logic;
signal \N__17047\ : std_logic;
signal \N__17044\ : std_logic;
signal \N__17041\ : std_logic;
signal \N__17036\ : std_logic;
signal \N__17029\ : std_logic;
signal \N__17028\ : std_logic;
signal \N__17027\ : std_logic;
signal \N__17026\ : std_logic;
signal \N__17023\ : std_logic;
signal \N__17020\ : std_logic;
signal \N__17015\ : std_logic;
signal \N__17008\ : std_logic;
signal \N__17005\ : std_logic;
signal \N__17004\ : std_logic;
signal \N__17001\ : std_logic;
signal \N__16998\ : std_logic;
signal \N__16995\ : std_logic;
signal \N__16992\ : std_logic;
signal \N__16987\ : std_logic;
signal \N__16986\ : std_logic;
signal \N__16983\ : std_logic;
signal \N__16980\ : std_logic;
signal \N__16975\ : std_logic;
signal \N__16974\ : std_logic;
signal \N__16971\ : std_logic;
signal \N__16968\ : std_logic;
signal \N__16965\ : std_logic;
signal \N__16962\ : std_logic;
signal \N__16959\ : std_logic;
signal \N__16956\ : std_logic;
signal \N__16953\ : std_logic;
signal \N__16950\ : std_logic;
signal \N__16947\ : std_logic;
signal \N__16944\ : std_logic;
signal \N__16941\ : std_logic;
signal \N__16938\ : std_logic;
signal \N__16935\ : std_logic;
signal \N__16932\ : std_logic;
signal \N__16929\ : std_logic;
signal \N__16926\ : std_logic;
signal \N__16923\ : std_logic;
signal \N__16920\ : std_logic;
signal \N__16917\ : std_logic;
signal \N__16914\ : std_logic;
signal \N__16911\ : std_logic;
signal \N__16908\ : std_logic;
signal \N__16905\ : std_logic;
signal \N__16902\ : std_logic;
signal \N__16899\ : std_logic;
signal \N__16896\ : std_logic;
signal \N__16893\ : std_logic;
signal \N__16890\ : std_logic;
signal \N__16887\ : std_logic;
signal \N__16884\ : std_logic;
signal \N__16881\ : std_logic;
signal \N__16878\ : std_logic;
signal \N__16875\ : std_logic;
signal \N__16872\ : std_logic;
signal \N__16869\ : std_logic;
signal \N__16866\ : std_logic;
signal \N__16863\ : std_logic;
signal \N__16860\ : std_logic;
signal \N__16857\ : std_logic;
signal \N__16854\ : std_logic;
signal \N__16851\ : std_logic;
signal \N__16848\ : std_logic;
signal \N__16845\ : std_logic;
signal \N__16842\ : std_logic;
signal \N__16839\ : std_logic;
signal \N__16836\ : std_logic;
signal \N__16833\ : std_logic;
signal \N__16830\ : std_logic;
signal \N__16827\ : std_logic;
signal \N__16824\ : std_logic;
signal \N__16821\ : std_logic;
signal \N__16818\ : std_logic;
signal \N__16815\ : std_logic;
signal \N__16812\ : std_logic;
signal \N__16809\ : std_logic;
signal \N__16806\ : std_logic;
signal \N__16803\ : std_logic;
signal \N__16800\ : std_logic;
signal \N__16797\ : std_logic;
signal \N__16794\ : std_logic;
signal \N__16791\ : std_logic;
signal \N__16788\ : std_logic;
signal \N__16785\ : std_logic;
signal \N__16782\ : std_logic;
signal \N__16779\ : std_logic;
signal \N__16776\ : std_logic;
signal \N__16773\ : std_logic;
signal \N__16770\ : std_logic;
signal \N__16765\ : std_logic;
signal \N__16762\ : std_logic;
signal \N__16761\ : std_logic;
signal \N__16760\ : std_logic;
signal \N__16757\ : std_logic;
signal \N__16756\ : std_logic;
signal \N__16755\ : std_logic;
signal \N__16752\ : std_logic;
signal \N__16749\ : std_logic;
signal \N__16746\ : std_logic;
signal \N__16743\ : std_logic;
signal \N__16740\ : std_logic;
signal \N__16729\ : std_logic;
signal \N__16726\ : std_logic;
signal \N__16723\ : std_logic;
signal \N__16720\ : std_logic;
signal \N__16719\ : std_logic;
signal \N__16718\ : std_logic;
signal \N__16717\ : std_logic;
signal \N__16714\ : std_logic;
signal \N__16713\ : std_logic;
signal \N__16712\ : std_logic;
signal \N__16709\ : std_logic;
signal \N__16706\ : std_logic;
signal \N__16705\ : std_logic;
signal \N__16702\ : std_logic;
signal \N__16699\ : std_logic;
signal \N__16694\ : std_logic;
signal \N__16689\ : std_logic;
signal \N__16686\ : std_logic;
signal \N__16683\ : std_logic;
signal \N__16678\ : std_logic;
signal \N__16675\ : std_logic;
signal \N__16668\ : std_logic;
signal \N__16663\ : std_logic;
signal \N__16660\ : std_logic;
signal \N__16657\ : std_logic;
signal \N__16654\ : std_logic;
signal \N__16653\ : std_logic;
signal \N__16650\ : std_logic;
signal \N__16647\ : std_logic;
signal \N__16642\ : std_logic;
signal \N__16639\ : std_logic;
signal \N__16638\ : std_logic;
signal \N__16635\ : std_logic;
signal \N__16632\ : std_logic;
signal \N__16629\ : std_logic;
signal \N__16626\ : std_logic;
signal \N__16623\ : std_logic;
signal \N__16620\ : std_logic;
signal \N__16617\ : std_logic;
signal \N__16614\ : std_logic;
signal \N__16611\ : std_logic;
signal \N__16608\ : std_logic;
signal \N__16605\ : std_logic;
signal \N__16602\ : std_logic;
signal \N__16599\ : std_logic;
signal \N__16596\ : std_logic;
signal \N__16593\ : std_logic;
signal \N__16590\ : std_logic;
signal \N__16587\ : std_logic;
signal \N__16584\ : std_logic;
signal \N__16581\ : std_logic;
signal \N__16578\ : std_logic;
signal \N__16575\ : std_logic;
signal \N__16572\ : std_logic;
signal \N__16569\ : std_logic;
signal \N__16566\ : std_logic;
signal \N__16563\ : std_logic;
signal \N__16560\ : std_logic;
signal \N__16557\ : std_logic;
signal \N__16554\ : std_logic;
signal \N__16551\ : std_logic;
signal \N__16548\ : std_logic;
signal \N__16545\ : std_logic;
signal \N__16542\ : std_logic;
signal \N__16539\ : std_logic;
signal \N__16536\ : std_logic;
signal \N__16533\ : std_logic;
signal \N__16530\ : std_logic;
signal \N__16527\ : std_logic;
signal \N__16524\ : std_logic;
signal \N__16521\ : std_logic;
signal \N__16518\ : std_logic;
signal \N__16515\ : std_logic;
signal \N__16512\ : std_logic;
signal \N__16509\ : std_logic;
signal \N__16506\ : std_logic;
signal \N__16503\ : std_logic;
signal \N__16500\ : std_logic;
signal \N__16497\ : std_logic;
signal \N__16494\ : std_logic;
signal \N__16491\ : std_logic;
signal \N__16488\ : std_logic;
signal \N__16485\ : std_logic;
signal \N__16482\ : std_logic;
signal \N__16479\ : std_logic;
signal \N__16476\ : std_logic;
signal \N__16473\ : std_logic;
signal \N__16470\ : std_logic;
signal \N__16467\ : std_logic;
signal \N__16464\ : std_logic;
signal \N__16461\ : std_logic;
signal \N__16458\ : std_logic;
signal \N__16455\ : std_logic;
signal \N__16452\ : std_logic;
signal \N__16449\ : std_logic;
signal \N__16446\ : std_logic;
signal \N__16443\ : std_logic;
signal \N__16440\ : std_logic;
signal \N__16435\ : std_logic;
signal \N__16432\ : std_logic;
signal \N__16429\ : std_logic;
signal \N__16426\ : std_logic;
signal \N__16423\ : std_logic;
signal \N__16420\ : std_logic;
signal \N__16417\ : std_logic;
signal \N__16414\ : std_logic;
signal \N__16413\ : std_logic;
signal \N__16410\ : std_logic;
signal \N__16407\ : std_logic;
signal \N__16404\ : std_logic;
signal \N__16401\ : std_logic;
signal \N__16398\ : std_logic;
signal \N__16393\ : std_logic;
signal \N__16392\ : std_logic;
signal \N__16389\ : std_logic;
signal \N__16386\ : std_logic;
signal \N__16381\ : std_logic;
signal \N__16378\ : std_logic;
signal \N__16377\ : std_logic;
signal \N__16374\ : std_logic;
signal \N__16371\ : std_logic;
signal \N__16366\ : std_logic;
signal \N__16363\ : std_logic;
signal \N__16360\ : std_logic;
signal \N__16357\ : std_logic;
signal \N__16354\ : std_logic;
signal \N__16351\ : std_logic;
signal \N__16348\ : std_logic;
signal \N__16345\ : std_logic;
signal \N__16342\ : std_logic;
signal \N__16341\ : std_logic;
signal \N__16338\ : std_logic;
signal \N__16335\ : std_logic;
signal \N__16332\ : std_logic;
signal \N__16327\ : std_logic;
signal \N__16324\ : std_logic;
signal \N__16321\ : std_logic;
signal \N__16320\ : std_logic;
signal \N__16317\ : std_logic;
signal \N__16314\ : std_logic;
signal \N__16309\ : std_logic;
signal \N__16308\ : std_logic;
signal \N__16305\ : std_logic;
signal \N__16302\ : std_logic;
signal \N__16299\ : std_logic;
signal \N__16296\ : std_logic;
signal \N__16293\ : std_logic;
signal \N__16290\ : std_logic;
signal \N__16287\ : std_logic;
signal \N__16284\ : std_logic;
signal \N__16281\ : std_logic;
signal \N__16278\ : std_logic;
signal \N__16275\ : std_logic;
signal \N__16272\ : std_logic;
signal \N__16269\ : std_logic;
signal \N__16266\ : std_logic;
signal \N__16263\ : std_logic;
signal \N__16260\ : std_logic;
signal \N__16257\ : std_logic;
signal \N__16254\ : std_logic;
signal \N__16251\ : std_logic;
signal \N__16248\ : std_logic;
signal \N__16245\ : std_logic;
signal \N__16242\ : std_logic;
signal \N__16239\ : std_logic;
signal \N__16236\ : std_logic;
signal \N__16233\ : std_logic;
signal \N__16230\ : std_logic;
signal \N__16227\ : std_logic;
signal \N__16224\ : std_logic;
signal \N__16221\ : std_logic;
signal \N__16218\ : std_logic;
signal \N__16215\ : std_logic;
signal \N__16212\ : std_logic;
signal \N__16209\ : std_logic;
signal \N__16206\ : std_logic;
signal \N__16203\ : std_logic;
signal \N__16200\ : std_logic;
signal \N__16197\ : std_logic;
signal \N__16194\ : std_logic;
signal \N__16191\ : std_logic;
signal \N__16188\ : std_logic;
signal \N__16185\ : std_logic;
signal \N__16182\ : std_logic;
signal \N__16179\ : std_logic;
signal \N__16176\ : std_logic;
signal \N__16173\ : std_logic;
signal \N__16170\ : std_logic;
signal \N__16167\ : std_logic;
signal \N__16164\ : std_logic;
signal \N__16161\ : std_logic;
signal \N__16158\ : std_logic;
signal \N__16155\ : std_logic;
signal \N__16152\ : std_logic;
signal \N__16149\ : std_logic;
signal \N__16146\ : std_logic;
signal \N__16143\ : std_logic;
signal \N__16140\ : std_logic;
signal \N__16137\ : std_logic;
signal \N__16134\ : std_logic;
signal \N__16131\ : std_logic;
signal \N__16128\ : std_logic;
signal \N__16125\ : std_logic;
signal \N__16122\ : std_logic;
signal \N__16119\ : std_logic;
signal \N__16116\ : std_logic;
signal \N__16113\ : std_logic;
signal \N__16110\ : std_logic;
signal \N__16107\ : std_logic;
signal \N__16104\ : std_logic;
signal \N__16101\ : std_logic;
signal \N__16098\ : std_logic;
signal \N__16093\ : std_logic;
signal \N__16090\ : std_logic;
signal \N__16087\ : std_logic;
signal \N__16084\ : std_logic;
signal \N__16081\ : std_logic;
signal \N__16078\ : std_logic;
signal \N__16075\ : std_logic;
signal \N__16072\ : std_logic;
signal \N__16069\ : std_logic;
signal \N__16066\ : std_logic;
signal \N__16063\ : std_logic;
signal \N__16060\ : std_logic;
signal \N__16057\ : std_logic;
signal \N__16054\ : std_logic;
signal \N__16051\ : std_logic;
signal \N__16048\ : std_logic;
signal \N__16045\ : std_logic;
signal \N__16042\ : std_logic;
signal \N__16039\ : std_logic;
signal \N__16038\ : std_logic;
signal \N__16037\ : std_logic;
signal \N__16036\ : std_logic;
signal \N__16033\ : std_logic;
signal \N__16030\ : std_logic;
signal \N__16029\ : std_logic;
signal \N__16026\ : std_logic;
signal \N__16025\ : std_logic;
signal \N__16022\ : std_logic;
signal \N__16019\ : std_logic;
signal \N__16016\ : std_logic;
signal \N__16013\ : std_logic;
signal \N__16010\ : std_logic;
signal \N__16007\ : std_logic;
signal \N__16004\ : std_logic;
signal \N__16001\ : std_logic;
signal \N__15996\ : std_logic;
signal \N__15993\ : std_logic;
signal \N__15990\ : std_logic;
signal \N__15983\ : std_logic;
signal \N__15978\ : std_logic;
signal \N__15973\ : std_logic;
signal \N__15970\ : std_logic;
signal \N__15967\ : std_logic;
signal \N__15964\ : std_logic;
signal \N__15961\ : std_logic;
signal \N__15958\ : std_logic;
signal \N__15955\ : std_logic;
signal \N__15952\ : std_logic;
signal \N__15949\ : std_logic;
signal \N__15948\ : std_logic;
signal \N__15945\ : std_logic;
signal \N__15942\ : std_logic;
signal \N__15939\ : std_logic;
signal \N__15934\ : std_logic;
signal \N__15931\ : std_logic;
signal \N__15930\ : std_logic;
signal \N__15929\ : std_logic;
signal \N__15928\ : std_logic;
signal \N__15927\ : std_logic;
signal \N__15924\ : std_logic;
signal \N__15923\ : std_logic;
signal \N__15922\ : std_logic;
signal \N__15921\ : std_logic;
signal \N__15918\ : std_logic;
signal \N__15915\ : std_logic;
signal \N__15908\ : std_logic;
signal \N__15901\ : std_logic;
signal \N__15892\ : std_logic;
signal \N__15891\ : std_logic;
signal \N__15890\ : std_logic;
signal \N__15889\ : std_logic;
signal \N__15888\ : std_logic;
signal \N__15887\ : std_logic;
signal \N__15886\ : std_logic;
signal \N__15885\ : std_logic;
signal \N__15882\ : std_logic;
signal \N__15879\ : std_logic;
signal \N__15872\ : std_logic;
signal \N__15865\ : std_logic;
signal \N__15856\ : std_logic;
signal \N__15853\ : std_logic;
signal \N__15852\ : std_logic;
signal \N__15849\ : std_logic;
signal \N__15848\ : std_logic;
signal \N__15845\ : std_logic;
signal \N__15844\ : std_logic;
signal \N__15843\ : std_logic;
signal \N__15842\ : std_logic;
signal \N__15839\ : std_logic;
signal \N__15836\ : std_logic;
signal \N__15833\ : std_logic;
signal \N__15830\ : std_logic;
signal \N__15827\ : std_logic;
signal \N__15824\ : std_logic;
signal \N__15821\ : std_logic;
signal \N__15818\ : std_logic;
signal \N__15815\ : std_logic;
signal \N__15808\ : std_logic;
signal \N__15807\ : std_logic;
signal \N__15806\ : std_logic;
signal \N__15803\ : std_logic;
signal \N__15796\ : std_logic;
signal \N__15795\ : std_logic;
signal \N__15792\ : std_logic;
signal \N__15789\ : std_logic;
signal \N__15786\ : std_logic;
signal \N__15783\ : std_logic;
signal \N__15776\ : std_logic;
signal \N__15769\ : std_logic;
signal \N__15766\ : std_logic;
signal \N__15763\ : std_logic;
signal \N__15762\ : std_logic;
signal \N__15761\ : std_logic;
signal \N__15760\ : std_logic;
signal \N__15759\ : std_logic;
signal \N__15758\ : std_logic;
signal \N__15757\ : std_logic;
signal \N__15756\ : std_logic;
signal \N__15755\ : std_logic;
signal \N__15752\ : std_logic;
signal \N__15749\ : std_logic;
signal \N__15746\ : std_logic;
signal \N__15739\ : std_logic;
signal \N__15732\ : std_logic;
signal \N__15721\ : std_logic;
signal \N__15720\ : std_logic;
signal \N__15719\ : std_logic;
signal \N__15716\ : std_logic;
signal \N__15713\ : std_logic;
signal \N__15712\ : std_logic;
signal \N__15709\ : std_logic;
signal \N__15704\ : std_logic;
signal \N__15701\ : std_logic;
signal \N__15698\ : std_logic;
signal \N__15693\ : std_logic;
signal \N__15690\ : std_logic;
signal \N__15687\ : std_logic;
signal \N__15684\ : std_logic;
signal \N__15681\ : std_logic;
signal \N__15678\ : std_logic;
signal \N__15675\ : std_logic;
signal \N__15670\ : std_logic;
signal \N__15667\ : std_logic;
signal \N__15664\ : std_logic;
signal \N__15661\ : std_logic;
signal \N__15658\ : std_logic;
signal \N__15655\ : std_logic;
signal \N__15652\ : std_logic;
signal \N__15649\ : std_logic;
signal \N__15648\ : std_logic;
signal \N__15645\ : std_logic;
signal \N__15642\ : std_logic;
signal \N__15639\ : std_logic;
signal \N__15636\ : std_logic;
signal \N__15633\ : std_logic;
signal \N__15630\ : std_logic;
signal \N__15627\ : std_logic;
signal \N__15624\ : std_logic;
signal \N__15621\ : std_logic;
signal \N__15618\ : std_logic;
signal \N__15615\ : std_logic;
signal \N__15612\ : std_logic;
signal \N__15609\ : std_logic;
signal \N__15606\ : std_logic;
signal \N__15603\ : std_logic;
signal \N__15600\ : std_logic;
signal \N__15597\ : std_logic;
signal \N__15594\ : std_logic;
signal \N__15591\ : std_logic;
signal \N__15588\ : std_logic;
signal \N__15585\ : std_logic;
signal \N__15582\ : std_logic;
signal \N__15579\ : std_logic;
signal \N__15576\ : std_logic;
signal \N__15573\ : std_logic;
signal \N__15570\ : std_logic;
signal \N__15567\ : std_logic;
signal \N__15564\ : std_logic;
signal \N__15561\ : std_logic;
signal \N__15558\ : std_logic;
signal \N__15555\ : std_logic;
signal \N__15552\ : std_logic;
signal \N__15549\ : std_logic;
signal \N__15546\ : std_logic;
signal \N__15543\ : std_logic;
signal \N__15540\ : std_logic;
signal \N__15537\ : std_logic;
signal \N__15534\ : std_logic;
signal \N__15531\ : std_logic;
signal \N__15528\ : std_logic;
signal \N__15525\ : std_logic;
signal \N__15522\ : std_logic;
signal \N__15519\ : std_logic;
signal \N__15516\ : std_logic;
signal \N__15513\ : std_logic;
signal \N__15510\ : std_logic;
signal \N__15507\ : std_logic;
signal \N__15504\ : std_logic;
signal \N__15501\ : std_logic;
signal \N__15498\ : std_logic;
signal \N__15495\ : std_logic;
signal \N__15492\ : std_logic;
signal \N__15489\ : std_logic;
signal \N__15486\ : std_logic;
signal \N__15483\ : std_logic;
signal \N__15480\ : std_logic;
signal \N__15477\ : std_logic;
signal \N__15474\ : std_logic;
signal \N__15471\ : std_logic;
signal \N__15468\ : std_logic;
signal \N__15465\ : std_logic;
signal \N__15462\ : std_logic;
signal \N__15459\ : std_logic;
signal \N__15456\ : std_logic;
signal \N__15453\ : std_logic;
signal \N__15450\ : std_logic;
signal \N__15445\ : std_logic;
signal \N__15442\ : std_logic;
signal \N__15441\ : std_logic;
signal \N__15440\ : std_logic;
signal \N__15435\ : std_logic;
signal \N__15432\ : std_logic;
signal \N__15429\ : std_logic;
signal \N__15426\ : std_logic;
signal \N__15423\ : std_logic;
signal \N__15420\ : std_logic;
signal \N__15417\ : std_logic;
signal \N__15414\ : std_logic;
signal \N__15411\ : std_logic;
signal \N__15408\ : std_logic;
signal \N__15403\ : std_logic;
signal \N__15400\ : std_logic;
signal \N__15397\ : std_logic;
signal \N__15396\ : std_logic;
signal \N__15393\ : std_logic;
signal \N__15390\ : std_logic;
signal \N__15387\ : std_logic;
signal \N__15384\ : std_logic;
signal \N__15381\ : std_logic;
signal \N__15378\ : std_logic;
signal \N__15375\ : std_logic;
signal \N__15372\ : std_logic;
signal \N__15369\ : std_logic;
signal \N__15366\ : std_logic;
signal \N__15363\ : std_logic;
signal \N__15360\ : std_logic;
signal \N__15357\ : std_logic;
signal \N__15354\ : std_logic;
signal \N__15351\ : std_logic;
signal \N__15348\ : std_logic;
signal \N__15345\ : std_logic;
signal \N__15342\ : std_logic;
signal \N__15339\ : std_logic;
signal \N__15336\ : std_logic;
signal \N__15333\ : std_logic;
signal \N__15330\ : std_logic;
signal \N__15327\ : std_logic;
signal \N__15324\ : std_logic;
signal \N__15321\ : std_logic;
signal \N__15318\ : std_logic;
signal \N__15315\ : std_logic;
signal \N__15312\ : std_logic;
signal \N__15309\ : std_logic;
signal \N__15306\ : std_logic;
signal \N__15303\ : std_logic;
signal \N__15300\ : std_logic;
signal \N__15297\ : std_logic;
signal \N__15294\ : std_logic;
signal \N__15291\ : std_logic;
signal \N__15288\ : std_logic;
signal \N__15285\ : std_logic;
signal \N__15282\ : std_logic;
signal \N__15279\ : std_logic;
signal \N__15276\ : std_logic;
signal \N__15273\ : std_logic;
signal \N__15270\ : std_logic;
signal \N__15267\ : std_logic;
signal \N__15264\ : std_logic;
signal \N__15261\ : std_logic;
signal \N__15258\ : std_logic;
signal \N__15255\ : std_logic;
signal \N__15252\ : std_logic;
signal \N__15249\ : std_logic;
signal \N__15246\ : std_logic;
signal \N__15243\ : std_logic;
signal \N__15240\ : std_logic;
signal \N__15237\ : std_logic;
signal \N__15234\ : std_logic;
signal \N__15231\ : std_logic;
signal \N__15228\ : std_logic;
signal \N__15225\ : std_logic;
signal \N__15222\ : std_logic;
signal \N__15219\ : std_logic;
signal \N__15216\ : std_logic;
signal \N__15213\ : std_logic;
signal \N__15210\ : std_logic;
signal \N__15207\ : std_logic;
signal \N__15204\ : std_logic;
signal \N__15201\ : std_logic;
signal \N__15198\ : std_logic;
signal \N__15195\ : std_logic;
signal \N__15192\ : std_logic;
signal \N__15189\ : std_logic;
signal \N__15186\ : std_logic;
signal \N__15185\ : std_logic;
signal \N__15182\ : std_logic;
signal \N__15179\ : std_logic;
signal \N__15176\ : std_logic;
signal \N__15171\ : std_logic;
signal \N__15166\ : std_logic;
signal \N__15163\ : std_logic;
signal \N__15162\ : std_logic;
signal \N__15159\ : std_logic;
signal \N__15156\ : std_logic;
signal \N__15153\ : std_logic;
signal \N__15150\ : std_logic;
signal \N__15147\ : std_logic;
signal \N__15144\ : std_logic;
signal \N__15141\ : std_logic;
signal \N__15138\ : std_logic;
signal \N__15135\ : std_logic;
signal \N__15132\ : std_logic;
signal \N__15129\ : std_logic;
signal \N__15126\ : std_logic;
signal \N__15123\ : std_logic;
signal \N__15120\ : std_logic;
signal \N__15117\ : std_logic;
signal \N__15114\ : std_logic;
signal \N__15111\ : std_logic;
signal \N__15108\ : std_logic;
signal \N__15105\ : std_logic;
signal \N__15102\ : std_logic;
signal \N__15099\ : std_logic;
signal \N__15096\ : std_logic;
signal \N__15093\ : std_logic;
signal \N__15090\ : std_logic;
signal \N__15087\ : std_logic;
signal \N__15084\ : std_logic;
signal \N__15081\ : std_logic;
signal \N__15078\ : std_logic;
signal \N__15075\ : std_logic;
signal \N__15072\ : std_logic;
signal \N__15069\ : std_logic;
signal \N__15066\ : std_logic;
signal \N__15063\ : std_logic;
signal \N__15060\ : std_logic;
signal \N__15057\ : std_logic;
signal \N__15054\ : std_logic;
signal \N__15051\ : std_logic;
signal \N__15048\ : std_logic;
signal \N__15045\ : std_logic;
signal \N__15042\ : std_logic;
signal \N__15039\ : std_logic;
signal \N__15036\ : std_logic;
signal \N__15033\ : std_logic;
signal \N__15030\ : std_logic;
signal \N__15027\ : std_logic;
signal \N__15024\ : std_logic;
signal \N__15021\ : std_logic;
signal \N__15018\ : std_logic;
signal \N__15015\ : std_logic;
signal \N__15012\ : std_logic;
signal \N__15009\ : std_logic;
signal \N__15006\ : std_logic;
signal \N__15003\ : std_logic;
signal \N__15000\ : std_logic;
signal \N__14997\ : std_logic;
signal \N__14994\ : std_logic;
signal \N__14991\ : std_logic;
signal \N__14988\ : std_logic;
signal \N__14985\ : std_logic;
signal \N__14982\ : std_logic;
signal \N__14979\ : std_logic;
signal \N__14976\ : std_logic;
signal \N__14973\ : std_logic;
signal \N__14970\ : std_logic;
signal \N__14967\ : std_logic;
signal \N__14964\ : std_logic;
signal \N__14961\ : std_logic;
signal \N__14958\ : std_logic;
signal \N__14955\ : std_logic;
signal \N__14954\ : std_logic;
signal \N__14951\ : std_logic;
signal \N__14948\ : std_logic;
signal \N__14945\ : std_logic;
signal \N__14942\ : std_logic;
signal \N__14939\ : std_logic;
signal \N__14932\ : std_logic;
signal \N__14929\ : std_logic;
signal \N__14926\ : std_logic;
signal \N__14925\ : std_logic;
signal \N__14922\ : std_logic;
signal \N__14919\ : std_logic;
signal \N__14916\ : std_logic;
signal \N__14913\ : std_logic;
signal \N__14910\ : std_logic;
signal \N__14907\ : std_logic;
signal \N__14904\ : std_logic;
signal \N__14901\ : std_logic;
signal \N__14898\ : std_logic;
signal \N__14895\ : std_logic;
signal \N__14892\ : std_logic;
signal \N__14889\ : std_logic;
signal \N__14886\ : std_logic;
signal \N__14883\ : std_logic;
signal \N__14880\ : std_logic;
signal \N__14877\ : std_logic;
signal \N__14874\ : std_logic;
signal \N__14871\ : std_logic;
signal \N__14868\ : std_logic;
signal \N__14865\ : std_logic;
signal \N__14862\ : std_logic;
signal \N__14859\ : std_logic;
signal \N__14856\ : std_logic;
signal \N__14853\ : std_logic;
signal \N__14850\ : std_logic;
signal \N__14847\ : std_logic;
signal \N__14844\ : std_logic;
signal \N__14841\ : std_logic;
signal \N__14838\ : std_logic;
signal \N__14835\ : std_logic;
signal \N__14832\ : std_logic;
signal \N__14829\ : std_logic;
signal \N__14826\ : std_logic;
signal \N__14823\ : std_logic;
signal \N__14820\ : std_logic;
signal \N__14817\ : std_logic;
signal \N__14814\ : std_logic;
signal \N__14811\ : std_logic;
signal \N__14808\ : std_logic;
signal \N__14805\ : std_logic;
signal \N__14802\ : std_logic;
signal \N__14799\ : std_logic;
signal \N__14796\ : std_logic;
signal \N__14793\ : std_logic;
signal \N__14790\ : std_logic;
signal \N__14787\ : std_logic;
signal \N__14784\ : std_logic;
signal \N__14781\ : std_logic;
signal \N__14778\ : std_logic;
signal \N__14775\ : std_logic;
signal \N__14772\ : std_logic;
signal \N__14769\ : std_logic;
signal \N__14766\ : std_logic;
signal \N__14763\ : std_logic;
signal \N__14760\ : std_logic;
signal \N__14757\ : std_logic;
signal \N__14754\ : std_logic;
signal \N__14751\ : std_logic;
signal \N__14748\ : std_logic;
signal \N__14745\ : std_logic;
signal \N__14742\ : std_logic;
signal \N__14739\ : std_logic;
signal \N__14736\ : std_logic;
signal \N__14733\ : std_logic;
signal \N__14730\ : std_logic;
signal \N__14727\ : std_logic;
signal \N__14724\ : std_logic;
signal \N__14723\ : std_logic;
signal \N__14720\ : std_logic;
signal \N__14717\ : std_logic;
signal \N__14714\ : std_logic;
signal \N__14711\ : std_logic;
signal \N__14708\ : std_logic;
signal \N__14701\ : std_logic;
signal \N__14698\ : std_logic;
signal \N__14695\ : std_logic;
signal \N__14692\ : std_logic;
signal \N__14689\ : std_logic;
signal \N__14686\ : std_logic;
signal \N__14683\ : std_logic;
signal \N__14680\ : std_logic;
signal \N__14677\ : std_logic;
signal \N__14674\ : std_logic;
signal \N__14671\ : std_logic;
signal \N__14668\ : std_logic;
signal \N__14665\ : std_logic;
signal \N__14662\ : std_logic;
signal \N__14659\ : std_logic;
signal \N__14656\ : std_logic;
signal \N__14653\ : std_logic;
signal \N__14650\ : std_logic;
signal \N__14647\ : std_logic;
signal \N__14644\ : std_logic;
signal \N__14641\ : std_logic;
signal \N__14638\ : std_logic;
signal \N__14635\ : std_logic;
signal \N__14632\ : std_logic;
signal \N__14629\ : std_logic;
signal \N__14626\ : std_logic;
signal \N__14623\ : std_logic;
signal \N__14620\ : std_logic;
signal \N__14617\ : std_logic;
signal \N__14614\ : std_logic;
signal \N__14611\ : std_logic;
signal \N__14608\ : std_logic;
signal \N__14605\ : std_logic;
signal \N__14604\ : std_logic;
signal \N__14601\ : std_logic;
signal \N__14598\ : std_logic;
signal \N__14595\ : std_logic;
signal \N__14592\ : std_logic;
signal \N__14587\ : std_logic;
signal \N__14584\ : std_logic;
signal \N__14581\ : std_logic;
signal \N__14578\ : std_logic;
signal \N__14575\ : std_logic;
signal \N__14572\ : std_logic;
signal \N__14569\ : std_logic;
signal \N__14566\ : std_logic;
signal \N__14563\ : std_logic;
signal \N__14560\ : std_logic;
signal \N__14557\ : std_logic;
signal \N__14554\ : std_logic;
signal \N__14551\ : std_logic;
signal \N__14548\ : std_logic;
signal \N__14545\ : std_logic;
signal \N__14542\ : std_logic;
signal \N__14539\ : std_logic;
signal \N__14536\ : std_logic;
signal \N__14533\ : std_logic;
signal \N__14530\ : std_logic;
signal \N__14527\ : std_logic;
signal \N__14524\ : std_logic;
signal \N__14521\ : std_logic;
signal \N__14520\ : std_logic;
signal \N__14517\ : std_logic;
signal \N__14514\ : std_logic;
signal \N__14513\ : std_logic;
signal \N__14508\ : std_logic;
signal \N__14505\ : std_logic;
signal \N__14502\ : std_logic;
signal \N__14499\ : std_logic;
signal \N__14496\ : std_logic;
signal \N__14493\ : std_logic;
signal \N__14490\ : std_logic;
signal \N__14487\ : std_logic;
signal \N__14482\ : std_logic;
signal \N__14479\ : std_logic;
signal \N__14476\ : std_logic;
signal \N__14473\ : std_logic;
signal \N__14470\ : std_logic;
signal \N__14467\ : std_logic;
signal \N__14464\ : std_logic;
signal \N__14463\ : std_logic;
signal \N__14462\ : std_logic;
signal \N__14459\ : std_logic;
signal \N__14456\ : std_logic;
signal \N__14453\ : std_logic;
signal \N__14450\ : std_logic;
signal \N__14447\ : std_logic;
signal \N__14444\ : std_logic;
signal \N__14441\ : std_logic;
signal \N__14438\ : std_logic;
signal \N__14435\ : std_logic;
signal \N__14432\ : std_logic;
signal \N__14429\ : std_logic;
signal \N__14426\ : std_logic;
signal \N__14419\ : std_logic;
signal \N__14416\ : std_logic;
signal \N__14415\ : std_logic;
signal \N__14412\ : std_logic;
signal \N__14411\ : std_logic;
signal \N__14408\ : std_logic;
signal \N__14405\ : std_logic;
signal \N__14402\ : std_logic;
signal \N__14399\ : std_logic;
signal \N__14396\ : std_logic;
signal \N__14393\ : std_logic;
signal \N__14390\ : std_logic;
signal \N__14387\ : std_logic;
signal \N__14384\ : std_logic;
signal \N__14381\ : std_logic;
signal \N__14378\ : std_logic;
signal \N__14375\ : std_logic;
signal \N__14372\ : std_logic;
signal \N__14367\ : std_logic;
signal \N__14364\ : std_logic;
signal \N__14359\ : std_logic;
signal \N__14356\ : std_logic;
signal \N__14353\ : std_logic;
signal \N__14352\ : std_logic;
signal \N__14351\ : std_logic;
signal \N__14348\ : std_logic;
signal \N__14345\ : std_logic;
signal \N__14342\ : std_logic;
signal \N__14339\ : std_logic;
signal \N__14336\ : std_logic;
signal \N__14333\ : std_logic;
signal \N__14330\ : std_logic;
signal \N__14327\ : std_logic;
signal \N__14324\ : std_logic;
signal \N__14321\ : std_logic;
signal \N__14318\ : std_logic;
signal \N__14315\ : std_logic;
signal \N__14310\ : std_logic;
signal \N__14305\ : std_logic;
signal \N__14304\ : std_logic;
signal \N__14301\ : std_logic;
signal \N__14300\ : std_logic;
signal \N__14297\ : std_logic;
signal \N__14294\ : std_logic;
signal \N__14291\ : std_logic;
signal \N__14288\ : std_logic;
signal \N__14285\ : std_logic;
signal \N__14282\ : std_logic;
signal \N__14279\ : std_logic;
signal \N__14276\ : std_logic;
signal \N__14273\ : std_logic;
signal \N__14270\ : std_logic;
signal \N__14267\ : std_logic;
signal \N__14264\ : std_logic;
signal \N__14261\ : std_logic;
signal \N__14254\ : std_logic;
signal \N__14251\ : std_logic;
signal \N__14248\ : std_logic;
signal \N__14245\ : std_logic;
signal \N__14244\ : std_logic;
signal \N__14243\ : std_logic;
signal \N__14240\ : std_logic;
signal \N__14237\ : std_logic;
signal \N__14234\ : std_logic;
signal \N__14231\ : std_logic;
signal \N__14228\ : std_logic;
signal \N__14225\ : std_logic;
signal \N__14222\ : std_logic;
signal \N__14219\ : std_logic;
signal \N__14216\ : std_logic;
signal \N__14213\ : std_logic;
signal \N__14210\ : std_logic;
signal \N__14207\ : std_logic;
signal \N__14204\ : std_logic;
signal \N__14201\ : std_logic;
signal \N__14198\ : std_logic;
signal \N__14193\ : std_logic;
signal \N__14188\ : std_logic;
signal \N__14185\ : std_logic;
signal \N__14182\ : std_logic;
signal \N__14181\ : std_logic;
signal \N__14178\ : std_logic;
signal \N__14175\ : std_logic;
signal \N__14172\ : std_logic;
signal \N__14171\ : std_logic;
signal \N__14168\ : std_logic;
signal \N__14165\ : std_logic;
signal \N__14162\ : std_logic;
signal \N__14159\ : std_logic;
signal \N__14156\ : std_logic;
signal \N__14153\ : std_logic;
signal \N__14150\ : std_logic;
signal \N__14147\ : std_logic;
signal \N__14144\ : std_logic;
signal \N__14141\ : std_logic;
signal \N__14138\ : std_logic;
signal \N__14135\ : std_logic;
signal \N__14132\ : std_logic;
signal \N__14127\ : std_logic;
signal \N__14122\ : std_logic;
signal \N__14121\ : std_logic;
signal \N__14118\ : std_logic;
signal \N__14115\ : std_logic;
signal \N__14110\ : std_logic;
signal \N__14107\ : std_logic;
signal \N__14106\ : std_logic;
signal \N__14103\ : std_logic;
signal \N__14100\ : std_logic;
signal \N__14095\ : std_logic;
signal \N__14094\ : std_logic;
signal \N__14091\ : std_logic;
signal \N__14088\ : std_logic;
signal \N__14085\ : std_logic;
signal \N__14082\ : std_logic;
signal \N__14079\ : std_logic;
signal \N__14076\ : std_logic;
signal \N__14073\ : std_logic;
signal \N__14070\ : std_logic;
signal \N__14067\ : std_logic;
signal \N__14064\ : std_logic;
signal \N__14061\ : std_logic;
signal \N__14058\ : std_logic;
signal \N__14055\ : std_logic;
signal \N__14052\ : std_logic;
signal \N__14049\ : std_logic;
signal \N__14046\ : std_logic;
signal \N__14043\ : std_logic;
signal \N__14040\ : std_logic;
signal \N__14037\ : std_logic;
signal \N__14034\ : std_logic;
signal \N__14031\ : std_logic;
signal \N__14028\ : std_logic;
signal \N__14025\ : std_logic;
signal \N__14022\ : std_logic;
signal \N__14019\ : std_logic;
signal \N__14016\ : std_logic;
signal \N__14013\ : std_logic;
signal \N__14010\ : std_logic;
signal \N__14007\ : std_logic;
signal \N__14004\ : std_logic;
signal \N__14001\ : std_logic;
signal \N__13998\ : std_logic;
signal \N__13995\ : std_logic;
signal \N__13992\ : std_logic;
signal \N__13989\ : std_logic;
signal \N__13986\ : std_logic;
signal \N__13983\ : std_logic;
signal \N__13980\ : std_logic;
signal \N__13977\ : std_logic;
signal \N__13974\ : std_logic;
signal \N__13971\ : std_logic;
signal \N__13968\ : std_logic;
signal \N__13965\ : std_logic;
signal \N__13962\ : std_logic;
signal \N__13959\ : std_logic;
signal \N__13956\ : std_logic;
signal \N__13953\ : std_logic;
signal \N__13950\ : std_logic;
signal \N__13947\ : std_logic;
signal \N__13944\ : std_logic;
signal \N__13941\ : std_logic;
signal \N__13938\ : std_logic;
signal \N__13935\ : std_logic;
signal \N__13932\ : std_logic;
signal \N__13929\ : std_logic;
signal \N__13926\ : std_logic;
signal \N__13923\ : std_logic;
signal \N__13920\ : std_logic;
signal \N__13917\ : std_logic;
signal \N__13914\ : std_logic;
signal \N__13911\ : std_logic;
signal \N__13908\ : std_logic;
signal \N__13905\ : std_logic;
signal \N__13902\ : std_logic;
signal \N__13899\ : std_logic;
signal \N__13896\ : std_logic;
signal \N__13893\ : std_logic;
signal \N__13890\ : std_logic;
signal \N__13887\ : std_logic;
signal \N__13884\ : std_logic;
signal \N__13881\ : std_logic;
signal \N__13876\ : std_logic;
signal \N__13873\ : std_logic;
signal \N__13870\ : std_logic;
signal \N__13867\ : std_logic;
signal \N__13864\ : std_logic;
signal \N__13861\ : std_logic;
signal \N__13858\ : std_logic;
signal \N__13855\ : std_logic;
signal \N__13852\ : std_logic;
signal \N__13849\ : std_logic;
signal \N__13846\ : std_logic;
signal \N__13843\ : std_logic;
signal \N__13840\ : std_logic;
signal \N__13837\ : std_logic;
signal \N__13836\ : std_logic;
signal \N__13835\ : std_logic;
signal \N__13834\ : std_logic;
signal \N__13827\ : std_logic;
signal \N__13824\ : std_logic;
signal \N__13821\ : std_logic;
signal \N__13816\ : std_logic;
signal \N__13813\ : std_logic;
signal \N__13812\ : std_logic;
signal \N__13811\ : std_logic;
signal \N__13808\ : std_logic;
signal \N__13807\ : std_logic;
signal \N__13804\ : std_logic;
signal \N__13797\ : std_logic;
signal \N__13792\ : std_logic;
signal \N__13789\ : std_logic;
signal \N__13786\ : std_logic;
signal \N__13785\ : std_logic;
signal \N__13784\ : std_logic;
signal \N__13783\ : std_logic;
signal \N__13780\ : std_logic;
signal \N__13773\ : std_logic;
signal \N__13768\ : std_logic;
signal \N__13765\ : std_logic;
signal \N__13762\ : std_logic;
signal \N__13761\ : std_logic;
signal \N__13758\ : std_logic;
signal \N__13755\ : std_logic;
signal \N__13754\ : std_logic;
signal \N__13753\ : std_logic;
signal \N__13748\ : std_logic;
signal \N__13745\ : std_logic;
signal \N__13742\ : std_logic;
signal \N__13739\ : std_logic;
signal \N__13736\ : std_logic;
signal \N__13733\ : std_logic;
signal \N__13726\ : std_logic;
signal \N__13723\ : std_logic;
signal \N__13720\ : std_logic;
signal \N__13717\ : std_logic;
signal \N__13714\ : std_logic;
signal \N__13711\ : std_logic;
signal \N__13708\ : std_logic;
signal \N__13705\ : std_logic;
signal \N__13702\ : std_logic;
signal \N__13699\ : std_logic;
signal \N__13696\ : std_logic;
signal \N__13693\ : std_logic;
signal \N__13690\ : std_logic;
signal \N__13687\ : std_logic;
signal \N__13684\ : std_logic;
signal \N__13683\ : std_logic;
signal \N__13682\ : std_logic;
signal \N__13681\ : std_logic;
signal \N__13678\ : std_logic;
signal \N__13673\ : std_logic;
signal \N__13670\ : std_logic;
signal \N__13663\ : std_logic;
signal \N__13660\ : std_logic;
signal \N__13659\ : std_logic;
signal \N__13656\ : std_logic;
signal \N__13655\ : std_logic;
signal \N__13654\ : std_logic;
signal \N__13651\ : std_logic;
signal \N__13646\ : std_logic;
signal \N__13643\ : std_logic;
signal \N__13636\ : std_logic;
signal \N__13633\ : std_logic;
signal \N__13632\ : std_logic;
signal \N__13631\ : std_logic;
signal \N__13630\ : std_logic;
signal \N__13627\ : std_logic;
signal \N__13624\ : std_logic;
signal \N__13621\ : std_logic;
signal \N__13618\ : std_logic;
signal \N__13609\ : std_logic;
signal \N__13606\ : std_logic;
signal \N__13605\ : std_logic;
signal \N__13604\ : std_logic;
signal \N__13603\ : std_logic;
signal \N__13600\ : std_logic;
signal \N__13593\ : std_logic;
signal \N__13588\ : std_logic;
signal \N__13585\ : std_logic;
signal \N__13584\ : std_logic;
signal \N__13583\ : std_logic;
signal \N__13582\ : std_logic;
signal \N__13579\ : std_logic;
signal \N__13574\ : std_logic;
signal \N__13571\ : std_logic;
signal \N__13564\ : std_logic;
signal \N__13561\ : std_logic;
signal \N__13560\ : std_logic;
signal \N__13559\ : std_logic;
signal \N__13558\ : std_logic;
signal \N__13555\ : std_logic;
signal \N__13550\ : std_logic;
signal \N__13547\ : std_logic;
signal \N__13540\ : std_logic;
signal \N__13537\ : std_logic;
signal \N__13536\ : std_logic;
signal \N__13535\ : std_logic;
signal \N__13534\ : std_logic;
signal \N__13529\ : std_logic;
signal \N__13526\ : std_logic;
signal \N__13523\ : std_logic;
signal \N__13516\ : std_logic;
signal \N__13513\ : std_logic;
signal \N__13510\ : std_logic;
signal \N__13509\ : std_logic;
signal \N__13508\ : std_logic;
signal \N__13507\ : std_logic;
signal \N__13504\ : std_logic;
signal \N__13501\ : std_logic;
signal \N__13496\ : std_logic;
signal \N__13489\ : std_logic;
signal \N__13486\ : std_logic;
signal \N__13485\ : std_logic;
signal \N__13482\ : std_logic;
signal \N__13479\ : std_logic;
signal \N__13476\ : std_logic;
signal \N__13475\ : std_logic;
signal \N__13474\ : std_logic;
signal \N__13471\ : std_logic;
signal \N__13468\ : std_logic;
signal \N__13465\ : std_logic;
signal \N__13462\ : std_logic;
signal \N__13455\ : std_logic;
signal \N__13452\ : std_logic;
signal \N__13449\ : std_logic;
signal \N__13446\ : std_logic;
signal \N__13443\ : std_logic;
signal \N__13440\ : std_logic;
signal \N__13435\ : std_logic;
signal \N__13432\ : std_logic;
signal \N__13429\ : std_logic;
signal \N__13426\ : std_logic;
signal \N__13425\ : std_logic;
signal \N__13424\ : std_logic;
signal \N__13419\ : std_logic;
signal \N__13416\ : std_logic;
signal \N__13413\ : std_logic;
signal \N__13408\ : std_logic;
signal \N__13407\ : std_logic;
signal \N__13404\ : std_logic;
signal \N__13401\ : std_logic;
signal \N__13396\ : std_logic;
signal \N__13393\ : std_logic;
signal \N__13390\ : std_logic;
signal \N__13389\ : std_logic;
signal \N__13388\ : std_logic;
signal \N__13381\ : std_logic;
signal \N__13378\ : std_logic;
signal \N__13375\ : std_logic;
signal \N__13374\ : std_logic;
signal \N__13373\ : std_logic;
signal \N__13366\ : std_logic;
signal \N__13363\ : std_logic;
signal \N__13360\ : std_logic;
signal \N__13357\ : std_logic;
signal \N__13356\ : std_logic;
signal \N__13353\ : std_logic;
signal \N__13350\ : std_logic;
signal \N__13345\ : std_logic;
signal \N__13344\ : std_logic;
signal \N__13343\ : std_logic;
signal \N__13342\ : std_logic;
signal \N__13333\ : std_logic;
signal \N__13330\ : std_logic;
signal \N__13327\ : std_logic;
signal \N__13326\ : std_logic;
signal \N__13321\ : std_logic;
signal \N__13318\ : std_logic;
signal \N__13315\ : std_logic;
signal \N__13312\ : std_logic;
signal \N__13309\ : std_logic;
signal \N__13306\ : std_logic;
signal \N__13303\ : std_logic;
signal \N__13300\ : std_logic;
signal \N__13297\ : std_logic;
signal \N__13294\ : std_logic;
signal \N__13291\ : std_logic;
signal \N__13288\ : std_logic;
signal \N__13285\ : std_logic;
signal \N__13282\ : std_logic;
signal \N__13279\ : std_logic;
signal \N__13276\ : std_logic;
signal \N__13273\ : std_logic;
signal \N__13270\ : std_logic;
signal \N__13267\ : std_logic;
signal \N__13264\ : std_logic;
signal \N__13261\ : std_logic;
signal \N__13258\ : std_logic;
signal \N__13255\ : std_logic;
signal \N__13254\ : std_logic;
signal \N__13253\ : std_logic;
signal \N__13250\ : std_logic;
signal \N__13245\ : std_logic;
signal \N__13240\ : std_logic;
signal \N__13237\ : std_logic;
signal \N__13234\ : std_logic;
signal \N__13231\ : std_logic;
signal \N__13228\ : std_logic;
signal \N__13225\ : std_logic;
signal \N__13222\ : std_logic;
signal \N__13221\ : std_logic;
signal \N__13220\ : std_logic;
signal \N__13217\ : std_logic;
signal \N__13212\ : std_logic;
signal \N__13207\ : std_logic;
signal \N__13206\ : std_logic;
signal \N__13203\ : std_logic;
signal \N__13200\ : std_logic;
signal \N__13197\ : std_logic;
signal \N__13194\ : std_logic;
signal \N__13191\ : std_logic;
signal \N__13188\ : std_logic;
signal \N__13185\ : std_logic;
signal \N__13182\ : std_logic;
signal \N__13179\ : std_logic;
signal \N__13176\ : std_logic;
signal \N__13173\ : std_logic;
signal \N__13170\ : std_logic;
signal \N__13167\ : std_logic;
signal \N__13164\ : std_logic;
signal \N__13161\ : std_logic;
signal \N__13158\ : std_logic;
signal \N__13155\ : std_logic;
signal \N__13152\ : std_logic;
signal \N__13149\ : std_logic;
signal \N__13146\ : std_logic;
signal \N__13143\ : std_logic;
signal \N__13140\ : std_logic;
signal \N__13137\ : std_logic;
signal \N__13134\ : std_logic;
signal \N__13131\ : std_logic;
signal \N__13128\ : std_logic;
signal \N__13125\ : std_logic;
signal \N__13122\ : std_logic;
signal \N__13119\ : std_logic;
signal \N__13116\ : std_logic;
signal \N__13113\ : std_logic;
signal \N__13110\ : std_logic;
signal \N__13107\ : std_logic;
signal \N__13104\ : std_logic;
signal \N__13101\ : std_logic;
signal \N__13098\ : std_logic;
signal \N__13095\ : std_logic;
signal \N__13092\ : std_logic;
signal \N__13089\ : std_logic;
signal \N__13086\ : std_logic;
signal \N__13083\ : std_logic;
signal \N__13080\ : std_logic;
signal \N__13077\ : std_logic;
signal \N__13074\ : std_logic;
signal \N__13071\ : std_logic;
signal \N__13068\ : std_logic;
signal \N__13065\ : std_logic;
signal \N__13062\ : std_logic;
signal \N__13059\ : std_logic;
signal \N__13056\ : std_logic;
signal \N__13053\ : std_logic;
signal \N__13050\ : std_logic;
signal \N__13047\ : std_logic;
signal \N__13044\ : std_logic;
signal \N__13041\ : std_logic;
signal \N__13038\ : std_logic;
signal \N__13035\ : std_logic;
signal \N__13032\ : std_logic;
signal \N__13029\ : std_logic;
signal \N__13026\ : std_logic;
signal \N__13023\ : std_logic;
signal \N__13020\ : std_logic;
signal \N__13017\ : std_logic;
signal \N__13014\ : std_logic;
signal \N__13011\ : std_logic;
signal \N__13008\ : std_logic;
signal \N__13005\ : std_logic;
signal \N__13002\ : std_logic;
signal \N__12999\ : std_logic;
signal \N__12996\ : std_logic;
signal \N__12993\ : std_logic;
signal \N__12990\ : std_logic;
signal \N__12987\ : std_logic;
signal \N__12982\ : std_logic;
signal \N__12979\ : std_logic;
signal \N__12976\ : std_logic;
signal \N__12973\ : std_logic;
signal \N__12970\ : std_logic;
signal \N__12967\ : std_logic;
signal \N__12964\ : std_logic;
signal \N__12963\ : std_logic;
signal \N__12960\ : std_logic;
signal \N__12957\ : std_logic;
signal \N__12952\ : std_logic;
signal \N__12949\ : std_logic;
signal \N__12948\ : std_logic;
signal \N__12945\ : std_logic;
signal \N__12942\ : std_logic;
signal \N__12939\ : std_logic;
signal \N__12936\ : std_logic;
signal \N__12933\ : std_logic;
signal \N__12930\ : std_logic;
signal \N__12927\ : std_logic;
signal \N__12924\ : std_logic;
signal \N__12921\ : std_logic;
signal \N__12918\ : std_logic;
signal \N__12915\ : std_logic;
signal \N__12912\ : std_logic;
signal \N__12909\ : std_logic;
signal \N__12906\ : std_logic;
signal \N__12903\ : std_logic;
signal \N__12900\ : std_logic;
signal \N__12897\ : std_logic;
signal \N__12894\ : std_logic;
signal \N__12891\ : std_logic;
signal \N__12888\ : std_logic;
signal \N__12885\ : std_logic;
signal \N__12882\ : std_logic;
signal \N__12879\ : std_logic;
signal \N__12876\ : std_logic;
signal \N__12873\ : std_logic;
signal \N__12870\ : std_logic;
signal \N__12867\ : std_logic;
signal \N__12864\ : std_logic;
signal \N__12861\ : std_logic;
signal \N__12858\ : std_logic;
signal \N__12855\ : std_logic;
signal \N__12852\ : std_logic;
signal \N__12849\ : std_logic;
signal \N__12846\ : std_logic;
signal \N__12843\ : std_logic;
signal \N__12840\ : std_logic;
signal \N__12837\ : std_logic;
signal \N__12834\ : std_logic;
signal \N__12831\ : std_logic;
signal \N__12828\ : std_logic;
signal \N__12825\ : std_logic;
signal \N__12822\ : std_logic;
signal \N__12819\ : std_logic;
signal \N__12816\ : std_logic;
signal \N__12813\ : std_logic;
signal \N__12810\ : std_logic;
signal \N__12807\ : std_logic;
signal \N__12804\ : std_logic;
signal \N__12801\ : std_logic;
signal \N__12798\ : std_logic;
signal \N__12795\ : std_logic;
signal \N__12792\ : std_logic;
signal \N__12789\ : std_logic;
signal \N__12786\ : std_logic;
signal \N__12783\ : std_logic;
signal \N__12780\ : std_logic;
signal \N__12777\ : std_logic;
signal \N__12774\ : std_logic;
signal \N__12771\ : std_logic;
signal \N__12768\ : std_logic;
signal \N__12765\ : std_logic;
signal \N__12762\ : std_logic;
signal \N__12759\ : std_logic;
signal \N__12756\ : std_logic;
signal \N__12753\ : std_logic;
signal \N__12750\ : std_logic;
signal \N__12747\ : std_logic;
signal \N__12744\ : std_logic;
signal \N__12741\ : std_logic;
signal \N__12736\ : std_logic;
signal \N__12733\ : std_logic;
signal \N__12730\ : std_logic;
signal \N__12727\ : std_logic;
signal \N__12724\ : std_logic;
signal \N__12721\ : std_logic;
signal \N__12718\ : std_logic;
signal \N__12715\ : std_logic;
signal \N__12712\ : std_logic;
signal \N__12709\ : std_logic;
signal \N__12706\ : std_logic;
signal \N__12703\ : std_logic;
signal \N__12700\ : std_logic;
signal \N__12697\ : std_logic;
signal \N__12694\ : std_logic;
signal \N__12691\ : std_logic;
signal \N__12688\ : std_logic;
signal \N__12685\ : std_logic;
signal \N__12682\ : std_logic;
signal \N__12679\ : std_logic;
signal \N__12676\ : std_logic;
signal \N__12673\ : std_logic;
signal \N__12670\ : std_logic;
signal \N__12667\ : std_logic;
signal \N__12664\ : std_logic;
signal \N__12661\ : std_logic;
signal \N__12658\ : std_logic;
signal \N__12657\ : std_logic;
signal \N__12656\ : std_logic;
signal \N__12653\ : std_logic;
signal \N__12650\ : std_logic;
signal \N__12647\ : std_logic;
signal \N__12646\ : std_logic;
signal \N__12643\ : std_logic;
signal \N__12638\ : std_logic;
signal \N__12635\ : std_logic;
signal \N__12632\ : std_logic;
signal \N__12627\ : std_logic;
signal \N__12624\ : std_logic;
signal \N__12621\ : std_logic;
signal \N__12618\ : std_logic;
signal \N__12615\ : std_logic;
signal \N__12610\ : std_logic;
signal \N__12607\ : std_logic;
signal \N__12606\ : std_logic;
signal \N__12605\ : std_logic;
signal \N__12602\ : std_logic;
signal \N__12599\ : std_logic;
signal \N__12598\ : std_logic;
signal \N__12595\ : std_logic;
signal \N__12592\ : std_logic;
signal \N__12589\ : std_logic;
signal \N__12586\ : std_logic;
signal \N__12583\ : std_logic;
signal \N__12578\ : std_logic;
signal \N__12575\ : std_logic;
signal \N__12570\ : std_logic;
signal \N__12567\ : std_logic;
signal \N__12562\ : std_logic;
signal \N__12559\ : std_logic;
signal \N__12556\ : std_logic;
signal \N__12553\ : std_logic;
signal \N__12550\ : std_logic;
signal \N__12547\ : std_logic;
signal \N__12546\ : std_logic;
signal \N__12545\ : std_logic;
signal \N__12544\ : std_logic;
signal \N__12543\ : std_logic;
signal \N__12532\ : std_logic;
signal \N__12529\ : std_logic;
signal \N__12526\ : std_logic;
signal \N__12523\ : std_logic;
signal \N__12520\ : std_logic;
signal \N__12517\ : std_logic;
signal \N__12516\ : std_logic;
signal \N__12513\ : std_logic;
signal \N__12512\ : std_logic;
signal \N__12509\ : std_logic;
signal \N__12508\ : std_logic;
signal \N__12507\ : std_logic;
signal \N__12506\ : std_logic;
signal \N__12503\ : std_logic;
signal \N__12500\ : std_logic;
signal \N__12491\ : std_logic;
signal \N__12484\ : std_logic;
signal \N__12481\ : std_logic;
signal \N__12478\ : std_logic;
signal \N__12475\ : std_logic;
signal \N__12472\ : std_logic;
signal \N__12469\ : std_logic;
signal \N__12468\ : std_logic;
signal \N__12465\ : std_logic;
signal \N__12462\ : std_logic;
signal \N__12459\ : std_logic;
signal \N__12456\ : std_logic;
signal \N__12453\ : std_logic;
signal \N__12450\ : std_logic;
signal \N__12447\ : std_logic;
signal \N__12444\ : std_logic;
signal \N__12441\ : std_logic;
signal \N__12438\ : std_logic;
signal \N__12435\ : std_logic;
signal \N__12432\ : std_logic;
signal \N__12429\ : std_logic;
signal \N__12426\ : std_logic;
signal \N__12423\ : std_logic;
signal \N__12420\ : std_logic;
signal \N__12417\ : std_logic;
signal \N__12414\ : std_logic;
signal \N__12411\ : std_logic;
signal \N__12408\ : std_logic;
signal \N__12405\ : std_logic;
signal \N__12402\ : std_logic;
signal \N__12399\ : std_logic;
signal \N__12396\ : std_logic;
signal \N__12393\ : std_logic;
signal \N__12390\ : std_logic;
signal \N__12387\ : std_logic;
signal \N__12384\ : std_logic;
signal \N__12381\ : std_logic;
signal \N__12378\ : std_logic;
signal \N__12375\ : std_logic;
signal \N__12372\ : std_logic;
signal \N__12369\ : std_logic;
signal \N__12366\ : std_logic;
signal \N__12363\ : std_logic;
signal \N__12360\ : std_logic;
signal \N__12357\ : std_logic;
signal \N__12354\ : std_logic;
signal \N__12351\ : std_logic;
signal \N__12348\ : std_logic;
signal \N__12345\ : std_logic;
signal \N__12342\ : std_logic;
signal \N__12339\ : std_logic;
signal \N__12336\ : std_logic;
signal \N__12333\ : std_logic;
signal \N__12330\ : std_logic;
signal \N__12327\ : std_logic;
signal \N__12324\ : std_logic;
signal \N__12321\ : std_logic;
signal \N__12318\ : std_logic;
signal \N__12315\ : std_logic;
signal \N__12312\ : std_logic;
signal \N__12309\ : std_logic;
signal \N__12306\ : std_logic;
signal \N__12303\ : std_logic;
signal \N__12300\ : std_logic;
signal \N__12297\ : std_logic;
signal \N__12294\ : std_logic;
signal \N__12291\ : std_logic;
signal \N__12288\ : std_logic;
signal \N__12285\ : std_logic;
signal \N__12282\ : std_logic;
signal \N__12279\ : std_logic;
signal \N__12276\ : std_logic;
signal \N__12273\ : std_logic;
signal \N__12270\ : std_logic;
signal \N__12267\ : std_logic;
signal \N__12264\ : std_logic;
signal \N__12261\ : std_logic;
signal \N__12258\ : std_logic;
signal \N__12253\ : std_logic;
signal \N__12250\ : std_logic;
signal \N__12247\ : std_logic;
signal \N__12244\ : std_logic;
signal \N__12241\ : std_logic;
signal \N__12238\ : std_logic;
signal \N__12237\ : std_logic;
signal \N__12236\ : std_logic;
signal \N__12235\ : std_logic;
signal \N__12234\ : std_logic;
signal \N__12231\ : std_logic;
signal \N__12222\ : std_logic;
signal \N__12219\ : std_logic;
signal \N__12214\ : std_logic;
signal \N__12213\ : std_logic;
signal \N__12210\ : std_logic;
signal \N__12207\ : std_logic;
signal \N__12204\ : std_logic;
signal \N__12201\ : std_logic;
signal \N__12198\ : std_logic;
signal \N__12195\ : std_logic;
signal \N__12192\ : std_logic;
signal \N__12189\ : std_logic;
signal \N__12186\ : std_logic;
signal \N__12183\ : std_logic;
signal \N__12180\ : std_logic;
signal \N__12177\ : std_logic;
signal \N__12174\ : std_logic;
signal \N__12171\ : std_logic;
signal \N__12168\ : std_logic;
signal \N__12165\ : std_logic;
signal \N__12162\ : std_logic;
signal \N__12159\ : std_logic;
signal \N__12156\ : std_logic;
signal \N__12153\ : std_logic;
signal \N__12150\ : std_logic;
signal \N__12147\ : std_logic;
signal \N__12144\ : std_logic;
signal \N__12141\ : std_logic;
signal \N__12138\ : std_logic;
signal \N__12135\ : std_logic;
signal \N__12132\ : std_logic;
signal \N__12129\ : std_logic;
signal \N__12126\ : std_logic;
signal \N__12123\ : std_logic;
signal \N__12120\ : std_logic;
signal \N__12117\ : std_logic;
signal \N__12114\ : std_logic;
signal \N__12111\ : std_logic;
signal \N__12108\ : std_logic;
signal \N__12105\ : std_logic;
signal \N__12102\ : std_logic;
signal \N__12099\ : std_logic;
signal \N__12096\ : std_logic;
signal \N__12093\ : std_logic;
signal \N__12090\ : std_logic;
signal \N__12087\ : std_logic;
signal \N__12084\ : std_logic;
signal \N__12081\ : std_logic;
signal \N__12078\ : std_logic;
signal \N__12075\ : std_logic;
signal \N__12072\ : std_logic;
signal \N__12069\ : std_logic;
signal \N__12066\ : std_logic;
signal \N__12063\ : std_logic;
signal \N__12060\ : std_logic;
signal \N__12057\ : std_logic;
signal \N__12054\ : std_logic;
signal \N__12051\ : std_logic;
signal \N__12048\ : std_logic;
signal \N__12045\ : std_logic;
signal \N__12042\ : std_logic;
signal \N__12039\ : std_logic;
signal \N__12036\ : std_logic;
signal \N__12033\ : std_logic;
signal \N__12030\ : std_logic;
signal \N__12027\ : std_logic;
signal \N__12024\ : std_logic;
signal \N__12021\ : std_logic;
signal \N__12018\ : std_logic;
signal \N__12015\ : std_logic;
signal \N__12012\ : std_logic;
signal \N__12009\ : std_logic;
signal \N__12006\ : std_logic;
signal \N__12003\ : std_logic;
signal \N__11998\ : std_logic;
signal \N__11995\ : std_logic;
signal \N__11992\ : std_logic;
signal \N__11989\ : std_logic;
signal \N__11988\ : std_logic;
signal \N__11987\ : std_logic;
signal \N__11986\ : std_logic;
signal \N__11983\ : std_logic;
signal \N__11978\ : std_logic;
signal \N__11975\ : std_logic;
signal \N__11968\ : std_logic;
signal \N__11965\ : std_logic;
signal \N__11962\ : std_logic;
signal \N__11959\ : std_logic;
signal \N__11958\ : std_logic;
signal \N__11955\ : std_logic;
signal \N__11952\ : std_logic;
signal \N__11949\ : std_logic;
signal \N__11946\ : std_logic;
signal \N__11943\ : std_logic;
signal \N__11940\ : std_logic;
signal \N__11937\ : std_logic;
signal \N__11934\ : std_logic;
signal \N__11931\ : std_logic;
signal \N__11928\ : std_logic;
signal \N__11925\ : std_logic;
signal \N__11922\ : std_logic;
signal \N__11919\ : std_logic;
signal \N__11916\ : std_logic;
signal \N__11913\ : std_logic;
signal \N__11910\ : std_logic;
signal \N__11907\ : std_logic;
signal \N__11904\ : std_logic;
signal \N__11901\ : std_logic;
signal \N__11898\ : std_logic;
signal \N__11895\ : std_logic;
signal \N__11892\ : std_logic;
signal \N__11889\ : std_logic;
signal \N__11886\ : std_logic;
signal \N__11883\ : std_logic;
signal \N__11880\ : std_logic;
signal \N__11877\ : std_logic;
signal \N__11874\ : std_logic;
signal \N__11871\ : std_logic;
signal \N__11868\ : std_logic;
signal \N__11865\ : std_logic;
signal \N__11862\ : std_logic;
signal \N__11859\ : std_logic;
signal \N__11856\ : std_logic;
signal \N__11853\ : std_logic;
signal \N__11850\ : std_logic;
signal \N__11847\ : std_logic;
signal \N__11844\ : std_logic;
signal \N__11841\ : std_logic;
signal \N__11838\ : std_logic;
signal \N__11835\ : std_logic;
signal \N__11832\ : std_logic;
signal \N__11829\ : std_logic;
signal \N__11826\ : std_logic;
signal \N__11823\ : std_logic;
signal \N__11820\ : std_logic;
signal \N__11817\ : std_logic;
signal \N__11814\ : std_logic;
signal \N__11811\ : std_logic;
signal \N__11808\ : std_logic;
signal \N__11805\ : std_logic;
signal \N__11802\ : std_logic;
signal \N__11799\ : std_logic;
signal \N__11796\ : std_logic;
signal \N__11793\ : std_logic;
signal \N__11790\ : std_logic;
signal \N__11787\ : std_logic;
signal \N__11784\ : std_logic;
signal \N__11781\ : std_logic;
signal \N__11778\ : std_logic;
signal \N__11775\ : std_logic;
signal \N__11772\ : std_logic;
signal \N__11769\ : std_logic;
signal \N__11766\ : std_logic;
signal \N__11763\ : std_logic;
signal \N__11760\ : std_logic;
signal \N__11757\ : std_logic;
signal \N__11754\ : std_logic;
signal \N__11751\ : std_logic;
signal \N__11748\ : std_logic;
signal \N__11745\ : std_logic;
signal \N__11742\ : std_logic;
signal \N__11739\ : std_logic;
signal \N__11734\ : std_logic;
signal \N__11731\ : std_logic;
signal \N__11728\ : std_logic;
signal \N__11725\ : std_logic;
signal \N__11722\ : std_logic;
signal \N__11719\ : std_logic;
signal \N__11716\ : std_logic;
signal \N__11713\ : std_logic;
signal \N__11710\ : std_logic;
signal \N__11709\ : std_logic;
signal \N__11706\ : std_logic;
signal \N__11703\ : std_logic;
signal \N__11700\ : std_logic;
signal \N__11695\ : std_logic;
signal \N__11692\ : std_logic;
signal \N__11691\ : std_logic;
signal \N__11688\ : std_logic;
signal \N__11685\ : std_logic;
signal \N__11682\ : std_logic;
signal \N__11679\ : std_logic;
signal \N__11676\ : std_logic;
signal \N__11673\ : std_logic;
signal \N__11668\ : std_logic;
signal \N__11665\ : std_logic;
signal \N__11662\ : std_logic;
signal \N__11659\ : std_logic;
signal \N__11656\ : std_logic;
signal \N__11655\ : std_logic;
signal \N__11652\ : std_logic;
signal \N__11649\ : std_logic;
signal \N__11646\ : std_logic;
signal \N__11643\ : std_logic;
signal \N__11640\ : std_logic;
signal \N__11637\ : std_logic;
signal \N__11634\ : std_logic;
signal \N__11631\ : std_logic;
signal \N__11628\ : std_logic;
signal \N__11625\ : std_logic;
signal \N__11622\ : std_logic;
signal \N__11619\ : std_logic;
signal \N__11616\ : std_logic;
signal \N__11613\ : std_logic;
signal \N__11610\ : std_logic;
signal \N__11607\ : std_logic;
signal \N__11604\ : std_logic;
signal \N__11601\ : std_logic;
signal \N__11598\ : std_logic;
signal \N__11595\ : std_logic;
signal \N__11592\ : std_logic;
signal \N__11589\ : std_logic;
signal \N__11586\ : std_logic;
signal \N__11583\ : std_logic;
signal \N__11580\ : std_logic;
signal \N__11577\ : std_logic;
signal \N__11574\ : std_logic;
signal \N__11571\ : std_logic;
signal \N__11568\ : std_logic;
signal \N__11565\ : std_logic;
signal \N__11562\ : std_logic;
signal \N__11559\ : std_logic;
signal \N__11556\ : std_logic;
signal \N__11553\ : std_logic;
signal \N__11550\ : std_logic;
signal \N__11547\ : std_logic;
signal \N__11544\ : std_logic;
signal \N__11541\ : std_logic;
signal \N__11538\ : std_logic;
signal \N__11535\ : std_logic;
signal \N__11532\ : std_logic;
signal \N__11529\ : std_logic;
signal \N__11526\ : std_logic;
signal \N__11523\ : std_logic;
signal \N__11520\ : std_logic;
signal \N__11517\ : std_logic;
signal \N__11514\ : std_logic;
signal \N__11511\ : std_logic;
signal \N__11508\ : std_logic;
signal \N__11505\ : std_logic;
signal \N__11502\ : std_logic;
signal \N__11499\ : std_logic;
signal \N__11496\ : std_logic;
signal \N__11493\ : std_logic;
signal \N__11490\ : std_logic;
signal \N__11487\ : std_logic;
signal \N__11484\ : std_logic;
signal \N__11481\ : std_logic;
signal \N__11478\ : std_logic;
signal \N__11475\ : std_logic;
signal \N__11472\ : std_logic;
signal \N__11469\ : std_logic;
signal \N__11466\ : std_logic;
signal \N__11463\ : std_logic;
signal \N__11460\ : std_logic;
signal \N__11457\ : std_logic;
signal \N__11454\ : std_logic;
signal \N__11451\ : std_logic;
signal \N__11448\ : std_logic;
signal \N__11445\ : std_logic;
signal \N__11440\ : std_logic;
signal \N__11437\ : std_logic;
signal \N__11434\ : std_logic;
signal \N__11431\ : std_logic;
signal \N__11428\ : std_logic;
signal \N__11427\ : std_logic;
signal \N__11424\ : std_logic;
signal \N__11421\ : std_logic;
signal \N__11418\ : std_logic;
signal \N__11415\ : std_logic;
signal \N__11412\ : std_logic;
signal \N__11409\ : std_logic;
signal \N__11406\ : std_logic;
signal \N__11403\ : std_logic;
signal \N__11400\ : std_logic;
signal \N__11397\ : std_logic;
signal \N__11394\ : std_logic;
signal \N__11391\ : std_logic;
signal \N__11388\ : std_logic;
signal \N__11385\ : std_logic;
signal \N__11382\ : std_logic;
signal \N__11379\ : std_logic;
signal \N__11376\ : std_logic;
signal \N__11373\ : std_logic;
signal \N__11370\ : std_logic;
signal \N__11367\ : std_logic;
signal \N__11364\ : std_logic;
signal \N__11361\ : std_logic;
signal \N__11358\ : std_logic;
signal \N__11355\ : std_logic;
signal \N__11352\ : std_logic;
signal \N__11349\ : std_logic;
signal \N__11346\ : std_logic;
signal \N__11343\ : std_logic;
signal \N__11340\ : std_logic;
signal \N__11337\ : std_logic;
signal \N__11334\ : std_logic;
signal \N__11331\ : std_logic;
signal \N__11328\ : std_logic;
signal \N__11325\ : std_logic;
signal \N__11322\ : std_logic;
signal \N__11319\ : std_logic;
signal \N__11316\ : std_logic;
signal \N__11313\ : std_logic;
signal \N__11310\ : std_logic;
signal \N__11307\ : std_logic;
signal \N__11304\ : std_logic;
signal \N__11301\ : std_logic;
signal \N__11298\ : std_logic;
signal \N__11295\ : std_logic;
signal \N__11292\ : std_logic;
signal \N__11289\ : std_logic;
signal \N__11286\ : std_logic;
signal \N__11283\ : std_logic;
signal \N__11280\ : std_logic;
signal \N__11277\ : std_logic;
signal \N__11274\ : std_logic;
signal \N__11271\ : std_logic;
signal \N__11268\ : std_logic;
signal \N__11265\ : std_logic;
signal \N__11262\ : std_logic;
signal \N__11259\ : std_logic;
signal \N__11256\ : std_logic;
signal \N__11253\ : std_logic;
signal \N__11250\ : std_logic;
signal \N__11247\ : std_logic;
signal \N__11244\ : std_logic;
signal \N__11241\ : std_logic;
signal \N__11238\ : std_logic;
signal \N__11235\ : std_logic;
signal \N__11232\ : std_logic;
signal \N__11229\ : std_logic;
signal \N__11226\ : std_logic;
signal \N__11223\ : std_logic;
signal \N__11220\ : std_logic;
signal \N__11217\ : std_logic;
signal \N__11212\ : std_logic;
signal \N__11209\ : std_logic;
signal \N__11208\ : std_logic;
signal \N__11205\ : std_logic;
signal \N__11202\ : std_logic;
signal \N__11199\ : std_logic;
signal \N__11196\ : std_logic;
signal \N__11193\ : std_logic;
signal \N__11190\ : std_logic;
signal \N__11187\ : std_logic;
signal \N__11184\ : std_logic;
signal \N__11181\ : std_logic;
signal \N__11178\ : std_logic;
signal \N__11175\ : std_logic;
signal \N__11172\ : std_logic;
signal \N__11169\ : std_logic;
signal \N__11166\ : std_logic;
signal \N__11163\ : std_logic;
signal \N__11160\ : std_logic;
signal \N__11157\ : std_logic;
signal \N__11154\ : std_logic;
signal \N__11151\ : std_logic;
signal \N__11148\ : std_logic;
signal \N__11145\ : std_logic;
signal \N__11142\ : std_logic;
signal \N__11139\ : std_logic;
signal \N__11136\ : std_logic;
signal \N__11133\ : std_logic;
signal \N__11130\ : std_logic;
signal \N__11127\ : std_logic;
signal \N__11124\ : std_logic;
signal \N__11121\ : std_logic;
signal \N__11118\ : std_logic;
signal \N__11115\ : std_logic;
signal \N__11112\ : std_logic;
signal \N__11109\ : std_logic;
signal \N__11106\ : std_logic;
signal \N__11103\ : std_logic;
signal \N__11100\ : std_logic;
signal \N__11097\ : std_logic;
signal \N__11094\ : std_logic;
signal \N__11091\ : std_logic;
signal \N__11088\ : std_logic;
signal \N__11085\ : std_logic;
signal \N__11082\ : std_logic;
signal \N__11079\ : std_logic;
signal \N__11076\ : std_logic;
signal \N__11073\ : std_logic;
signal \N__11070\ : std_logic;
signal \N__11067\ : std_logic;
signal \N__11064\ : std_logic;
signal \N__11061\ : std_logic;
signal \N__11058\ : std_logic;
signal \N__11055\ : std_logic;
signal \N__11052\ : std_logic;
signal \N__11049\ : std_logic;
signal \N__11046\ : std_logic;
signal \N__11043\ : std_logic;
signal \N__11040\ : std_logic;
signal \N__11037\ : std_logic;
signal \N__11034\ : std_logic;
signal \N__11031\ : std_logic;
signal \N__11028\ : std_logic;
signal \N__11025\ : std_logic;
signal \N__11022\ : std_logic;
signal \N__11019\ : std_logic;
signal \N__11016\ : std_logic;
signal \N__11013\ : std_logic;
signal \N__11010\ : std_logic;
signal \N__11007\ : std_logic;
signal \N__11004\ : std_logic;
signal \N__10999\ : std_logic;
signal \N__10996\ : std_logic;
signal \N__10993\ : std_logic;
signal \N__10990\ : std_logic;
signal \N__10987\ : std_logic;
signal \N__10984\ : std_logic;
signal \N__10981\ : std_logic;
signal \N__10978\ : std_logic;
signal \N__10975\ : std_logic;
signal \N__10972\ : std_logic;
signal \N__10969\ : std_logic;
signal \N__10966\ : std_logic;
signal \N__10963\ : std_logic;
signal \N__10960\ : std_logic;
signal \N__10957\ : std_logic;
signal \N__10954\ : std_logic;
signal \N__10951\ : std_logic;
signal \N__10948\ : std_logic;
signal \N__10945\ : std_logic;
signal \N__10942\ : std_logic;
signal \N__10939\ : std_logic;
signal \N__10936\ : std_logic;
signal \N__10933\ : std_logic;
signal \N__10930\ : std_logic;
signal \N__10927\ : std_logic;
signal \N__10924\ : std_logic;
signal \N__10923\ : std_logic;
signal \N__10922\ : std_logic;
signal \N__10919\ : std_logic;
signal \N__10916\ : std_logic;
signal \N__10913\ : std_logic;
signal \N__10910\ : std_logic;
signal \N__10903\ : std_logic;
signal \N__10902\ : std_logic;
signal \N__10901\ : std_logic;
signal \N__10898\ : std_logic;
signal \N__10895\ : std_logic;
signal \N__10892\ : std_logic;
signal \N__10885\ : std_logic;
signal \N__10882\ : std_logic;
signal \N__10879\ : std_logic;
signal \N__10876\ : std_logic;
signal \N__10873\ : std_logic;
signal \N__10870\ : std_logic;
signal \N__10869\ : std_logic;
signal \N__10866\ : std_logic;
signal \N__10863\ : std_logic;
signal \N__10860\ : std_logic;
signal \N__10857\ : std_logic;
signal \N__10854\ : std_logic;
signal \N__10851\ : std_logic;
signal \N__10848\ : std_logic;
signal \N__10845\ : std_logic;
signal \N__10842\ : std_logic;
signal \N__10839\ : std_logic;
signal \N__10836\ : std_logic;
signal \N__10833\ : std_logic;
signal \N__10830\ : std_logic;
signal \N__10827\ : std_logic;
signal \N__10824\ : std_logic;
signal \N__10821\ : std_logic;
signal \N__10818\ : std_logic;
signal \N__10815\ : std_logic;
signal \N__10812\ : std_logic;
signal \N__10809\ : std_logic;
signal \N__10806\ : std_logic;
signal \N__10803\ : std_logic;
signal \N__10800\ : std_logic;
signal \N__10797\ : std_logic;
signal \N__10794\ : std_logic;
signal \N__10791\ : std_logic;
signal \N__10788\ : std_logic;
signal \N__10785\ : std_logic;
signal \N__10782\ : std_logic;
signal \N__10779\ : std_logic;
signal \N__10776\ : std_logic;
signal \N__10773\ : std_logic;
signal \N__10770\ : std_logic;
signal \N__10767\ : std_logic;
signal \N__10764\ : std_logic;
signal \N__10761\ : std_logic;
signal \N__10758\ : std_logic;
signal \N__10755\ : std_logic;
signal \N__10752\ : std_logic;
signal \N__10749\ : std_logic;
signal \N__10746\ : std_logic;
signal \N__10743\ : std_logic;
signal \N__10740\ : std_logic;
signal \N__10737\ : std_logic;
signal \N__10734\ : std_logic;
signal \N__10731\ : std_logic;
signal \N__10728\ : std_logic;
signal \N__10725\ : std_logic;
signal \N__10722\ : std_logic;
signal \N__10719\ : std_logic;
signal \N__10716\ : std_logic;
signal \N__10713\ : std_logic;
signal \N__10710\ : std_logic;
signal \N__10707\ : std_logic;
signal \N__10704\ : std_logic;
signal \N__10701\ : std_logic;
signal \N__10698\ : std_logic;
signal \N__10695\ : std_logic;
signal \N__10692\ : std_logic;
signal \N__10689\ : std_logic;
signal \N__10686\ : std_logic;
signal \N__10683\ : std_logic;
signal \N__10680\ : std_logic;
signal \N__10677\ : std_logic;
signal \N__10674\ : std_logic;
signal \N__10671\ : std_logic;
signal \N__10668\ : std_logic;
signal \N__10665\ : std_logic;
signal \N__10660\ : std_logic;
signal \N__10657\ : std_logic;
signal \N__10654\ : std_logic;
signal \N__10651\ : std_logic;
signal \N__10648\ : std_logic;
signal \N__10645\ : std_logic;
signal \N__10642\ : std_logic;
signal \N__10639\ : std_logic;
signal \N__10636\ : std_logic;
signal \N__10633\ : std_logic;
signal \N__10630\ : std_logic;
signal \N__10627\ : std_logic;
signal \N__10624\ : std_logic;
signal \N__10623\ : std_logic;
signal \N__10620\ : std_logic;
signal \N__10617\ : std_logic;
signal \N__10612\ : std_logic;
signal \N__10609\ : std_logic;
signal \N__10608\ : std_logic;
signal \N__10605\ : std_logic;
signal \N__10602\ : std_logic;
signal \N__10597\ : std_logic;
signal \N__10594\ : std_logic;
signal \N__10591\ : std_logic;
signal \N__10588\ : std_logic;
signal \N__10585\ : std_logic;
signal \N__10584\ : std_logic;
signal \N__10581\ : std_logic;
signal \N__10578\ : std_logic;
signal \N__10575\ : std_logic;
signal \N__10572\ : std_logic;
signal \N__10569\ : std_logic;
signal \N__10566\ : std_logic;
signal \N__10561\ : std_logic;
signal \N__10560\ : std_logic;
signal \N__10559\ : std_logic;
signal \N__10556\ : std_logic;
signal \N__10555\ : std_logic;
signal \N__10552\ : std_logic;
signal \N__10549\ : std_logic;
signal \N__10546\ : std_logic;
signal \N__10543\ : std_logic;
signal \N__10534\ : std_logic;
signal \N__10531\ : std_logic;
signal \N__10528\ : std_logic;
signal \N__10527\ : std_logic;
signal \N__10524\ : std_logic;
signal \N__10521\ : std_logic;
signal \N__10520\ : std_logic;
signal \N__10517\ : std_logic;
signal \N__10516\ : std_logic;
signal \N__10513\ : std_logic;
signal \N__10510\ : std_logic;
signal \N__10507\ : std_logic;
signal \N__10504\ : std_logic;
signal \N__10495\ : std_logic;
signal \N__10494\ : std_logic;
signal \N__10491\ : std_logic;
signal \N__10488\ : std_logic;
signal \N__10483\ : std_logic;
signal \N__10482\ : std_logic;
signal \N__10481\ : std_logic;
signal \N__10478\ : std_logic;
signal \N__10475\ : std_logic;
signal \N__10472\ : std_logic;
signal \N__10465\ : std_logic;
signal \N__10462\ : std_logic;
signal \N__10459\ : std_logic;
signal \N__10456\ : std_logic;
signal \N__10453\ : std_logic;
signal \N__10450\ : std_logic;
signal \N__10447\ : std_logic;
signal \N__10444\ : std_logic;
signal \N__10443\ : std_logic;
signal \N__10440\ : std_logic;
signal \N__10437\ : std_logic;
signal \N__10432\ : std_logic;
signal \N__10429\ : std_logic;
signal \N__10428\ : std_logic;
signal \N__10427\ : std_logic;
signal \N__10424\ : std_logic;
signal \N__10423\ : std_logic;
signal \N__10420\ : std_logic;
signal \N__10417\ : std_logic;
signal \N__10412\ : std_logic;
signal \N__10405\ : std_logic;
signal \N__10402\ : std_logic;
signal \N__10401\ : std_logic;
signal \N__10400\ : std_logic;
signal \N__10399\ : std_logic;
signal \N__10396\ : std_logic;
signal \N__10393\ : std_logic;
signal \N__10388\ : std_logic;
signal \N__10381\ : std_logic;
signal \N__10378\ : std_logic;
signal \N__10375\ : std_logic;
signal \N__10372\ : std_logic;
signal \N__10371\ : std_logic;
signal \N__10370\ : std_logic;
signal \N__10367\ : std_logic;
signal \N__10364\ : std_logic;
signal \N__10361\ : std_logic;
signal \N__10354\ : std_logic;
signal \N__10351\ : std_logic;
signal \N__10350\ : std_logic;
signal \N__10349\ : std_logic;
signal \N__10346\ : std_logic;
signal \N__10341\ : std_logic;
signal \N__10336\ : std_logic;
signal \N__10333\ : std_logic;
signal \N__10330\ : std_logic;
signal \N__10327\ : std_logic;
signal \N__10324\ : std_logic;
signal \N__10321\ : std_logic;
signal \N__10318\ : std_logic;
signal \N__10315\ : std_logic;
signal \N__10312\ : std_logic;
signal \N__10309\ : std_logic;
signal \N__10306\ : std_logic;
signal \N__10303\ : std_logic;
signal \N__10300\ : std_logic;
signal \N__10297\ : std_logic;
signal \N__10294\ : std_logic;
signal \N__10291\ : std_logic;
signal \N__10290\ : std_logic;
signal \N__10285\ : std_logic;
signal \N__10282\ : std_logic;
signal \N__10279\ : std_logic;
signal \N__10276\ : std_logic;
signal \N__10273\ : std_logic;
signal \N__10270\ : std_logic;
signal \N__10269\ : std_logic;
signal \N__10266\ : std_logic;
signal \N__10263\ : std_logic;
signal \N__10262\ : std_logic;
signal \N__10257\ : std_logic;
signal \N__10254\ : std_logic;
signal \N__10253\ : std_logic;
signal \N__10248\ : std_logic;
signal \N__10245\ : std_logic;
signal \N__10240\ : std_logic;
signal \N__10237\ : std_logic;
signal \N__10234\ : std_logic;
signal \N__10231\ : std_logic;
signal \N__10228\ : std_logic;
signal \N__10227\ : std_logic;
signal \N__10226\ : std_logic;
signal \N__10225\ : std_logic;
signal \N__10222\ : std_logic;
signal \N__10219\ : std_logic;
signal \N__10216\ : std_logic;
signal \N__10213\ : std_logic;
signal \N__10206\ : std_logic;
signal \N__10203\ : std_logic;
signal \N__10198\ : std_logic;
signal \N__10195\ : std_logic;
signal \N__10192\ : std_logic;
signal \N__10189\ : std_logic;
signal \N__10188\ : std_logic;
signal \N__10185\ : std_logic;
signal \N__10182\ : std_logic;
signal \N__10181\ : std_logic;
signal \N__10180\ : std_logic;
signal \N__10175\ : std_logic;
signal \N__10172\ : std_logic;
signal \N__10169\ : std_logic;
signal \N__10164\ : std_logic;
signal \N__10161\ : std_logic;
signal \N__10158\ : std_logic;
signal \N__10155\ : std_logic;
signal \N__10152\ : std_logic;
signal \N__10149\ : std_logic;
signal \N__10146\ : std_logic;
signal \N__10143\ : std_logic;
signal \N__10140\ : std_logic;
signal \N__10135\ : std_logic;
signal \N__10132\ : std_logic;
signal \N__10129\ : std_logic;
signal \N__10126\ : std_logic;
signal \N__10123\ : std_logic;
signal \N__10120\ : std_logic;
signal \N__10117\ : std_logic;
signal \N__10114\ : std_logic;
signal \N__10113\ : std_logic;
signal \N__10112\ : std_logic;
signal \N__10109\ : std_logic;
signal \N__10106\ : std_logic;
signal \N__10105\ : std_logic;
signal \N__10102\ : std_logic;
signal \N__10099\ : std_logic;
signal \N__10096\ : std_logic;
signal \N__10093\ : std_logic;
signal \N__10090\ : std_logic;
signal \N__10083\ : std_logic;
signal \N__10078\ : std_logic;
signal \N__10075\ : std_logic;
signal \N__10072\ : std_logic;
signal \N__10069\ : std_logic;
signal \N__10066\ : std_logic;
signal \N__10063\ : std_logic;
signal \N__10060\ : std_logic;
signal \N__10057\ : std_logic;
signal \N__10054\ : std_logic;
signal \N__10051\ : std_logic;
signal \N__10048\ : std_logic;
signal \N__10047\ : std_logic;
signal \N__10044\ : std_logic;
signal \N__10041\ : std_logic;
signal \N__10040\ : std_logic;
signal \N__10037\ : std_logic;
signal \N__10034\ : std_logic;
signal \N__10031\ : std_logic;
signal \N__10026\ : std_logic;
signal \N__10023\ : std_logic;
signal \N__10020\ : std_logic;
signal \N__10017\ : std_logic;
signal \N__10012\ : std_logic;
signal \N__10009\ : std_logic;
signal \N__10006\ : std_logic;
signal \N__10003\ : std_logic;
signal \N__10000\ : std_logic;
signal \N__9997\ : std_logic;
signal \N__9994\ : std_logic;
signal \N__9991\ : std_logic;
signal \N__9988\ : std_logic;
signal \N__9985\ : std_logic;
signal \N__9982\ : std_logic;
signal \N__9979\ : std_logic;
signal \N__9976\ : std_logic;
signal \N__9975\ : std_logic;
signal \N__9972\ : std_logic;
signal \N__9969\ : std_logic;
signal \N__9966\ : std_logic;
signal \N__9963\ : std_logic;
signal \N__9960\ : std_logic;
signal \N__9957\ : std_logic;
signal \N__9954\ : std_logic;
signal \N__9951\ : std_logic;
signal \N__9948\ : std_logic;
signal \N__9945\ : std_logic;
signal \N__9942\ : std_logic;
signal \N__9939\ : std_logic;
signal \N__9936\ : std_logic;
signal \N__9933\ : std_logic;
signal \N__9930\ : std_logic;
signal \N__9927\ : std_logic;
signal \N__9924\ : std_logic;
signal \N__9921\ : std_logic;
signal \N__9918\ : std_logic;
signal \N__9915\ : std_logic;
signal \N__9912\ : std_logic;
signal \N__9909\ : std_logic;
signal \N__9906\ : std_logic;
signal \N__9903\ : std_logic;
signal \N__9900\ : std_logic;
signal \N__9897\ : std_logic;
signal \N__9894\ : std_logic;
signal \N__9891\ : std_logic;
signal \N__9888\ : std_logic;
signal \N__9885\ : std_logic;
signal \N__9882\ : std_logic;
signal \N__9879\ : std_logic;
signal \N__9876\ : std_logic;
signal \N__9873\ : std_logic;
signal \N__9870\ : std_logic;
signal \N__9867\ : std_logic;
signal \N__9864\ : std_logic;
signal \N__9861\ : std_logic;
signal \N__9858\ : std_logic;
signal \N__9855\ : std_logic;
signal \N__9852\ : std_logic;
signal \N__9849\ : std_logic;
signal \N__9846\ : std_logic;
signal \N__9843\ : std_logic;
signal \N__9840\ : std_logic;
signal \N__9837\ : std_logic;
signal \N__9834\ : std_logic;
signal \N__9831\ : std_logic;
signal \N__9828\ : std_logic;
signal \N__9825\ : std_logic;
signal \N__9822\ : std_logic;
signal \N__9819\ : std_logic;
signal \N__9816\ : std_logic;
signal \N__9813\ : std_logic;
signal \N__9810\ : std_logic;
signal \N__9807\ : std_logic;
signal \N__9804\ : std_logic;
signal \N__9801\ : std_logic;
signal \N__9798\ : std_logic;
signal \N__9795\ : std_logic;
signal \N__9792\ : std_logic;
signal \N__9789\ : std_logic;
signal \N__9786\ : std_logic;
signal \N__9783\ : std_logic;
signal \N__9780\ : std_logic;
signal \N__9777\ : std_logic;
signal \N__9772\ : std_logic;
signal \N__9769\ : std_logic;
signal \N__9768\ : std_logic;
signal \N__9765\ : std_logic;
signal \N__9762\ : std_logic;
signal \N__9757\ : std_logic;
signal \N__9754\ : std_logic;
signal \N__9751\ : std_logic;
signal \N__9748\ : std_logic;
signal \N__9745\ : std_logic;
signal \N__9742\ : std_logic;
signal \N__9739\ : std_logic;
signal \N__9736\ : std_logic;
signal \N__9733\ : std_logic;
signal \N__9730\ : std_logic;
signal \N__9727\ : std_logic;
signal \N__9724\ : std_logic;
signal \N__9721\ : std_logic;
signal \N__9718\ : std_logic;
signal \N__9715\ : std_logic;
signal \N__9712\ : std_logic;
signal \N__9709\ : std_logic;
signal \N__9706\ : std_logic;
signal \N__9703\ : std_logic;
signal \N__9700\ : std_logic;
signal \N__9697\ : std_logic;
signal \N__9694\ : std_logic;
signal \N__9691\ : std_logic;
signal \N__9688\ : std_logic;
signal \N__9685\ : std_logic;
signal \N__9682\ : std_logic;
signal \N__9679\ : std_logic;
signal \N__9676\ : std_logic;
signal \N__9673\ : std_logic;
signal \N__9672\ : std_logic;
signal \N__9669\ : std_logic;
signal \N__9666\ : std_logic;
signal \N__9663\ : std_logic;
signal \N__9660\ : std_logic;
signal \N__9657\ : std_logic;
signal \N__9654\ : std_logic;
signal \N__9651\ : std_logic;
signal \N__9648\ : std_logic;
signal \N__9643\ : std_logic;
signal \N__9640\ : std_logic;
signal \N__9637\ : std_logic;
signal \N__9634\ : std_logic;
signal \N__9631\ : std_logic;
signal \N__9628\ : std_logic;
signal \N__9625\ : std_logic;
signal \N__9622\ : std_logic;
signal \N__9621\ : std_logic;
signal \N__9620\ : std_logic;
signal \N__9619\ : std_logic;
signal \N__9616\ : std_logic;
signal \N__9613\ : std_logic;
signal \N__9610\ : std_logic;
signal \N__9607\ : std_logic;
signal \N__9598\ : std_logic;
signal \N__9595\ : std_logic;
signal \N__9594\ : std_logic;
signal \N__9593\ : std_logic;
signal \N__9592\ : std_logic;
signal \N__9589\ : std_logic;
signal \N__9586\ : std_logic;
signal \N__9583\ : std_logic;
signal \N__9580\ : std_logic;
signal \N__9577\ : std_logic;
signal \N__9568\ : std_logic;
signal \N__9565\ : std_logic;
signal \N__9564\ : std_logic;
signal \N__9563\ : std_logic;
signal \N__9562\ : std_logic;
signal \N__9559\ : std_logic;
signal \N__9556\ : std_logic;
signal \N__9553\ : std_logic;
signal \N__9550\ : std_logic;
signal \N__9541\ : std_logic;
signal \N__9538\ : std_logic;
signal \N__9537\ : std_logic;
signal \N__9536\ : std_logic;
signal \N__9535\ : std_logic;
signal \N__9532\ : std_logic;
signal \N__9527\ : std_logic;
signal \N__9524\ : std_logic;
signal \N__9517\ : std_logic;
signal \N__9514\ : std_logic;
signal \N__9513\ : std_logic;
signal \N__9512\ : std_logic;
signal \N__9509\ : std_logic;
signal \N__9506\ : std_logic;
signal \N__9503\ : std_logic;
signal \N__9496\ : std_logic;
signal \N__9493\ : std_logic;
signal \N__9492\ : std_logic;
signal \N__9489\ : std_logic;
signal \N__9488\ : std_logic;
signal \N__9485\ : std_logic;
signal \N__9482\ : std_logic;
signal \N__9479\ : std_logic;
signal \N__9472\ : std_logic;
signal \N__9469\ : std_logic;
signal \N__9468\ : std_logic;
signal \N__9467\ : std_logic;
signal \N__9466\ : std_logic;
signal \N__9463\ : std_logic;
signal \N__9458\ : std_logic;
signal \N__9455\ : std_logic;
signal \N__9448\ : std_logic;
signal \N__9445\ : std_logic;
signal \N__9444\ : std_logic;
signal \N__9443\ : std_logic;
signal \N__9442\ : std_logic;
signal \N__9439\ : std_logic;
signal \N__9436\ : std_logic;
signal \N__9433\ : std_logic;
signal \N__9430\ : std_logic;
signal \N__9421\ : std_logic;
signal \N__9418\ : std_logic;
signal \N__9415\ : std_logic;
signal \N__9412\ : std_logic;
signal \N__9409\ : std_logic;
signal \N__9406\ : std_logic;
signal \N__9403\ : std_logic;
signal \N__9400\ : std_logic;
signal \N__9397\ : std_logic;
signal \N__9394\ : std_logic;
signal \N__9391\ : std_logic;
signal \N__9388\ : std_logic;
signal \N__9385\ : std_logic;
signal \N__9382\ : std_logic;
signal \N__9379\ : std_logic;
signal \N__9376\ : std_logic;
signal \N__9373\ : std_logic;
signal \N__9370\ : std_logic;
signal \N__9367\ : std_logic;
signal \N__9364\ : std_logic;
signal \N__9361\ : std_logic;
signal \N__9358\ : std_logic;
signal \N__9355\ : std_logic;
signal \N__9352\ : std_logic;
signal \N__9349\ : std_logic;
signal \N__9346\ : std_logic;
signal \N__9343\ : std_logic;
signal \N__9340\ : std_logic;
signal \N__9337\ : std_logic;
signal \N__9334\ : std_logic;
signal \N__9331\ : std_logic;
signal \N__9328\ : std_logic;
signal \N__9325\ : std_logic;
signal \N__9322\ : std_logic;
signal \N__9319\ : std_logic;
signal \N__9316\ : std_logic;
signal \N__9313\ : std_logic;
signal \N__9310\ : std_logic;
signal \N__9309\ : std_logic;
signal \N__9308\ : std_logic;
signal \N__9307\ : std_logic;
signal \N__9304\ : std_logic;
signal \N__9301\ : std_logic;
signal \N__9298\ : std_logic;
signal \N__9295\ : std_logic;
signal \N__9286\ : std_logic;
signal \N__9283\ : std_logic;
signal \N__9280\ : std_logic;
signal \N__9277\ : std_logic;
signal \N__9274\ : std_logic;
signal \N__9271\ : std_logic;
signal \N__9268\ : std_logic;
signal \N__9265\ : std_logic;
signal \N__9262\ : std_logic;
signal \N__9259\ : std_logic;
signal \N__9256\ : std_logic;
signal \N__9253\ : std_logic;
signal \N__9250\ : std_logic;
signal \N__9247\ : std_logic;
signal \N__9244\ : std_logic;
signal \N__9241\ : std_logic;
signal \N__9238\ : std_logic;
signal \N__9235\ : std_logic;
signal \N__9232\ : std_logic;
signal \N__9229\ : std_logic;
signal \N__9226\ : std_logic;
signal \N__9223\ : std_logic;
signal \N__9220\ : std_logic;
signal \N__9217\ : std_logic;
signal \N__9214\ : std_logic;
signal \N__9211\ : std_logic;
signal \N__9208\ : std_logic;
signal \N__9205\ : std_logic;
signal \N__9202\ : std_logic;
signal \N__9199\ : std_logic;
signal \N__9196\ : std_logic;
signal \N__9193\ : std_logic;
signal \N__9190\ : std_logic;
signal \N__9187\ : std_logic;
signal \N__9184\ : std_logic;
signal \N__9181\ : std_logic;
signal \N__9178\ : std_logic;
signal \N__9175\ : std_logic;
signal \N__9172\ : std_logic;
signal \N__9169\ : std_logic;
signal \N__9166\ : std_logic;
signal \N__9163\ : std_logic;
signal \N__9160\ : std_logic;
signal \N__9157\ : std_logic;
signal \N__9154\ : std_logic;
signal \N__9151\ : std_logic;
signal \N__9148\ : std_logic;
signal \N__9145\ : std_logic;
signal \N__9142\ : std_logic;
signal \N__9139\ : std_logic;
signal \N__9136\ : std_logic;
signal \N__9133\ : std_logic;
signal \N__9130\ : std_logic;
signal \N__9127\ : std_logic;
signal \N__9124\ : std_logic;
signal \N__9121\ : std_logic;
signal \N__9118\ : std_logic;
signal \N__9115\ : std_logic;
signal \N__9112\ : std_logic;
signal \N__9109\ : std_logic;
signal \N__9106\ : std_logic;
signal \N__9103\ : std_logic;
signal \N__9100\ : std_logic;
signal \N__9097\ : std_logic;
signal \N__9094\ : std_logic;
signal \N__9091\ : std_logic;
signal \N__9088\ : std_logic;
signal \N__9085\ : std_logic;
signal \N__9082\ : std_logic;
signal \N__9079\ : std_logic;
signal \N__9076\ : std_logic;
signal \N__9073\ : std_logic;
signal \N__9070\ : std_logic;
signal \N__9067\ : std_logic;
signal \N__9064\ : std_logic;
signal \N__9061\ : std_logic;
signal \N__9058\ : std_logic;
signal \N__9055\ : std_logic;
signal \N__9052\ : std_logic;
signal \N__9049\ : std_logic;
signal \N__9046\ : std_logic;
signal \N__9043\ : std_logic;
signal \N__9040\ : std_logic;
signal \N__9037\ : std_logic;
signal \N__9034\ : std_logic;
signal \N__9031\ : std_logic;
signal \N__9028\ : std_logic;
signal \N__9025\ : std_logic;
signal \N__9022\ : std_logic;
signal \N__9019\ : std_logic;
signal \N__9016\ : std_logic;
signal \N__9013\ : std_logic;
signal \N__9010\ : std_logic;
signal \N__9009\ : std_logic;
signal \N__9006\ : std_logic;
signal \N__9003\ : std_logic;
signal \N__8998\ : std_logic;
signal \N__8997\ : std_logic;
signal \N__8994\ : std_logic;
signal \N__8991\ : std_logic;
signal \N__8990\ : std_logic;
signal \N__8985\ : std_logic;
signal \N__8982\ : std_logic;
signal \N__8979\ : std_logic;
signal \N__8976\ : std_logic;
signal \N__8975\ : std_logic;
signal \N__8974\ : std_logic;
signal \N__8969\ : std_logic;
signal \N__8966\ : std_logic;
signal \N__8963\ : std_logic;
signal \N__8958\ : std_logic;
signal \N__8955\ : std_logic;
signal \N__8954\ : std_logic;
signal \N__8951\ : std_logic;
signal \N__8948\ : std_logic;
signal \N__8945\ : std_logic;
signal \N__8942\ : std_logic;
signal \N__8941\ : std_logic;
signal \N__8938\ : std_logic;
signal \N__8935\ : std_logic;
signal \N__8932\ : std_logic;
signal \N__8929\ : std_logic;
signal \N__8924\ : std_logic;
signal \N__8919\ : std_logic;
signal \N__8916\ : std_logic;
signal \N__8913\ : std_logic;
signal \N__8910\ : std_logic;
signal \N__8907\ : std_logic;
signal \N__8902\ : std_logic;
signal \N__8899\ : std_logic;
signal \N__8896\ : std_logic;
signal \N__8893\ : std_logic;
signal \N__8890\ : std_logic;
signal \N__8887\ : std_logic;
signal \N__8884\ : std_logic;
signal \N__8883\ : std_logic;
signal \N__8880\ : std_logic;
signal \N__8877\ : std_logic;
signal \N__8876\ : std_logic;
signal \N__8875\ : std_logic;
signal \N__8870\ : std_logic;
signal \N__8867\ : std_logic;
signal \N__8864\ : std_logic;
signal \N__8857\ : std_logic;
signal \N__8856\ : std_logic;
signal \N__8855\ : std_logic;
signal \N__8852\ : std_logic;
signal \N__8849\ : std_logic;
signal \N__8846\ : std_logic;
signal \N__8841\ : std_logic;
signal \N__8840\ : std_logic;
signal \N__8839\ : std_logic;
signal \N__8836\ : std_logic;
signal \N__8833\ : std_logic;
signal \N__8830\ : std_logic;
signal \N__8827\ : std_logic;
signal \N__8824\ : std_logic;
signal \N__8821\ : std_logic;
signal \N__8818\ : std_logic;
signal \N__8815\ : std_logic;
signal \N__8812\ : std_logic;
signal \N__8809\ : std_logic;
signal \N__8806\ : std_logic;
signal \N__8803\ : std_logic;
signal \N__8800\ : std_logic;
signal \N__8797\ : std_logic;
signal \N__8794\ : std_logic;
signal \N__8791\ : std_logic;
signal \N__8788\ : std_logic;
signal \N__8783\ : std_logic;
signal \N__8780\ : std_logic;
signal \N__8773\ : std_logic;
signal \N__8772\ : std_logic;
signal \N__8769\ : std_logic;
signal \N__8766\ : std_logic;
signal \N__8765\ : std_logic;
signal \N__8760\ : std_logic;
signal \N__8757\ : std_logic;
signal \N__8752\ : std_logic;
signal \N__8751\ : std_logic;
signal \N__8750\ : std_logic;
signal \N__8747\ : std_logic;
signal \N__8744\ : std_logic;
signal \N__8743\ : std_logic;
signal \N__8740\ : std_logic;
signal \N__8735\ : std_logic;
signal \N__8732\ : std_logic;
signal \N__8729\ : std_logic;
signal \N__8726\ : std_logic;
signal \N__8723\ : std_logic;
signal \N__8722\ : std_logic;
signal \N__8719\ : std_logic;
signal \N__8716\ : std_logic;
signal \N__8713\ : std_logic;
signal \N__8710\ : std_logic;
signal \N__8707\ : std_logic;
signal \N__8704\ : std_logic;
signal \N__8701\ : std_logic;
signal \N__8698\ : std_logic;
signal \N__8697\ : std_logic;
signal \N__8694\ : std_logic;
signal \N__8691\ : std_logic;
signal \N__8688\ : std_logic;
signal \N__8685\ : std_logic;
signal \N__8682\ : std_logic;
signal \N__8671\ : std_logic;
signal \N__8668\ : std_logic;
signal \N__8667\ : std_logic;
signal \N__8666\ : std_logic;
signal \N__8665\ : std_logic;
signal \N__8662\ : std_logic;
signal \N__8659\ : std_logic;
signal \N__8656\ : std_logic;
signal \N__8653\ : std_logic;
signal \N__8650\ : std_logic;
signal \N__8649\ : std_logic;
signal \N__8646\ : std_logic;
signal \N__8643\ : std_logic;
signal \N__8642\ : std_logic;
signal \N__8639\ : std_logic;
signal \N__8636\ : std_logic;
signal \N__8633\ : std_logic;
signal \N__8630\ : std_logic;
signal \N__8627\ : std_logic;
signal \N__8626\ : std_logic;
signal \N__8625\ : std_logic;
signal \N__8622\ : std_logic;
signal \N__8619\ : std_logic;
signal \N__8616\ : std_logic;
signal \N__8613\ : std_logic;
signal \N__8610\ : std_logic;
signal \N__8607\ : std_logic;
signal \N__8604\ : std_logic;
signal \N__8601\ : std_logic;
signal \N__8598\ : std_logic;
signal \N__8595\ : std_logic;
signal \N__8588\ : std_logic;
signal \N__8583\ : std_logic;
signal \N__8580\ : std_logic;
signal \N__8577\ : std_logic;
signal \N__8574\ : std_logic;
signal \N__8567\ : std_logic;
signal \N__8564\ : std_logic;
signal \N__8557\ : std_logic;
signal \N__8556\ : std_logic;
signal \N__8553\ : std_logic;
signal \N__8550\ : std_logic;
signal \N__8547\ : std_logic;
signal \N__8546\ : std_logic;
signal \N__8543\ : std_logic;
signal \N__8540\ : std_logic;
signal \N__8537\ : std_logic;
signal \N__8536\ : std_logic;
signal \N__8533\ : std_logic;
signal \N__8528\ : std_logic;
signal \N__8525\ : std_logic;
signal \N__8522\ : std_logic;
signal \N__8521\ : std_logic;
signal \N__8516\ : std_logic;
signal \N__8515\ : std_logic;
signal \N__8512\ : std_logic;
signal \N__8509\ : std_logic;
signal \N__8508\ : std_logic;
signal \N__8505\ : std_logic;
signal \N__8502\ : std_logic;
signal \N__8497\ : std_logic;
signal \N__8494\ : std_logic;
signal \N__8489\ : std_logic;
signal \N__8484\ : std_logic;
signal \N__8483\ : std_logic;
signal \N__8480\ : std_logic;
signal \N__8477\ : std_logic;
signal \N__8474\ : std_logic;
signal \N__8471\ : std_logic;
signal \N__8466\ : std_logic;
signal \N__8463\ : std_logic;
signal \N__8460\ : std_logic;
signal \N__8455\ : std_logic;
signal \N__8452\ : std_logic;
signal \N__8451\ : std_logic;
signal \N__8448\ : std_logic;
signal \N__8447\ : std_logic;
signal \N__8444\ : std_logic;
signal \N__8441\ : std_logic;
signal \N__8440\ : std_logic;
signal \N__8437\ : std_logic;
signal \N__8434\ : std_logic;
signal \N__8433\ : std_logic;
signal \N__8430\ : std_logic;
signal \N__8427\ : std_logic;
signal \N__8424\ : std_logic;
signal \N__8421\ : std_logic;
signal \N__8418\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8412\ : std_logic;
signal \N__8411\ : std_logic;
signal \N__8408\ : std_logic;
signal \N__8403\ : std_logic;
signal \N__8400\ : std_logic;
signal \N__8397\ : std_logic;
signal \N__8394\ : std_logic;
signal \N__8391\ : std_logic;
signal \N__8386\ : std_logic;
signal \N__8381\ : std_logic;
signal \N__8380\ : std_logic;
signal \N__8377\ : std_logic;
signal \N__8374\ : std_logic;
signal \N__8371\ : std_logic;
signal \N__8368\ : std_logic;
signal \N__8363\ : std_logic;
signal \N__8358\ : std_logic;
signal \N__8355\ : std_logic;
signal \N__8352\ : std_logic;
signal \N__8347\ : std_logic;
signal \N__8346\ : std_logic;
signal \N__8343\ : std_logic;
signal \N__8340\ : std_logic;
signal \N__8337\ : std_logic;
signal \N__8336\ : std_logic;
signal \N__8335\ : std_logic;
signal \N__8332\ : std_logic;
signal \N__8329\ : std_logic;
signal \N__8326\ : std_logic;
signal \N__8325\ : std_logic;
signal \N__8322\ : std_logic;
signal \N__8321\ : std_logic;
signal \N__8318\ : std_logic;
signal \N__8313\ : std_logic;
signal \N__8310\ : std_logic;
signal \N__8307\ : std_logic;
signal \N__8304\ : std_logic;
signal \N__8301\ : std_logic;
signal \N__8296\ : std_logic;
signal \N__8293\ : std_logic;
signal \N__8290\ : std_logic;
signal \N__8289\ : std_logic;
signal \N__8286\ : std_logic;
signal \N__8283\ : std_logic;
signal \N__8280\ : std_logic;
signal \N__8277\ : std_logic;
signal \N__8274\ : std_logic;
signal \N__8271\ : std_logic;
signal \N__8268\ : std_logic;
signal \N__8265\ : std_logic;
signal \N__8262\ : std_logic;
signal \N__8259\ : std_logic;
signal \N__8258\ : std_logic;
signal \N__8255\ : std_logic;
signal \N__8252\ : std_logic;
signal \N__8245\ : std_logic;
signal \N__8242\ : std_logic;
signal \N__8237\ : std_logic;
signal \N__8234\ : std_logic;
signal \N__8231\ : std_logic;
signal \N__8228\ : std_logic;
signal \N__8225\ : std_logic;
signal \N__8222\ : std_logic;
signal \N__8215\ : std_logic;
signal \N__8214\ : std_logic;
signal \N__8211\ : std_logic;
signal \N__8208\ : std_logic;
signal \N__8207\ : std_logic;
signal \N__8206\ : std_logic;
signal \N__8203\ : std_logic;
signal \N__8200\ : std_logic;
signal \N__8197\ : std_logic;
signal \N__8194\ : std_logic;
signal \N__8193\ : std_logic;
signal \N__8190\ : std_logic;
signal \N__8187\ : std_logic;
signal \N__8184\ : std_logic;
signal \N__8183\ : std_logic;
signal \N__8182\ : std_logic;
signal \N__8179\ : std_logic;
signal \N__8176\ : std_logic;
signal \N__8175\ : std_logic;
signal \N__8172\ : std_logic;
signal \N__8169\ : std_logic;
signal \N__8166\ : std_logic;
signal \N__8163\ : std_logic;
signal \N__8160\ : std_logic;
signal \N__8157\ : std_logic;
signal \N__8154\ : std_logic;
signal \N__8151\ : std_logic;
signal \N__8146\ : std_logic;
signal \N__8143\ : std_logic;
signal \N__8140\ : std_logic;
signal \N__8137\ : std_logic;
signal \N__8130\ : std_logic;
signal \N__8125\ : std_logic;
signal \N__8122\ : std_logic;
signal \N__8119\ : std_logic;
signal \N__8116\ : std_logic;
signal \N__8109\ : std_logic;
signal \TVP_VIDEO_c_3\ : std_logic;
signal \VCCG0\ : std_logic;
signal \TVP_VIDEO_c_5\ : std_logic;
signal \TVP_VIDEO_c_4\ : std_logic;
signal \GNDG0\ : std_logic;
signal \TVP_VIDEO_c_7\ : std_logic;
signal \TVP_VIDEO_c_6\ : std_logic;
signal \TVP_VIDEO_c_8\ : std_logic;
signal \TVP_VIDEO_c_9\ : std_logic;
signal \TVP_VIDEO_c_2\ : std_logic;
signal \receive_module.rx_counter.n12_cascade_\ : std_logic;
signal \receive_module.rx_counter.n3938_cascade_\ : std_logic;
signal \receive_module.rx_counter.n3938\ : std_logic;
signal \receive_module.rx_counter.n13\ : std_logic;
signal \receive_module.rx_counter.n3176_cascade_\ : std_logic;
signal \receive_module.rx_counter.n3208\ : std_logic;
signal \line_buffer.n675\ : std_logic;
signal \line_buffer.n683\ : std_logic;
signal \line_buffer.n611\ : std_logic;
signal \line_buffer.n4170_cascade_\ : std_logic;
signal \line_buffer.n619\ : std_logic;
signal \line_buffer.n643\ : std_logic;
signal \line_buffer.n651\ : std_logic;
signal \line_buffer.n687\ : std_logic;
signal \line_buffer.n679\ : std_logic;
signal \line_buffer.n4152\ : std_logic;
signal \line_buffer.n554\ : std_logic;
signal \line_buffer.n546\ : std_logic;
signal \line_buffer.n4155_cascade_\ : std_logic;
signal \line_buffer.n4173\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_95\ : std_logic;
signal \line_buffer.n680\ : std_logic;
signal \line_buffer.n688\ : std_logic;
signal \bfn_10_9_0_\ : std_logic;
signal \receive_module.rx_counter.n3669\ : std_logic;
signal \receive_module.rx_counter.n3670\ : std_logic;
signal \receive_module.rx_counter.n3671\ : std_logic;
signal \receive_module.rx_counter.n3672\ : std_logic;
signal \receive_module.rx_counter.n3673\ : std_logic;
signal \receive_module.rx_counter.n3674\ : std_logic;
signal \receive_module.rx_counter.n3675\ : std_logic;
signal \receive_module.rx_counter.n3676\ : std_logic;
signal \bfn_10_10_0_\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_84\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_83\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_90\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_89\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_88\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_87\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_92\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_91\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_86\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_85\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_94\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_93\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_96\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_97\ : std_logic;
signal \line_buffer.n624\ : std_logic;
signal \line_buffer.n4122\ : std_logic;
signal \line_buffer.n616\ : std_logic;
signal \receive_module.rx_counter.Y_0\ : std_logic;
signal \bfn_11_9_0_\ : std_logic;
signal \receive_module.rx_counter.Y_1\ : std_logic;
signal \receive_module.rx_counter.n3711\ : std_logic;
signal \receive_module.rx_counter.Y_2\ : std_logic;
signal \receive_module.rx_counter.n3712\ : std_logic;
signal \receive_module.rx_counter.Y_3\ : std_logic;
signal \receive_module.rx_counter.n3713\ : std_logic;
signal \receive_module.rx_counter.Y_4\ : std_logic;
signal \receive_module.rx_counter.n3714\ : std_logic;
signal \receive_module.rx_counter.Y_5\ : std_logic;
signal \receive_module.rx_counter.n3715\ : std_logic;
signal \receive_module.rx_counter.Y_6\ : std_logic;
signal \receive_module.rx_counter.n3716\ : std_logic;
signal \receive_module.rx_counter.Y_7\ : std_logic;
signal \receive_module.rx_counter.n3717\ : std_logic;
signal \receive_module.rx_counter.n3718\ : std_logic;
signal \receive_module.rx_counter.Y_8\ : std_logic;
signal \bfn_11_10_0_\ : std_logic;
signal \receive_module.rx_counter.n3979\ : std_logic;
signal \receive_module.rx_counter.O_VISIBLE_N_89\ : std_logic;
signal \DEBUG_c_6\ : std_logic;
signal \transmit_module.video_signal_controller.SYNC_BUFF1\ : std_logic;
signal \transmit_module.video_signal_controller.n3987_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.n4_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.n3935\ : std_logic;
signal \transmit_module.video_signal_controller.n3935_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.n6\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_98\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_76\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_73\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_82\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_75\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_74\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_77\ : std_logic;
signal n1996 : std_logic;
signal \INVADV_R__i1C_net\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_70\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_72\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_71\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_63\ : std_logic;
signal n18 : std_logic;
signal \receive_module.rx_counter.PULSE_1HZ_N_97\ : std_logic;
signal \receive_module.n4212_cascade_\ : std_logic;
signal \receive_module.n4213_cascade_\ : std_logic;
signal \receive_module.rx_counter.n3204\ : std_logic;
signal n659 : std_logic;
signal \DEBUG_c_0\ : std_logic;
signal n691 : std_logic;
signal \line_buffer.n626\ : std_logic;
signal \line_buffer.n561\ : std_logic;
signal \transmit_module.video_signal_controller.n3978_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.n4052\ : std_logic;
signal \transmit_module.video_signal_controller.n4216_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.n12\ : std_logic;
signal \transmit_module.video_signal_controller.n2274_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.SYNC_BUFF2\ : std_logic;
signal \transmit_module.video_signal_controller.n3226\ : std_logic;
signal \transmit_module.video_signal_controller.n2260\ : std_logic;
signal \transmit_module.video_signal_controller.n3917\ : std_logic;
signal \transmit_module.video_signal_controller.n2260_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.n4217\ : std_logic;
signal \transmit_module.video_signal_controller.n18_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.n2219\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_0\ : std_logic;
signal \bfn_12_16_0_\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_1\ : std_logic;
signal \transmit_module.video_signal_controller.n3677\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_2\ : std_logic;
signal \transmit_module.video_signal_controller.n3678\ : std_logic;
signal \transmit_module.video_signal_controller.n3679\ : std_logic;
signal \transmit_module.video_signal_controller.n3680\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_5\ : std_logic;
signal \transmit_module.video_signal_controller.n3681\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_6\ : std_logic;
signal \transmit_module.video_signal_controller.n3682\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_7\ : std_logic;
signal \transmit_module.video_signal_controller.n3683\ : std_logic;
signal \transmit_module.video_signal_controller.n3684\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_8\ : std_logic;
signal \bfn_12_17_0_\ : std_logic;
signal \transmit_module.video_signal_controller.n3685\ : std_logic;
signal \transmit_module.video_signal_controller.n3686\ : std_logic;
signal \transmit_module.video_signal_controller.n3687\ : std_logic;
signal \transmit_module.video_signal_controller.n2594\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_3\ : std_logic;
signal \transmit_module.video_signal_controller.n4215\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_4\ : std_logic;
signal \transmit_module.video_signal_controller.n3892\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_9\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_VISIBLE_Y_N_553_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.n3936\ : std_logic;
signal \transmit_module.n3926_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_11\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_10\ : std_logic;
signal \transmit_module.video_signal_controller.n4218\ : std_logic;
signal \transmit_module.n219_cascade_\ : std_logic;
signal n28 : std_logic;
signal n4210 : std_logic;
signal \n4210_cascade_\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_64\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_67\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_81\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_69\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_68\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_78\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_62\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_66\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_65\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_80\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_79\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_57\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_10\ : std_logic;
signal \transmit_module.n209\ : std_logic;
signal \transmit_module.n178\ : std_logic;
signal \transmit_module.n209_cascade_\ : std_logic;
signal n2283 : std_logic;
signal \old_HS\ : std_logic;
signal \RX_ADDR_3\ : std_logic;
signal \bfn_13_10_0_\ : std_logic;
signal \RX_ADDR_4\ : std_logic;
signal \receive_module.rx_counter.n3650\ : std_logic;
signal \RX_ADDR_5\ : std_logic;
signal \receive_module.rx_counter.n3651\ : std_logic;
signal \receive_module.rx_counter.n3652\ : std_logic;
signal \receive_module.rx_counter.n3653\ : std_logic;
signal \receive_module.rx_counter.n3654\ : std_logic;
signal \receive_module.rx_counter.n3655\ : std_logic;
signal \receive_module.O_X_9\ : std_logic;
signal \receive_module.rx_counter.n4\ : std_logic;
signal \receive_module.O_Y_0\ : std_logic;
signal \receive_module.O_X_6\ : std_logic;
signal \RX_ADDR_6\ : std_logic;
signal \bfn_13_11_0_\ : std_logic;
signal \receive_module.O_X_7\ : std_logic;
signal \receive_module.O_Y_1\ : std_logic;
signal \RX_ADDR_7\ : std_logic;
signal \receive_module.n3699\ : std_logic;
signal \receive_module.O_Y_2\ : std_logic;
signal \receive_module.O_X_8\ : std_logic;
signal \RX_ADDR_8\ : std_logic;
signal \receive_module.n3700\ : std_logic;
signal \receive_module.n7\ : std_logic;
signal \receive_module.O_Y_3\ : std_logic;
signal \RX_ADDR_9\ : std_logic;
signal \receive_module.n3701\ : std_logic;
signal \receive_module.n6\ : std_logic;
signal \receive_module.O_Y_4\ : std_logic;
signal \RX_ADDR_10\ : std_logic;
signal \receive_module.n3702\ : std_logic;
signal \receive_module.n5\ : std_logic;
signal \receive_module.O_Y_5\ : std_logic;
signal \receive_module.n3703\ : std_logic;
signal \receive_module.n4\ : std_logic;
signal \receive_module.O_Y_6\ : std_logic;
signal \receive_module.n3704\ : std_logic;
signal \receive_module.n3\ : std_logic;
signal \receive_module.O_Y_7\ : std_logic;
signal \receive_module.n3705\ : std_logic;
signal \line_buffer.n627\ : std_logic;
signal \line_buffer.n562\ : std_logic;
signal n690 : std_logic;
signal \db5.COUNTER_3\ : std_logic;
signal \db5.NEXT_COUNTER_3\ : std_logic;
signal \db5.COUNTER_2\ : std_logic;
signal \db5.NEXT_COUNTER_2\ : std_logic;
signal \db5.COUNTER_1\ : std_logic;
signal \db5.NEXT_COUNTER_1\ : std_logic;
signal \db5.COUNTER_0\ : std_logic;
signal \db5.NEXT_COUNTER_0\ : std_logic;
signal \INVdb5.NEXT_COUNTER__i3C_net\ : std_logic;
signal \db5.n4221\ : std_logic;
signal \transmit_module.video_signal_controller.n3997\ : std_logic;
signal \transmit_module.video_signal_controller.n3196\ : std_logic;
signal \line_buffer.n655\ : std_logic;
signal \line_buffer.n647\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_0\ : std_logic;
signal \bfn_13_15_0_\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_1\ : std_logic;
signal \transmit_module.video_signal_controller.n3688\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_2\ : std_logic;
signal \transmit_module.video_signal_controller.n3689\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_3\ : std_logic;
signal \transmit_module.video_signal_controller.n3690\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_4\ : std_logic;
signal \transmit_module.video_signal_controller.n3691\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_5\ : std_logic;
signal \transmit_module.video_signal_controller.n3692\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_6\ : std_logic;
signal \transmit_module.video_signal_controller.n3693\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_7\ : std_logic;
signal \transmit_module.video_signal_controller.n3694\ : std_logic;
signal \transmit_module.video_signal_controller.n3695\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_8\ : std_logic;
signal \bfn_13_16_0_\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_9\ : std_logic;
signal \transmit_module.video_signal_controller.n3696\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_10\ : std_logic;
signal \transmit_module.video_signal_controller.n3697\ : std_logic;
signal \transmit_module.video_signal_controller.n3698\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_11\ : std_logic;
signal \transmit_module.video_signal_controller.n2274\ : std_logic;
signal \line_buffer.n4102\ : std_logic;
signal \line_buffer.n648\ : std_logic;
signal \line_buffer.n656\ : std_logic;
signal \transmit_module.n186\ : std_logic;
signal \transmit_module.n4211_cascade_\ : std_logic;
signal \transmit_module.n217\ : std_logic;
signal n26 : std_logic;
signal \line_buffer.n559\ : std_logic;
signal \line_buffer.n4182\ : std_logic;
signal \line_buffer.n551\ : std_logic;
signal \line_buffer.n4185_cascade_\ : std_logic;
signal \line_buffer.n4125\ : std_logic;
signal n1995 : std_logic;
signal \TX_DATA_2\ : std_logic;
signal n1994 : std_logic;
signal n1993 : std_logic;
signal n1992 : std_logic;
signal n1991 : std_logic;
signal \TX_DATA_6\ : std_logic;
signal n1990 : std_logic;
signal \TX_DATA_7\ : std_logic;
signal \ADV_B_c\ : std_logic;
signal \INVADV_R__i2C_net\ : std_logic;
signal n2587 : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_43\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_44\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_46\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_45\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_47\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_48\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_53\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_52\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_49\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_54\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_51\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_50\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_56\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_55\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_59\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_58\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_61\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_60\ : std_logic;
signal \line_buffer.n558\ : std_logic;
signal \line_buffer.n550\ : std_logic;
signal \line_buffer.n4101\ : std_logic;
signal n22 : std_logic;
signal \receive_module.rx_counter.n5_cascade_\ : std_logic;
signal \TVP_HSYNC_c\ : std_logic;
signal \receive_module.rx_counter.n4_adj_576\ : std_logic;
signal \RX_ADDR_0\ : std_logic;
signal \bfn_14_9_0_\ : std_logic;
signal \RX_ADDR_1\ : std_logic;
signal \receive_module.rx_counter.n3720\ : std_logic;
signal \RX_ADDR_2\ : std_logic;
signal \receive_module.rx_counter.n3721\ : std_logic;
signal \receive_module.rx_counter.n3722\ : std_logic;
signal \receive_module.rx_counter.n3723\ : std_logic;
signal \receive_module.rx_counter.n3724\ : std_logic;
signal \receive_module.rx_counter.n3725\ : std_logic;
signal \receive_module.rx_counter.n3726\ : std_logic;
signal \receive_module.rx_counter.n3727\ : std_logic;
signal \bfn_14_10_0_\ : std_logic;
signal \receive_module.rx_counter.n3728\ : std_logic;
signal n4214 : std_logic;
signal \RX_ADDR_11\ : std_logic;
signal \RX_ADDR_12\ : std_logic;
signal \DEBUG_c_5\ : std_logic;
signal \DEBUG_c_3\ : std_logic;
signal n658 : std_logic;
signal \transmit_module.X_DELTA_PATTERN_13\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_9\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_12\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_11\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_10\ : std_logic;
signal \line_buffer.n4072\ : std_logic;
signal \line_buffer.n4134\ : std_logic;
signal \transmit_module.n2361\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_2\ : std_logic;
signal \transmit_module.n219\ : std_logic;
signal \transmit_module.n179_cascade_\ : std_logic;
signal \transmit_module.n213\ : std_logic;
signal \transmit_module.n179\ : std_logic;
signal \transmit_module.n210\ : std_logic;
signal n19 : std_logic;
signal \transmit_module.n180\ : std_logic;
signal \transmit_module.n211\ : std_logic;
signal n20 : std_logic;
signal \transmit_module.old_VGA_HS\ : std_logic;
signal \ADV_HSYNC_c\ : std_logic;
signal \transmit_module.n181\ : std_logic;
signal \transmit_module.n212\ : std_logic;
signal \transmit_module.n181_cascade_\ : std_logic;
signal n21 : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_7\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_6\ : std_logic;
signal \transmit_module.n182\ : std_logic;
signal \receive_module.rx_counter.FRAME_COUNTER_0\ : std_logic;
signal \bfn_15_8_0_\ : std_logic;
signal \receive_module.rx_counter.FRAME_COUNTER_1\ : std_logic;
signal \receive_module.rx_counter.n3706\ : std_logic;
signal \receive_module.rx_counter.FRAME_COUNTER_2\ : std_logic;
signal \receive_module.rx_counter.n3707\ : std_logic;
signal \receive_module.rx_counter.FRAME_COUNTER_3\ : std_logic;
signal \receive_module.rx_counter.n3708\ : std_logic;
signal \receive_module.rx_counter.FRAME_COUNTER_4\ : std_logic;
signal \receive_module.rx_counter.n3709\ : std_logic;
signal \receive_module.rx_counter.n3710\ : std_logic;
signal \receive_module.rx_counter.FRAME_COUNTER_5\ : std_logic;
signal \receive_module.rx_counter.n2605\ : std_logic;
signal \receive_module.rx_counter.old_VS\ : std_logic;
signal \TVP_VSYNC_c\ : std_logic;
signal \receive_module.rx_counter.X_5\ : std_logic;
signal \receive_module.rx_counter.X_4\ : std_logic;
signal \receive_module.rx_counter.X_3\ : std_logic;
signal \receive_module.rx_counter.X_8\ : std_logic;
signal \receive_module.rx_counter.X_9\ : std_logic;
signal \receive_module.rx_counter.n4219\ : std_logic;
signal \receive_module.rx_counter.X_7\ : std_logic;
signal \receive_module.rx_counter.n4_adj_575_cascade_\ : std_logic;
signal \receive_module.rx_counter.X_6\ : std_logic;
signal \receive_module.rx_counter.O_VISIBLE_N_86\ : std_logic;
signal \receive_module.rx_counter.n11\ : std_logic;
signal \LED_c\ : std_logic;
signal \receive_module.rx_counter.n4222\ : std_logic;
signal \line_buffer.n623\ : std_logic;
signal \line_buffer.n615\ : std_logic;
signal \line_buffer.n4071\ : std_logic;
signal \line_buffer.n646\ : std_logic;
signal \line_buffer.n654\ : std_logic;
signal \line_buffer.n549\ : std_logic;
signal \line_buffer.n4176_cascade_\ : std_logic;
signal \line_buffer.n557\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_8\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_7\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_6\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_14\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_2\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_1\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_3\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_15\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_5\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_4\ : std_logic;
signal \transmit_module.n2315\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_0\ : std_logic;
signal \transmit_module.n204\ : std_logic;
signal \bfn_15_17_0_\ : std_logic;
signal \transmit_module.n3656\ : std_logic;
signal \transmit_module.TX_ADDR_2\ : std_logic;
signal \transmit_module.n202\ : std_logic;
signal \transmit_module.n3657\ : std_logic;
signal \transmit_module.n201\ : std_logic;
signal \transmit_module.n3658\ : std_logic;
signal \transmit_module.n3659\ : std_logic;
signal \transmit_module.n3660\ : std_logic;
signal \transmit_module.TX_ADDR_6\ : std_logic;
signal \transmit_module.n198\ : std_logic;
signal \transmit_module.n3661\ : std_logic;
signal \transmit_module.TX_ADDR_7\ : std_logic;
signal \transmit_module.n197\ : std_logic;
signal \transmit_module.n3662\ : std_logic;
signal \transmit_module.n3663\ : std_logic;
signal \transmit_module.n196\ : std_logic;
signal \bfn_15_18_0_\ : std_logic;
signal \transmit_module.n195\ : std_logic;
signal \transmit_module.n3664\ : std_logic;
signal \transmit_module.TX_ADDR_10\ : std_logic;
signal \transmit_module.n194\ : std_logic;
signal \transmit_module.n3665\ : std_logic;
signal \transmit_module.n3666\ : std_logic;
signal \transmit_module.n3667\ : std_logic;
signal \transmit_module.n3668\ : std_logic;
signal \transmit_module.TX_ADDR_8\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_8\ : std_logic;
signal \transmit_module.n203\ : std_logic;
signal \transmit_module.n218_cascade_\ : std_logic;
signal \transmit_module.n188\ : std_logic;
signal \transmit_module.TX_ADDR_0\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_0\ : std_logic;
signal \transmit_module.TX_ADDR_3\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_3\ : std_logic;
signal \transmit_module.n193\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_11\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_1\ : std_logic;
signal \transmit_module.TX_ADDR_1\ : std_logic;
signal \transmit_module.n187\ : std_logic;
signal \transmit_module.n218\ : std_logic;
signal n27 : std_logic;
signal \line_buffer.n678\ : std_logic;
signal \line_buffer.n686\ : std_logic;
signal \line_buffer.n614\ : std_logic;
signal \line_buffer.n4188_cascade_\ : std_logic;
signal \line_buffer.n622\ : std_logic;
signal \line_buffer.n4191_cascade_\ : std_logic;
signal \line_buffer.n4179\ : std_logic;
signal \TX_DATA_5\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_18\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_21\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_20\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_19\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_1\ : std_logic;
signal \transmit_module.TX_ADDR_9\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_9\ : std_logic;
signal \transmit_module.n200\ : std_logic;
signal \transmit_module.n215_cascade_\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_5\ : std_logic;
signal \transmit_module.n191\ : std_logic;
signal \transmit_module.BRAM_ADDR_13_N_258_13\ : std_logic;
signal \transmit_module.n199\ : std_logic;
signal \transmit_module.n3910\ : std_logic;
signal \transmit_module.n214_cascade_\ : std_logic;
signal \transmit_module.TX_ADDR_5\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_4\ : std_logic;
signal \transmit_module.TX_ADDR_4\ : std_logic;
signal \transmit_module.n184\ : std_logic;
signal \transmit_module.n215\ : std_logic;
signal n24 : std_logic;
signal \transmit_module.n183\ : std_logic;
signal \transmit_module.n214\ : std_logic;
signal n23 : std_logic;
signal \transmit_module.n4220\ : std_logic;
signal \transmit_module.n192\ : std_logic;
signal \transmit_module.n3926\ : std_logic;
signal \transmit_module.n2277\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_42\ : std_logic;
signal \DEBUG_c_1_c\ : std_logic;
signal \GB_BUFFER_DEBUG_c_1_c_THRU_CO\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_29\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_31\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_30\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_12\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_32\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_13\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_14\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_26\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_25\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_28\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_27\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_0\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_99\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_37\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_36\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_38\ : std_logic;
signal \transmit_module.n185\ : std_logic;
signal \transmit_module.n216\ : std_logic;
signal \transmit_module.n4211\ : std_logic;
signal n25 : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_12\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_13\ : std_logic;
signal \transmit_module.n2305\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_39\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_41\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_40\ : std_logic;
signal \line_buffer.n620\ : std_logic;
signal \line_buffer.n612\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_6\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_5\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_7\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_11\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_10\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_9\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_8\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_15\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_4\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_17\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_16\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_3\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_2\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_22\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_24\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_23\ : std_logic;
signal \transmit_module.n4224\ : std_logic;
signal \line_buffer.n642\ : std_logic;
signal \line_buffer.n650\ : std_logic;
signal \line_buffer.n545\ : std_logic;
signal \line_buffer.n4164_cascade_\ : std_logic;
signal \line_buffer.n553\ : std_logic;
signal \line_buffer.n4167_cascade_\ : std_logic;
signal \TX_DATA_1\ : std_logic;
signal \line_buffer.n4065\ : std_logic;
signal \line_buffer.n684\ : std_logic;
signal \line_buffer.n676\ : std_logic;
signal \line_buffer.n4066\ : std_logic;
signal \line_buffer.n555\ : std_logic;
signal \line_buffer.n547\ : std_logic;
signal \line_buffer.n4074_cascade_\ : std_logic;
signal \line_buffer.n4128\ : std_logic;
signal \TX_DATA_3\ : std_logic;
signal \line_buffer.n652\ : std_logic;
signal \line_buffer.n644\ : std_logic;
signal \line_buffer.n4075\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_33\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_35\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_34\ : std_logic;
signal \transmit_module.n4225\ : std_logic;
signal \ADV_VSYNC_c\ : std_logic;
signal \line_buffer.n617\ : std_logic;
signal \line_buffer.n609\ : std_logic;
signal \line_buffer.n610\ : std_logic;
signal \line_buffer.n618\ : std_logic;
signal \line_buffer.n4161\ : std_logic;
signal \line_buffer.n673\ : std_logic;
signal \line_buffer.n681\ : std_logic;
signal \line_buffer.n4146\ : std_logic;
signal \line_buffer.n4149\ : std_logic;
signal \TX_DATA_0\ : std_logic;
signal \line_buffer.n621\ : std_logic;
signal \line_buffer.n613\ : std_logic;
signal \line_buffer.n653\ : std_logic;
signal \line_buffer.n645\ : std_logic;
signal \line_buffer.n4062\ : std_logic;
signal \line_buffer.n4078\ : std_logic;
signal \DEBUG_c_2\ : std_logic;
signal \line_buffer.n4140\ : std_logic;
signal \TX_DATA_4\ : std_logic;
signal \ADV_CLK_c\ : std_logic;
signal \line_buffer.n641\ : std_logic;
signal \line_buffer.n649\ : std_logic;
signal \line_buffer.n552\ : std_logic;
signal \line_buffer.n4116\ : std_logic;
signal \line_buffer.n544\ : std_logic;
signal \line_buffer.n4119\ : std_logic;
signal \line_buffer.n548\ : std_logic;
signal \line_buffer.n556\ : std_logic;
signal \line_buffer.n4077\ : std_logic;
signal \line_buffer.n674\ : std_logic;
signal \TX_ADDR_12\ : std_logic;
signal \line_buffer.n682\ : std_logic;
signal \line_buffer.n4158\ : std_logic;
signal \line_buffer.n685\ : std_logic;
signal \line_buffer.n677\ : std_logic;
signal \TX_ADDR_11\ : std_logic;
signal \line_buffer.n4063\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \TVP_CLK_wire\ : std_logic;
signal \ADV_CLK_wire\ : std_logic;
signal \TVP_VIDEO_wire\ : std_logic_vector(9 downto 0);
signal \ADV_G_wire\ : std_logic_vector(7 downto 0);
signal \ADV_R_wire\ : std_logic_vector(7 downto 0);
signal \ADV_B_wire\ : std_logic_vector(7 downto 0);
signal \ADV_SYNC_N_wire\ : std_logic;
signal \TVP_HSYNC_wire\ : std_logic;
signal \TVP_VSYNC_wire\ : std_logic;
signal \ADV_BLANK_N_wire\ : std_logic;
signal \LED_wire\ : std_logic;
signal \ADV_HSYNC_wire\ : std_logic;
signal \ADV_VSYNC_wire\ : std_logic;
signal \tx_pll.TX_PLL_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);
signal \line_buffer.mem2_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem2_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem2_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem2_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem2_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem14_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem14_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem14_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem14_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem14_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem5_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem5_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem5_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem5_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem5_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem11_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem11_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem11_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem11_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem11_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem21_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem21_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem21_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem21_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem21_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem12_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem12_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem12_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem12_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem12_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem18_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem18_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem18_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem18_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem18_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem24_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem24_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem24_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem24_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem24_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem15_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem15_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem15_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem15_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem15_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem27_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem27_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem27_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem27_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem27_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem4_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem4_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem4_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem4_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem4_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem16_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem16_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem16_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem16_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem16_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem30_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem30_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem30_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem30_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem30_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem7_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem7_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem7_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem7_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem7_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem20_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem20_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem20_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem20_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem20_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem13_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem13_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem13_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem13_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem13_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem19_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem19_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem19_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem19_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem19_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem23_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem23_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem23_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem23_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem23_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem26_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem26_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem26_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem26_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem26_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem3_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem3_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem3_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem3_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem3_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem17_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem17_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem17_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem17_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem17_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem31_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem31_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem31_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem31_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem31_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem9_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem9_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem9_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem9_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem9_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem29_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem29_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem29_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem29_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem29_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem6_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem6_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem6_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem6_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem6_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem10_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem10_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem10_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem10_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem10_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem22_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem22_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem22_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem22_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem22_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem25_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem25_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem25_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem25_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem25_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem8_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem8_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem8_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem8_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem8_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem28_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem28_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem28_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem28_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem28_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    \TVP_CLK_wire\ <= TVP_CLK;
    ADV_CLK <= \ADV_CLK_wire\;
    \TVP_VIDEO_wire\ <= TVP_VIDEO;
    ADV_G <= \ADV_G_wire\;
    ADV_R <= \ADV_R_wire\;
    ADV_B <= \ADV_B_wire\;
    ADV_SYNC_N <= \ADV_SYNC_N_wire\;
    \TVP_HSYNC_wire\ <= TVP_HSYNC;
    \TVP_VSYNC_wire\ <= TVP_VSYNC;
    ADV_BLANK_N <= \ADV_BLANK_N_wire\;
    LED <= \LED_wire\;
    ADV_HSYNC <= \ADV_HSYNC_wire\;
    ADV_VSYNC <= \ADV_VSYNC_wire\;
    \tx_pll.TX_PLL_inst_DYNAMICDELAY_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.n559\ <= \line_buffer.mem2_physical_RDATA_wire\(11);
    \line_buffer.n558\ <= \line_buffer.mem2_physical_RDATA_wire\(3);
    \line_buffer.mem2_physical_RADDR_wire\ <= \N__9840\&\N__16167\&\N__16833\&\N__16497\&\N__15513\&\N__18567\&\N__18801\&\N__19971\&\N__13950\&\N__18126\&\N__10740\;
    \line_buffer.mem2_physical_WADDR_wire\ <= \N__12804\&\N__13062\&\N__11814\&\N__12072\&\N__12339\&\N__11067\&\N__11292\&\N__11526\&\N__14790\&\N__15021\&\N__15252\;
    \line_buffer.mem2_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem2_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8743\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8855\&'0'&'0'&'0';
    \line_buffer.n646\ <= \line_buffer.mem14_physical_RDATA_wire\(11);
    \line_buffer.n645\ <= \line_buffer.mem14_physical_RDATA_wire\(3);
    \line_buffer.mem14_physical_RADDR_wire\ <= \N__9912\&\N__16239\&\N__16905\&\N__16569\&\N__15585\&\N__18639\&\N__18873\&\N__20043\&\N__14022\&\N__18198\&\N__10812\;
    \line_buffer.mem14_physical_WADDR_wire\ <= \N__12876\&\N__13134\&\N__11886\&\N__12144\&\N__12411\&\N__11139\&\N__11364\&\N__11598\&\N__14862\&\N__15093\&\N__15324\;
    \line_buffer.mem14_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem14_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8666\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8536\&'0'&'0'&'0';
    \line_buffer.n656\ <= \line_buffer.mem5_physical_RDATA_wire\(11);
    \line_buffer.n655\ <= \line_buffer.mem5_physical_RDATA_wire\(3);
    \line_buffer.mem5_physical_RADDR_wire\ <= \N__9843\&\N__16176\&\N__16842\&\N__16506\&\N__15516\&\N__18582\&\N__18810\&\N__19986\&\N__13965\&\N__18129\&\N__10737\;
    \line_buffer.mem5_physical_WADDR_wire\ <= \N__12825\&\N__13077\&\N__11829\&\N__12081\&\N__12336\&\N__11076\&\N__11295\&\N__11523\&\N__14793\&\N__15030\&\N__15267\;
    \line_buffer.mem5_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem5_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8765\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8876\&'0'&'0'&'0';
    \line_buffer.n614\ <= \line_buffer.mem11_physical_RDATA_wire\(11);
    \line_buffer.n613\ <= \line_buffer.mem11_physical_RDATA_wire\(3);
    \line_buffer.mem11_physical_RADDR_wire\ <= \N__9948\&\N__16275\&\N__16941\&\N__16605\&\N__15621\&\N__18675\&\N__18909\&\N__20079\&\N__14058\&\N__18234\&\N__10848\;
    \line_buffer.mem11_physical_WADDR_wire\ <= \N__12912\&\N__13170\&\N__11922\&\N__12180\&\N__12447\&\N__11175\&\N__11400\&\N__11634\&\N__14898\&\N__15129\&\N__15360\;
    \line_buffer.mem11_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem11_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8626\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8515\&'0'&'0'&'0';
    \line_buffer.n676\ <= \line_buffer.mem21_physical_RDATA_wire\(11);
    \line_buffer.n675\ <= \line_buffer.mem21_physical_RDATA_wire\(3);
    \line_buffer.mem21_physical_RADDR_wire\ <= \N__9816\&\N__16143\&\N__16809\&\N__16473\&\N__15489\&\N__18543\&\N__18777\&\N__19947\&\N__13926\&\N__18102\&\N__10716\;
    \line_buffer.mem21_physical_WADDR_wire\ <= \N__12780\&\N__13038\&\N__11790\&\N__12048\&\N__12315\&\N__11043\&\N__11268\&\N__11502\&\N__14766\&\N__14997\&\N__15228\;
    \line_buffer.mem21_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem21_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8447\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8347\&'0'&'0'&'0';
    \line_buffer.n612\ <= \line_buffer.mem12_physical_RDATA_wire\(11);
    \line_buffer.n611\ <= \line_buffer.mem12_physical_RDATA_wire\(3);
    \line_buffer.mem12_physical_RADDR_wire\ <= \N__9936\&\N__16263\&\N__16929\&\N__16593\&\N__15609\&\N__18663\&\N__18897\&\N__20067\&\N__14046\&\N__18222\&\N__10836\;
    \line_buffer.mem12_physical_WADDR_wire\ <= \N__12900\&\N__13158\&\N__11910\&\N__12168\&\N__12435\&\N__11163\&\N__11388\&\N__11622\&\N__14886\&\N__15117\&\N__15348\;
    \line_buffer.mem12_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem12_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8417\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8335\&'0'&'0'&'0';
    \line_buffer.n555\ <= \line_buffer.mem18_physical_RDATA_wire\(11);
    \line_buffer.n554\ <= \line_buffer.mem18_physical_RDATA_wire\(3);
    \line_buffer.mem18_physical_RADDR_wire\ <= \N__9864\&\N__16191\&\N__16857\&\N__16521\&\N__15537\&\N__18591\&\N__18825\&\N__19995\&\N__13974\&\N__18150\&\N__10764\;
    \line_buffer.mem18_physical_WADDR_wire\ <= \N__12828\&\N__13086\&\N__11838\&\N__12096\&\N__12363\&\N__11091\&\N__11316\&\N__11550\&\N__14814\&\N__15045\&\N__15276\;
    \line_buffer.mem18_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem18_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8451\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8336\&'0'&'0'&'0';
    \line_buffer.n620\ <= \line_buffer.mem24_physical_RDATA_wire\(11);
    \line_buffer.n619\ <= \line_buffer.mem24_physical_RDATA_wire\(3);
    \line_buffer.mem24_physical_RADDR_wire\ <= \N__9963\&\N__16296\&\N__16962\&\N__16626\&\N__15636\&\N__18702\&\N__18930\&\N__20106\&\N__14085\&\N__18249\&\N__10857\;
    \line_buffer.mem24_physical_WADDR_wire\ <= \N__12945\&\N__13197\&\N__11949\&\N__12201\&\N__12456\&\N__11196\&\N__11415\&\N__11643\&\N__14913\&\N__15150\&\N__15387\;
    \line_buffer.mem24_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem24_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8380\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8258\&'0'&'0'&'0';
    \line_buffer.n648\ <= \line_buffer.mem1_physical_RDATA_wire\(11);
    \line_buffer.n647\ <= \line_buffer.mem1_physical_RDATA_wire\(3);
    \line_buffer.mem1_physical_RADDR_wire\ <= \N__9972\&\N__16299\&\N__16965\&\N__16629\&\N__15645\&\N__18699\&\N__18933\&\N__20103\&\N__14082\&\N__18258\&\N__10870\;
    \line_buffer.mem1_physical_WADDR_wire\ <= \N__12936\&\N__13194\&\N__11946\&\N__12204\&\N__12469\&\N__11199\&\N__11424\&\N__11656\&\N__14922\&\N__15153\&\N__15384\;
    \line_buffer.mem1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8722\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8840\&'0'&'0'&'0';
    \line_buffer.n644\ <= \line_buffer.mem15_physical_RDATA_wire\(11);
    \line_buffer.n643\ <= \line_buffer.mem15_physical_RDATA_wire\(3);
    \line_buffer.mem15_physical_RADDR_wire\ <= \N__9900\&\N__16227\&\N__16893\&\N__16557\&\N__15573\&\N__18627\&\N__18861\&\N__20031\&\N__14010\&\N__18186\&\N__10800\;
    \line_buffer.mem15_physical_WADDR_wire\ <= \N__12864\&\N__13122\&\N__11874\&\N__12132\&\N__12399\&\N__11127\&\N__11352\&\N__11586\&\N__14850\&\N__15081\&\N__15312\;
    \line_buffer.mem15_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem15_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8433\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8325\&'0'&'0'&'0';
    \line_buffer.n652\ <= \line_buffer.mem27_physical_RDATA_wire\(11);
    \line_buffer.n651\ <= \line_buffer.mem27_physical_RDATA_wire\(3);
    \line_buffer.mem27_physical_RADDR_wire\ <= \N__9927\&\N__16260\&\N__16926\&\N__16590\&\N__15600\&\N__18666\&\N__18894\&\N__20070\&\N__14049\&\N__18213\&\N__10821\;
    \line_buffer.mem27_physical_WADDR_wire\ <= \N__12909\&\N__13161\&\N__11913\&\N__12165\&\N__12420\&\N__11160\&\N__11379\&\N__11607\&\N__14877\&\N__15114\&\N__15351\;
    \line_buffer.mem27_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem27_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8411\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8289\&'0'&'0'&'0';
    \line_buffer.n624\ <= \line_buffer.mem4_physical_RDATA_wire\(11);
    \line_buffer.n623\ <= \line_buffer.mem4_physical_RDATA_wire\(3);
    \line_buffer.mem4_physical_RADDR_wire\ <= \N__9855\&\N__16188\&\N__16854\&\N__16518\&\N__15528\&\N__18594\&\N__18822\&\N__19998\&\N__13977\&\N__18141\&\N__10749\;
    \line_buffer.mem4_physical_WADDR_wire\ <= \N__12837\&\N__13089\&\N__11841\&\N__12093\&\N__12348\&\N__11088\&\N__11307\&\N__11535\&\N__14805\&\N__15042\&\N__15279\;
    \line_buffer.mem4_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem4_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8750\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8875\&'0'&'0'&'0';
    \line_buffer.n642\ <= \line_buffer.mem16_physical_RDATA_wire\(11);
    \line_buffer.n641\ <= \line_buffer.mem16_physical_RDATA_wire\(3);
    \line_buffer.mem16_physical_RADDR_wire\ <= \N__9888\&\N__16215\&\N__16881\&\N__16545\&\N__15561\&\N__18615\&\N__18849\&\N__20019\&\N__13998\&\N__18174\&\N__10788\;
    \line_buffer.mem16_physical_WADDR_wire\ <= \N__12852\&\N__13110\&\N__11862\&\N__12120\&\N__12387\&\N__11115\&\N__11340\&\N__11574\&\N__14838\&\N__15069\&\N__15300\;
    \line_buffer.mem16_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem16_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8214\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8997\&'0'&'0'&'0';
    \line_buffer.n684\ <= \line_buffer.mem30_physical_RDATA_wire\(11);
    \line_buffer.n683\ <= \line_buffer.mem30_physical_RDATA_wire\(3);
    \line_buffer.mem30_physical_RADDR_wire\ <= \N__9879\&\N__16212\&\N__16878\&\N__16542\&\N__15552\&\N__18618\&\N__18846\&\N__20022\&\N__14001\&\N__18165\&\N__10773\;
    \line_buffer.mem30_physical_WADDR_wire\ <= \N__12861\&\N__13113\&\N__11865\&\N__12117\&\N__12372\&\N__11112\&\N__11331\&\N__11559\&\N__14829\&\N__15066\&\N__15303\;
    \line_buffer.mem30_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem30_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8440\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8321\&'0'&'0'&'0';
    \line_buffer.n551\ <= \line_buffer.mem7_physical_RDATA_wire\(11);
    \line_buffer.n550\ <= \line_buffer.mem7_physical_RDATA_wire\(3);
    \line_buffer.mem7_physical_RADDR_wire\ <= \N__9819\&\N__16152\&\N__16818\&\N__16482\&\N__15492\&\N__18558\&\N__18786\&\N__19962\&\N__13941\&\N__18105\&\N__10713\;
    \line_buffer.mem7_physical_WADDR_wire\ <= \N__12801\&\N__13053\&\N__11805\&\N__12057\&\N__12312\&\N__11052\&\N__11271\&\N__11499\&\N__14769\&\N__15006\&\N__15243\;
    \line_buffer.mem7_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem7_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8773\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8884\&'0'&'0'&'0';
    \line_buffer.n678\ <= \line_buffer.mem20_physical_RDATA_wire\(11);
    \line_buffer.n677\ <= \line_buffer.mem20_physical_RDATA_wire\(3);
    \line_buffer.mem20_physical_RADDR_wire\ <= \N__9828\&\N__16155\&\N__16821\&\N__16485\&\N__15501\&\N__18555\&\N__18789\&\N__19959\&\N__13938\&\N__18114\&\N__10728\;
    \line_buffer.mem20_physical_WADDR_wire\ <= \N__12792\&\N__13050\&\N__11802\&\N__12060\&\N__12327\&\N__11055\&\N__11280\&\N__11514\&\N__14778\&\N__15009\&\N__15240\;
    \line_buffer.mem20_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem20_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8665\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8557\&'0'&'0'&'0';
    \line_buffer.n610\ <= \line_buffer.mem13_physical_RDATA_wire\(11);
    \line_buffer.n609\ <= \line_buffer.mem13_physical_RDATA_wire\(3);
    \line_buffer.mem13_physical_RADDR_wire\ <= \N__9924\&\N__16251\&\N__16917\&\N__16581\&\N__15597\&\N__18651\&\N__18885\&\N__20055\&\N__14034\&\N__18210\&\N__10824\;
    \line_buffer.mem13_physical_WADDR_wire\ <= \N__12888\&\N__13146\&\N__11898\&\N__12156\&\N__12423\&\N__11151\&\N__11376\&\N__11610\&\N__14874\&\N__15105\&\N__15336\;
    \line_buffer.mem13_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem13_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8193\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8990\&'0'&'0'&'0';
    \line_buffer.n553\ <= \line_buffer.mem19_physical_RDATA_wire\(11);
    \line_buffer.n552\ <= \line_buffer.mem19_physical_RDATA_wire\(3);
    \line_buffer.mem19_physical_RADDR_wire\ <= \N__9852\&\N__16179\&\N__16845\&\N__16509\&\N__15525\&\N__18579\&\N__18813\&\N__19983\&\N__13962\&\N__18138\&\N__10752\;
    \line_buffer.mem19_physical_WADDR_wire\ <= \N__12816\&\N__13074\&\N__11826\&\N__12084\&\N__12351\&\N__11079\&\N__11304\&\N__11538\&\N__14802\&\N__15033\&\N__15264\;
    \line_buffer.mem19_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem19_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8206\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__9009\&'0'&'0'&'0';
    \line_buffer.n622\ <= \line_buffer.mem23_physical_RDATA_wire\(11);
    \line_buffer.n621\ <= \line_buffer.mem23_physical_RDATA_wire\(3);
    \line_buffer.mem23_physical_RADDR_wire\ <= \N__9975\&\N__16308\&\N__16974\&\N__16638\&\N__15648\&\N__18712\&\N__18942\&\N__20116\&\N__14095\&\N__18261\&\N__10869\;
    \line_buffer.mem23_physical_WADDR_wire\ <= \N__12952\&\N__13207\&\N__11959\&\N__12213\&\N__12468\&\N__11208\&\N__11427\&\N__11655\&\N__14925\&\N__15162\&\N__15397\;
    \line_buffer.mem23_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem23_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8642\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8483\&'0'&'0'&'0';
    \line_buffer.n616\ <= \line_buffer.mem0_physical_RDATA_wire\(11);
    \line_buffer.n615\ <= \line_buffer.mem0_physical_RDATA_wire\(3);
    \line_buffer.mem0_physical_RADDR_wire\ <= \N__9979\&\N__16309\&\N__16975\&\N__16639\&\N__15652\&\N__18711\&\N__18943\&\N__20115\&\N__14094\&\N__18265\&\N__10876\;
    \line_buffer.mem0_physical_WADDR_wire\ <= \N__12948\&\N__13206\&\N__11958\&\N__12214\&\N__12475\&\N__11209\&\N__11431\&\N__11662\&\N__14929\&\N__15163\&\N__15396\;
    \line_buffer.mem0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8697\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8839\&'0'&'0'&'0';
    \line_buffer.n654\ <= \line_buffer.mem26_physical_RDATA_wire\(11);
    \line_buffer.n653\ <= \line_buffer.mem26_physical_RDATA_wire\(3);
    \line_buffer.mem26_physical_RADDR_wire\ <= \N__9939\&\N__16272\&\N__16938\&\N__16602\&\N__15612\&\N__18678\&\N__18906\&\N__20082\&\N__14061\&\N__18225\&\N__10833\;
    \line_buffer.mem26_physical_WADDR_wire\ <= \N__12921\&\N__13173\&\N__11925\&\N__12177\&\N__12432\&\N__11172\&\N__11391\&\N__11619\&\N__14889\&\N__15126\&\N__15363\;
    \line_buffer.mem26_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem26_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8625\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8508\&'0'&'0'&'0';
    \line_buffer.n680\ <= \line_buffer.mem3_physical_RDATA_wire\(11);
    \line_buffer.n679\ <= \line_buffer.mem3_physical_RDATA_wire\(3);
    \line_buffer.mem3_physical_RADDR_wire\ <= \N__9891\&\N__16224\&\N__16890\&\N__16554\&\N__15564\&\N__18630\&\N__18858\&\N__20034\&\N__14013\&\N__18177\&\N__10785\;
    \line_buffer.mem3_physical_WADDR_wire\ <= \N__12873\&\N__13125\&\N__11877\&\N__12129\&\N__12384\&\N__11124\&\N__11343\&\N__11571\&\N__14841\&\N__15078\&\N__15315\;
    \line_buffer.mem3_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem3_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8751\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8856\&'0'&'0'&'0';
    \line_buffer.n557\ <= \line_buffer.mem17_physical_RDATA_wire\(11);
    \line_buffer.n556\ <= \line_buffer.mem17_physical_RDATA_wire\(3);
    \line_buffer.mem17_physical_RADDR_wire\ <= \N__9876\&\N__16203\&\N__16869\&\N__16533\&\N__15549\&\N__18603\&\N__18837\&\N__20007\&\N__13986\&\N__18162\&\N__10776\;
    \line_buffer.mem17_physical_WADDR_wire\ <= \N__12840\&\N__13098\&\N__11850\&\N__12108\&\N__12375\&\N__11103\&\N__11328\&\N__11562\&\N__14826\&\N__15057\&\N__15288\;
    \line_buffer.mem17_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem17_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8649\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8546\&'0'&'0'&'0';
    \line_buffer.n682\ <= \line_buffer.mem31_physical_RDATA_wire\(11);
    \line_buffer.n681\ <= \line_buffer.mem31_physical_RDATA_wire\(3);
    \line_buffer.mem31_physical_RADDR_wire\ <= \N__9867\&\N__16200\&\N__16866\&\N__16530\&\N__15540\&\N__18606\&\N__18834\&\N__20010\&\N__13989\&\N__18153\&\N__10761\;
    \line_buffer.mem31_physical_WADDR_wire\ <= \N__12849\&\N__13101\&\N__11853\&\N__12105\&\N__12360\&\N__11100\&\N__11319\&\N__11547\&\N__14817\&\N__15054\&\N__15291\;
    \line_buffer.mem31_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem31_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8183\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8974\&'0'&'0'&'0';
    \line_buffer.n547\ <= \line_buffer.mem9_physical_RDATA_wire\(11);
    \line_buffer.n546\ <= \line_buffer.mem9_physical_RDATA_wire\(3);
    \line_buffer.mem9_physical_RADDR_wire\ <= \N__9795\&\N__16128\&\N__16794\&\N__16458\&\N__15468\&\N__18534\&\N__18762\&\N__19938\&\N__13917\&\N__18081\&\N__10689\;
    \line_buffer.mem9_physical_WADDR_wire\ <= \N__12777\&\N__13029\&\N__11781\&\N__12033\&\N__12288\&\N__11028\&\N__11247\&\N__11475\&\N__14745\&\N__14982\&\N__15219\;
    \line_buffer.mem9_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem9_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8455\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8346\&'0'&'0'&'0';
    \line_buffer.n686\ <= \line_buffer.mem29_physical_RDATA_wire\(11);
    \line_buffer.n685\ <= \line_buffer.mem29_physical_RDATA_wire\(3);
    \line_buffer.mem29_physical_RADDR_wire\ <= \N__9903\&\N__16236\&\N__16902\&\N__16566\&\N__15576\&\N__18642\&\N__18870\&\N__20046\&\N__14025\&\N__18189\&\N__10797\;
    \line_buffer.mem29_physical_WADDR_wire\ <= \N__12885\&\N__13137\&\N__11889\&\N__12141\&\N__12396\&\N__11136\&\N__11355\&\N__11583\&\N__14853\&\N__15090\&\N__15327\;
    \line_buffer.mem29_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem29_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8667\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8521\&'0'&'0'&'0';
    \line_buffer.n688\ <= \line_buffer.mem6_physical_RDATA_wire\(11);
    \line_buffer.n687\ <= \line_buffer.mem6_physical_RDATA_wire\(3);
    \line_buffer.mem6_physical_RADDR_wire\ <= \N__9831\&\N__16164\&\N__16830\&\N__16494\&\N__15504\&\N__18570\&\N__18798\&\N__19974\&\N__13953\&\N__18117\&\N__10725\;
    \line_buffer.mem6_physical_WADDR_wire\ <= \N__12813\&\N__13065\&\N__11817\&\N__12069\&\N__12324\&\N__11064\&\N__11283\&\N__11511\&\N__14781\&\N__15018\&\N__15255\;
    \line_buffer.mem6_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem6_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8772\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8883\&'0'&'0'&'0';
    \line_buffer.n545\ <= \line_buffer.mem10_physical_RDATA_wire\(11);
    \line_buffer.n544\ <= \line_buffer.mem10_physical_RDATA_wire\(3);
    \line_buffer.mem10_physical_RADDR_wire\ <= \N__9960\&\N__16287\&\N__16953\&\N__16617\&\N__15633\&\N__18687\&\N__18921\&\N__20091\&\N__14070\&\N__18246\&\N__10860\;
    \line_buffer.mem10_physical_WADDR_wire\ <= \N__12924\&\N__13182\&\N__11934\&\N__12192\&\N__12459\&\N__11187\&\N__11412\&\N__11646\&\N__14910\&\N__15141\&\N__15372\;
    \line_buffer.mem10_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem10_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8207\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8975\&'0'&'0'&'0';
    \line_buffer.n674\ <= \line_buffer.mem22_physical_RDATA_wire\(11);
    \line_buffer.n673\ <= \line_buffer.mem22_physical_RDATA_wire\(3);
    \line_buffer.mem22_physical_RADDR_wire\ <= \N__9804\&\N__16131\&\N__16797\&\N__16461\&\N__15477\&\N__18531\&\N__18765\&\N__19935\&\N__13914\&\N__18090\&\N__10704\;
    \line_buffer.mem22_physical_WADDR_wire\ <= \N__12768\&\N__13026\&\N__11778\&\N__12036\&\N__12303\&\N__11031\&\N__11256\&\N__11490\&\N__14754\&\N__14985\&\N__15216\;
    \line_buffer.mem22_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem22_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8215\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__9016\&'0'&'0'&'0';
    \line_buffer.n618\ <= \line_buffer.mem25_physical_RDATA_wire\(11);
    \line_buffer.n617\ <= \line_buffer.mem25_physical_RDATA_wire\(3);
    \line_buffer.mem25_physical_RADDR_wire\ <= \N__9951\&\N__16284\&\N__16950\&\N__16614\&\N__15624\&\N__18690\&\N__18918\&\N__20094\&\N__14073\&\N__18237\&\N__10845\;
    \line_buffer.mem25_physical_WADDR_wire\ <= \N__12933\&\N__13185\&\N__11937\&\N__12189\&\N__12444\&\N__11184\&\N__11403\&\N__11631\&\N__14901\&\N__15138\&\N__15375\;
    \line_buffer.mem25_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem25_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8182\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8941\&'0'&'0'&'0';
    \line_buffer.n549\ <= \line_buffer.mem8_physical_RDATA_wire\(11);
    \line_buffer.n548\ <= \line_buffer.mem8_physical_RDATA_wire\(3);
    \line_buffer.mem8_physical_RADDR_wire\ <= \N__9807\&\N__16140\&\N__16806\&\N__16470\&\N__15480\&\N__18546\&\N__18774\&\N__19950\&\N__13929\&\N__18093\&\N__10701\;
    \line_buffer.mem8_physical_WADDR_wire\ <= \N__12789\&\N__13041\&\N__11793\&\N__12045\&\N__12300\&\N__11040\&\N__11259\&\N__11487\&\N__14757\&\N__14994\&\N__15231\;
    \line_buffer.mem8_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem8_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8671\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8556\&'0'&'0'&'0';
    \line_buffer.n650\ <= \line_buffer.mem28_physical_RDATA_wire\(11);
    \line_buffer.n649\ <= \line_buffer.mem28_physical_RDATA_wire\(3);
    \line_buffer.mem28_physical_RADDR_wire\ <= \N__9915\&\N__16248\&\N__16914\&\N__16578\&\N__15588\&\N__18654\&\N__18882\&\N__20058\&\N__14037\&\N__18201\&\N__10809\;
    \line_buffer.mem28_physical_WADDR_wire\ <= \N__12897\&\N__13149\&\N__11901\&\N__12153\&\N__12408\&\N__11148\&\N__11367\&\N__11595\&\N__14865\&\N__15102\&\N__15339\;
    \line_buffer.mem28_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem28_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8175\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__8954\&'0'&'0'&'0';

    \tx_pll.TX_PLL_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "010",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "100",
            DIVF => "0100110",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            LATCHINPUTVALUE => '0',
            SCLK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => \ADV_CLK_c\,
            REFERENCECLK => \N__19215\,
            RESETB => \N__23324\,
            BYPASS => \GNDG0\,
            SDI => '0',
            DYNAMICDELAY => \tx_pll.TX_PLL_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => OPEN
        );

    \line_buffer.mem2_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem2_physical_RDATA_wire\,
            RADDR => \line_buffer.mem2_physical_RADDR_wire\,
            WADDR => \line_buffer.mem2_physical_WADDR_wire\,
            MASK => \line_buffer.mem2_physical_MASK_wire\,
            WDATA => \line_buffer.mem2_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22387\,
            RE => \N__23189\,
            WCLKE => 'H',
            WCLK => \N__19361\,
            WE => \N__12610\
        );

    \line_buffer.mem14_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem14_physical_RDATA_wire\,
            RADDR => \line_buffer.mem14_physical_RADDR_wire\,
            WADDR => \line_buffer.mem14_physical_WADDR_wire\,
            MASK => \line_buffer.mem14_physical_MASK_wire\,
            WDATA => \line_buffer.mem14_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22623\,
            RE => \N__23261\,
            WCLKE => 'H',
            WCLK => \N__19346\,
            WE => \N__15712\
        );

    \line_buffer.mem5_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem5_physical_RDATA_wire\,
            RADDR => \line_buffer.mem5_physical_RADDR_wire\,
            WADDR => \line_buffer.mem5_physical_WADDR_wire\,
            MASK => \line_buffer.mem5_physical_MASK_wire\,
            WDATA => \line_buffer.mem5_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__21959\,
            RE => \N__23281\,
            WCLKE => 'H',
            WCLK => \N__19360\,
            WE => \N__10120\
        );

    \line_buffer.mem11_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem11_physical_RDATA_wire\,
            RADDR => \line_buffer.mem11_physical_RADDR_wire\,
            WADDR => \line_buffer.mem11_physical_WADDR_wire\,
            MASK => \line_buffer.mem11_physical_MASK_wire\,
            WDATA => \line_buffer.mem11_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22676\,
            RE => \N__23344\,
            WCLKE => 'H',
            WCLK => \N__19333\,
            WE => \N__10227\
        );

    \line_buffer.mem21_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem21_physical_RDATA_wire\,
            RADDR => \line_buffer.mem21_physical_RADDR_wire\,
            WADDR => \line_buffer.mem21_physical_WADDR_wire\,
            MASK => \line_buffer.mem21_physical_MASK_wire\,
            WDATA => \line_buffer.mem21_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22386\,
            RE => \N__23138\,
            WCLKE => 'H',
            WCLK => \N__19365\,
            WE => \N__13486\
        );

    \line_buffer.mem12_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem12_physical_RDATA_wire\,
            RADDR => \line_buffer.mem12_physical_RADDR_wire\,
            WADDR => \line_buffer.mem12_physical_WADDR_wire\,
            MASK => \line_buffer.mem12_physical_MASK_wire\,
            WDATA => \line_buffer.mem12_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22655\,
            RE => \N__23311\,
            WCLKE => 'H',
            WCLK => \N__19341\,
            WE => \N__10226\
        );

    \line_buffer.mem18_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem18_physical_RDATA_wire\,
            RADDR => \line_buffer.mem18_physical_RADDR_wire\,
            WADDR => \line_buffer.mem18_physical_WADDR_wire\,
            MASK => \line_buffer.mem18_physical_MASK_wire\,
            WDATA => \line_buffer.mem18_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22516\,
            RE => \N__23124\,
            WCLKE => 'H',
            WCLK => \N__19354\,
            WE => \N__12606\
        );

    \line_buffer.mem24_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem24_physical_RDATA_wire\,
            RADDR => \line_buffer.mem24_physical_RADDR_wire\,
            WADDR => \line_buffer.mem24_physical_WADDR_wire\,
            MASK => \line_buffer.mem24_physical_MASK_wire\,
            WDATA => \line_buffer.mem24_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22407\,
            RE => \N__23394\,
            WCLKE => 'H',
            WCLK => \N__19328\,
            WE => \N__12656\
        );

    \line_buffer.mem1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem1_physical_RDATA_wire\,
            RADDR => \line_buffer.mem1_physical_RADDR_wire\,
            WADDR => \line_buffer.mem1_physical_WADDR_wire\,
            MASK => \line_buffer.mem1_physical_MASK_wire\,
            WDATA => \line_buffer.mem1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22688\,
            RE => \N__23370\,
            WCLKE => 'H',
            WCLK => \N__19325\,
            WE => \N__15719\
        );

    \line_buffer.mem15_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem15_physical_RDATA_wire\,
            RADDR => \line_buffer.mem15_physical_RADDR_wire\,
            WADDR => \line_buffer.mem15_physical_WADDR_wire\,
            MASK => \line_buffer.mem15_physical_MASK_wire\,
            WDATA => \line_buffer.mem15_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22622\,
            RE => \N__23260\,
            WCLKE => 'H',
            WCLK => \N__19348\,
            WE => \N__15720\
        );

    \line_buffer.mem27_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem27_physical_RDATA_wire\,
            RADDR => \line_buffer.mem27_physical_RADDR_wire\,
            WADDR => \line_buffer.mem27_physical_WADDR_wire\,
            MASK => \line_buffer.mem27_physical_MASK_wire\,
            WDATA => \line_buffer.mem27_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22640\,
            RE => \N__23373\,
            WCLKE => 'H',
            WCLK => \N__19343\,
            WE => \N__10113\
        );

    \line_buffer.mem4_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem4_physical_RDATA_wire\,
            RADDR => \line_buffer.mem4_physical_RADDR_wire\,
            WADDR => \line_buffer.mem4_physical_WADDR_wire\,
            MASK => \line_buffer.mem4_physical_MASK_wire\,
            WDATA => \line_buffer.mem4_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22488\,
            RE => \N__23282\,
            WCLKE => 'H',
            WCLK => \N__19355\,
            WE => \N__12658\
        );

    \line_buffer.mem16_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem16_physical_RDATA_wire\,
            RADDR => \line_buffer.mem16_physical_RADDR_wire\,
            WADDR => \line_buffer.mem16_physical_WADDR_wire\,
            MASK => \line_buffer.mem16_physical_MASK_wire\,
            WDATA => \line_buffer.mem16_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22583\,
            RE => \N__23192\,
            WCLKE => 'H',
            WCLK => \N__19350\,
            WE => \N__15721\
        );

    \line_buffer.mem30_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem30_physical_RDATA_wire\,
            RADDR => \line_buffer.mem30_physical_RADDR_wire\,
            WADDR => \line_buffer.mem30_physical_WADDR_wire\,
            MASK => \line_buffer.mem30_physical_MASK_wire\,
            WDATA => \line_buffer.mem30_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22579\,
            RE => \N__23326\,
            WCLKE => 'H',
            WCLK => \N__19351\,
            WE => \N__10262\
        );

    \line_buffer.mem7_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem7_physical_RDATA_wire\,
            RADDR => \line_buffer.mem7_physical_RADDR_wire\,
            WADDR => \line_buffer.mem7_physical_WADDR_wire\,
            MASK => \line_buffer.mem7_physical_MASK_wire\,
            WDATA => \line_buffer.mem7_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22020\,
            RE => \N__23228\,
            WCLKE => 'H',
            WCLK => \N__19364\,
            WE => \N__10181\
        );

    \line_buffer.mem20_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem20_physical_RDATA_wire\,
            RADDR => \line_buffer.mem20_physical_RADDR_wire\,
            WADDR => \line_buffer.mem20_physical_WADDR_wire\,
            MASK => \line_buffer.mem20_physical_MASK_wire\,
            WDATA => \line_buffer.mem20_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22205\,
            RE => \N__23190\,
            WCLKE => 'H',
            WCLK => \N__19363\,
            WE => \N__13475\
        );

    \line_buffer.mem13_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem13_physical_RDATA_wire\,
            RADDR => \line_buffer.mem13_physical_RADDR_wire\,
            WADDR => \line_buffer.mem13_physical_WADDR_wire\,
            MASK => \line_buffer.mem13_physical_MASK_wire\,
            WDATA => \line_buffer.mem13_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22654\,
            RE => \N__23310\,
            WCLKE => 'H',
            WCLK => \N__19344\,
            WE => \N__10225\
        );

    \line_buffer.mem19_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem19_physical_RDATA_wire\,
            RADDR => \line_buffer.mem19_physical_RADDR_wire\,
            WADDR => \line_buffer.mem19_physical_WADDR_wire\,
            MASK => \line_buffer.mem19_physical_MASK_wire\,
            WDATA => \line_buffer.mem19_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22515\,
            RE => \N__23117\,
            WCLKE => 'H',
            WCLK => \N__19359\,
            WE => \N__12605\
        );

    \line_buffer.mem23_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem23_physical_RDATA_wire\,
            RADDR => \line_buffer.mem23_physical_RADDR_wire\,
            WADDR => \line_buffer.mem23_physical_WADDR_wire\,
            MASK => \line_buffer.mem23_physical_MASK_wire\,
            WDATA => \line_buffer.mem23_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22690\,
            RE => \N__23395\,
            WCLKE => 'H',
            WCLK => \N__19323\,
            WE => \N__12657\
        );

    \line_buffer.mem0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem0_physical_RDATA_wire\,
            RADDR => \line_buffer.mem0_physical_RADDR_wire\,
            WADDR => \line_buffer.mem0_physical_WADDR_wire\,
            MASK => \line_buffer.mem0_physical_MASK_wire\,
            WDATA => \line_buffer.mem0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22689\,
            RE => \N__23371\,
            WCLKE => 'H',
            WCLK => \N__19321\,
            WE => \N__10234\
        );

    \line_buffer.mem26_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem26_physical_RDATA_wire\,
            RADDR => \line_buffer.mem26_physical_RADDR_wire\,
            WADDR => \line_buffer.mem26_physical_WADDR_wire\,
            MASK => \line_buffer.mem26_physical_MASK_wire\,
            WDATA => \line_buffer.mem26_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22668\,
            RE => \N__23386\,
            WCLKE => 'H',
            WCLK => \N__19337\,
            WE => \N__10112\
        );

    \line_buffer.mem3_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem3_physical_RDATA_wire\,
            RADDR => \line_buffer.mem3_physical_RADDR_wire\,
            WADDR => \line_buffer.mem3_physical_WADDR_wire\,
            MASK => \line_buffer.mem3_physical_MASK_wire\,
            WDATA => \line_buffer.mem3_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22538\,
            RE => \N__23352\,
            WCLKE => 'H',
            WCLK => \N__19349\,
            WE => \N__13474\
        );

    \line_buffer.mem17_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem17_physical_RDATA_wire\,
            RADDR => \line_buffer.mem17_physical_RADDR_wire\,
            WADDR => \line_buffer.mem17_physical_WADDR_wire\,
            MASK => \line_buffer.mem17_physical_MASK_wire\,
            WDATA => \line_buffer.mem17_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22582\,
            RE => \N__23191\,
            WCLKE => 'H',
            WCLK => \N__19352\,
            WE => \N__12598\
        );

    \line_buffer.mem31_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem31_physical_RDATA_wire\,
            RADDR => \line_buffer.mem31_physical_RADDR_wire\,
            WADDR => \line_buffer.mem31_physical_WADDR_wire\,
            MASK => \line_buffer.mem31_physical_MASK_wire\,
            WDATA => \line_buffer.mem31_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22436\,
            RE => \N__23325\,
            WCLKE => 'H',
            WCLK => \N__19353\,
            WE => \N__10269\
        );

    \line_buffer.mem9_physical\ : SB_RAM40_4K
    generic map (
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem9_physical_RDATA_wire\,
            RADDR => \line_buffer.mem9_physical_RADDR_wire\,
            WADDR => \line_buffer.mem9_physical_WADDR_wire\,
            MASK => \line_buffer.mem9_physical_MASK_wire\,
            WDATA => \line_buffer.mem9_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22037\,
            RE => \N__23343\,
            WCLKE => 'H',
            WCLK => \N__19368\,
            WE => \N__10189\
        );

    \line_buffer.mem29_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem29_physical_RDATA_wire\,
            RADDR => \line_buffer.mem29_physical_RADDR_wire\,
            WADDR => \line_buffer.mem29_physical_WADDR_wire\,
            MASK => \line_buffer.mem29_physical_MASK_wire\,
            WDATA => \line_buffer.mem29_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22675\,
            RE => \N__23353\,
            WCLKE => 'H',
            WCLK => \N__19347\,
            WE => \N__10253\
        );

    \line_buffer.mem6_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem6_physical_RDATA_wire\,
            RADDR => \line_buffer.mem6_physical_RADDR_wire\,
            WADDR => \line_buffer.mem6_physical_WADDR_wire\,
            MASK => \line_buffer.mem6_physical_MASK_wire\,
            WDATA => \line_buffer.mem6_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22408\,
            RE => \N__23227\,
            WCLKE => 'H',
            WCLK => \N__19362\,
            WE => \N__10273\
        );

    \line_buffer.mem10_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem10_physical_RDATA_wire\,
            RADDR => \line_buffer.mem10_physical_RADDR_wire\,
            WADDR => \line_buffer.mem10_physical_WADDR_wire\,
            MASK => \line_buffer.mem10_physical_MASK_wire\,
            WDATA => \line_buffer.mem10_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22677\,
            RE => \N__23345\,
            WCLKE => 'H',
            WCLK => \N__19331\,
            WE => \N__10180\
        );

    \line_buffer.mem22_physical\ : SB_RAM40_4K
    generic map (
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem22_physical_RDATA_wire\,
            RADDR => \line_buffer.mem22_physical_RADDR_wire\,
            WADDR => \line_buffer.mem22_physical_WADDR_wire\,
            MASK => \line_buffer.mem22_physical_MASK_wire\,
            WDATA => \line_buffer.mem22_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22239\,
            RE => \N__23139\,
            WCLKE => 'H',
            WCLK => \N__19367\,
            WE => \N__13485\
        );

    \line_buffer.mem25_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem25_physical_RDATA_wire\,
            RADDR => \line_buffer.mem25_physical_RADDR_wire\,
            WADDR => \line_buffer.mem25_physical_WADDR_wire\,
            MASK => \line_buffer.mem25_physical_MASK_wire\,
            WDATA => \line_buffer.mem25_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22684\,
            RE => \N__23387\,
            WCLKE => 'H',
            WCLK => \N__19332\,
            WE => \N__12646\
        );

    \line_buffer.mem8_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem8_physical_RDATA_wire\,
            RADDR => \line_buffer.mem8_physical_RADDR_wire\,
            WADDR => \line_buffer.mem8_physical_WADDR_wire\,
            MASK => \line_buffer.mem8_physical_MASK_wire\,
            WDATA => \line_buffer.mem8_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22225\,
            RE => \N__23299\,
            WCLKE => 'H',
            WCLK => \N__19366\,
            WE => \N__10188\
        );

    \line_buffer.mem28_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \line_buffer.mem28_physical_RDATA_wire\,
            RADDR => \line_buffer.mem28_physical_RADDR_wire\,
            WADDR => \line_buffer.mem28_physical_WADDR_wire\,
            MASK => \line_buffer.mem28_physical_MASK_wire\,
            WDATA => \line_buffer.mem28_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22600\,
            RE => \N__23372\,
            WCLKE => 'H',
            WCLK => \N__19345\,
            WE => \N__10105\
        );

    \DEBUG_c_1_pad_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__24374\,
            GLOBALBUFFEROUTPUT => \DEBUG_c_1_c\
        );

    \DEBUG_c_1_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24376\,
            DIN => \N__24375\,
            DOUT => \N__24374\,
            PACKAGEPIN => \TVP_CLK_wire\
        );

    \DEBUG_c_1_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24376\,
            PADOUT => \N__24375\,
            PADIN => \N__24374\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24365\,
            DIN => \N__24364\,
            DOUT => \N__24363\,
            PACKAGEPIN => \ADV_CLK_wire\
        );

    \ADV_CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24365\,
            PADOUT => \N__24364\,
            PADIN => \N__24363\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__22536\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24356\,
            DIN => \N__24355\,
            DOUT => \N__24354\,
            PACKAGEPIN => DEBUG(3)
        );

    \DEBUG_pad_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24356\,
            PADOUT => \N__24355\,
            PADIN => \N__24354\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__15769\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_VIDEO_pad_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24347\,
            DIN => \N__24346\,
            DOUT => \N__24345\,
            PACKAGEPIN => \TVP_VIDEO_wire\(2)
        );

    \TVP_VIDEO_pad_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24347\,
            PADOUT => \N__24346\,
            PADIN => \N__24345\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_VIDEO_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24338\,
            DIN => \N__24337\,
            DOUT => \N__24336\,
            PACKAGEPIN => \ADV_G_wire\(5)
        );

    \ADV_G_pad_5_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24338\,
            PADOUT => \N__24337\,
            PADIN => \N__24336\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__14304\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24329\,
            DIN => \N__24328\,
            DOUT => \N__24327\,
            PACKAGEPIN => \ADV_R_wire\(3)
        );

    \ADV_R_pad_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24329\,
            PADOUT => \N__24328\,
            PADIN => \N__24327\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__14415\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24320\,
            DIN => \N__24319\,
            DOUT => \N__24318\,
            PACKAGEPIN => \ADV_G_wire\(1)
        );

    \ADV_G_pad_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24320\,
            PADOUT => \N__24319\,
            PADIN => \N__24318\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__14524\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24311\,
            DIN => \N__24310\,
            DOUT => \N__24309\,
            PACKAGEPIN => \ADV_R_wire\(0)
        );

    \ADV_R_pad_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24311\,
            PADOUT => \N__24310\,
            PADIN => \N__24309\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10047\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24302\,
            DIN => \N__24301\,
            DOUT => \N__24300\,
            PACKAGEPIN => DEBUG(2)
        );

    \DEBUG_pad_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24302\,
            PADOUT => \N__24301\,
            PADIN => \N__24300\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__22873\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_VIDEO_pad_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24293\,
            DIN => \N__24292\,
            DOUT => \N__24291\,
            PACKAGEPIN => \TVP_VIDEO_wire\(3)
        );

    \TVP_VIDEO_pad_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24293\,
            PADOUT => \N__24292\,
            PADIN => \N__24291\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_VIDEO_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24284\,
            DIN => \N__24283\,
            DOUT => \N__24282\,
            PACKAGEPIN => \ADV_G_wire\(4)
        );

    \ADV_G_pad_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24284\,
            PADOUT => \N__24283\,
            PADIN => \N__24282\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__14351\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24275\,
            DIN => \N__24274\,
            DOUT => \N__24273\,
            PACKAGEPIN => \ADV_R_wire\(5)
        );

    \ADV_R_pad_5_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24275\,
            PADOUT => \N__24274\,
            PADIN => \N__24273\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__14300\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_VIDEO_pad_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24266\,
            DIN => \N__24265\,
            DOUT => \N__24264\,
            PACKAGEPIN => \TVP_VIDEO_wire\(9)
        );

    \TVP_VIDEO_pad_9_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24266\,
            PADOUT => \N__24265\,
            PADIN => \N__24264\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_VIDEO_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24257\,
            DIN => \N__24256\,
            DOUT => \N__24255\,
            PACKAGEPIN => DEBUG(1)
        );

    \DEBUG_pad_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24257\,
            PADOUT => \N__24256\,
            PADIN => \N__24255\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__19222\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24248\,
            DIN => \N__24247\,
            DOUT => \N__24246\,
            PACKAGEPIN => \ADV_B_wire\(1)
        );

    \ADV_B_pad_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24248\,
            PADOUT => \N__24247\,
            PADIN => \N__24246\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__14513\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_SYNC_N_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24239\,
            DIN => \N__24238\,
            DOUT => \N__24237\,
            PACKAGEPIN => \ADV_SYNC_N_wire\
        );

    \ADV_SYNC_N_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24239\,
            PADOUT => \N__24238\,
            PADIN => \N__24237\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24230\,
            DIN => \N__24229\,
            DOUT => \N__24228\,
            PACKAGEPIN => \ADV_B_wire\(6)
        );

    \ADV_B_pad_6_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24230\,
            PADOUT => \N__24229\,
            PADIN => \N__24228\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__14245\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24221\,
            DIN => \N__24220\,
            DOUT => \N__24219\,
            PACKAGEPIN => DEBUG(6)
        );

    \DEBUG_pad_6_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24221\,
            PADOUT => \N__24220\,
            PADIN => \N__24219\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9676\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_VIDEO_pad_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24212\,
            DIN => \N__24211\,
            DOUT => \N__24210\,
            PACKAGEPIN => \TVP_VIDEO_wire\(7)
        );

    \TVP_VIDEO_pad_7_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24212\,
            PADOUT => \N__24211\,
            PADIN => \N__24210\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_VIDEO_c_7\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24203\,
            DIN => \N__24202\,
            DOUT => \N__24201\,
            PACKAGEPIN => \ADV_G_wire\(0)
        );

    \ADV_G_pad_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24203\,
            PADOUT => \N__24202\,
            PADIN => \N__24201\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10054\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24194\,
            DIN => \N__24193\,
            DOUT => \N__24192\,
            PACKAGEPIN => \ADV_R_wire\(1)
        );

    \ADV_R_pad_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24194\,
            PADOUT => \N__24193\,
            PADIN => \N__24192\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__14520\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24185\,
            DIN => \N__24184\,
            DOUT => \N__24183\,
            PACKAGEPIN => DEBUG(5)
        );

    \DEBUG_pad_5_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24185\,
            PADOUT => \N__24184\,
            PADIN => \N__24183\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__15856\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_HSYNC_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24176\,
            DIN => \N__24175\,
            DOUT => \N__24174\,
            PACKAGEPIN => \TVP_HSYNC_wire\
        );

    \TVP_HSYNC_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24176\,
            PADOUT => \N__24175\,
            PADIN => \N__24174\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_HSYNC_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24167\,
            DIN => \N__24166\,
            DOUT => \N__24165\,
            PACKAGEPIN => \ADV_G_wire\(7)
        );

    \ADV_G_pad_7_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24167\,
            PADOUT => \N__24166\,
            PADIN => \N__24165\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__14171\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24158\,
            DIN => \N__24157\,
            DOUT => \N__24156\,
            PACKAGEPIN => \ADV_R_wire\(6)
        );

    \ADV_R_pad_6_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24158\,
            PADOUT => \N__24157\,
            PADIN => \N__24156\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__14243\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_VSYNC_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24149\,
            DIN => \N__24148\,
            DOUT => \N__24147\,
            PACKAGEPIN => \TVP_VSYNC_wire\
        );

    \TVP_VSYNC_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24149\,
            PADOUT => \N__24148\,
            PADIN => \N__24147\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_VSYNC_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_BLANK_N_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24140\,
            DIN => \N__24139\,
            DOUT => \N__24138\,
            PACKAGEPIN => \ADV_BLANK_N_wire\
        );

    \ADV_BLANK_N_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24140\,
            PADOUT => \N__24139\,
            PADIN => \N__24138\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__23323\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24131\,
            DIN => \N__24130\,
            DOUT => \N__24129\,
            PACKAGEPIN => DEBUG(0)
        );

    \DEBUG_pad_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24131\,
            PADOUT => \N__24130\,
            PADIN => \N__24129\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10075\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24122\,
            DIN => \N__24121\,
            DOUT => \N__24120\,
            PACKAGEPIN => \ADV_B_wire\(2)
        );

    \ADV_B_pad_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24122\,
            PADOUT => \N__24121\,
            PADIN => \N__24120\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__14463\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24113\,
            DIN => \N__24112\,
            DOUT => \N__24111\,
            PACKAGEPIN => \ADV_B_wire\(7)
        );

    \ADV_B_pad_7_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24113\,
            PADOUT => \N__24112\,
            PADIN => \N__24111\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__14182\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LED_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24104\,
            DIN => \N__24103\,
            DOUT => \N__24102\,
            PACKAGEPIN => \LED_wire\
        );

    \LED_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24104\,
            PADOUT => \N__24103\,
            PADIN => \N__24102\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__17359\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_VIDEO_pad_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24095\,
            DIN => \N__24094\,
            DOUT => \N__24093\,
            PACKAGEPIN => \TVP_VIDEO_wire\(4)
        );

    \TVP_VIDEO_pad_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24095\,
            PADOUT => \N__24094\,
            PADIN => \N__24093\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_VIDEO_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24086\,
            DIN => \N__24085\,
            DOUT => \N__24084\,
            PACKAGEPIN => \ADV_G_wire\(3)
        );

    \ADV_G_pad_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24086\,
            PADOUT => \N__24085\,
            PADIN => \N__24084\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__14411\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_HSYNC_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24077\,
            DIN => \N__24076\,
            DOUT => \N__24075\,
            PACKAGEPIN => \ADV_HSYNC_wire\
        );

    \ADV_HSYNC_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24077\,
            PADOUT => \N__24076\,
            PADIN => \N__24075\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__16729\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24068\,
            DIN => \N__24067\,
            DOUT => \N__24066\,
            PACKAGEPIN => \ADV_R_wire\(2)
        );

    \ADV_R_pad_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24068\,
            PADOUT => \N__24067\,
            PADIN => \N__24066\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__14462\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24059\,
            DIN => \N__24058\,
            DOUT => \N__24057\,
            PACKAGEPIN => \ADV_B_wire\(4)
        );

    \ADV_B_pad_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24059\,
            PADOUT => \N__24058\,
            PADIN => \N__24057\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__14359\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24050\,
            DIN => \N__24049\,
            DOUT => \N__24048\,
            PACKAGEPIN => DEBUG(4)
        );

    \DEBUG_pad_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24050\,
            PADOUT => \N__24049\,
            PADIN => \N__24048\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10657\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24041\,
            DIN => \N__24040\,
            DOUT => \N__24039\,
            PACKAGEPIN => \ADV_G_wire\(6)
        );

    \ADV_G_pad_6_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24041\,
            PADOUT => \N__24040\,
            PADIN => \N__24039\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__14244\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24032\,
            DIN => \N__24031\,
            DOUT => \N__24030\,
            PACKAGEPIN => \ADV_R_wire\(7)
        );

    \ADV_R_pad_7_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24032\,
            PADOUT => \N__24031\,
            PADIN => \N__24030\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__14181\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24023\,
            DIN => \N__24022\,
            DOUT => \N__24021\,
            PACKAGEPIN => \ADV_B_wire\(3)
        );

    \ADV_B_pad_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24023\,
            PADOUT => \N__24022\,
            PADIN => \N__24021\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__14416\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24014\,
            DIN => \N__24013\,
            DOUT => \N__24012\,
            PACKAGEPIN => \ADV_R_wire\(4)
        );

    \ADV_R_pad_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24014\,
            PADOUT => \N__24013\,
            PADIN => \N__24012\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__14352\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_VIDEO_pad_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24005\,
            DIN => \N__24004\,
            DOUT => \N__24003\,
            PACKAGEPIN => \TVP_VIDEO_wire\(8)
        );

    \TVP_VIDEO_pad_8_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24005\,
            PADOUT => \N__24004\,
            PADIN => \N__24003\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_VIDEO_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23996\,
            DIN => \N__23995\,
            DOUT => \N__23994\,
            PACKAGEPIN => \ADV_B_wire\(0)
        );

    \ADV_B_pad_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23996\,
            PADOUT => \N__23995\,
            PADIN => \N__23994\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10040\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_VIDEO_pad_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__23987\,
            DIN => \N__23986\,
            DOUT => \N__23985\,
            PACKAGEPIN => \TVP_VIDEO_wire\(5)
        );

    \TVP_VIDEO_pad_5_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23987\,
            PADOUT => \N__23986\,
            PADIN => \N__23985\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_VIDEO_c_5\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23978\,
            DIN => \N__23977\,
            DOUT => \N__23976\,
            PACKAGEPIN => \ADV_G_wire\(2)
        );

    \ADV_G_pad_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23978\,
            PADOUT => \N__23977\,
            PADIN => \N__23976\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__14464\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_VSYNC_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23969\,
            DIN => \N__23968\,
            DOUT => \N__23967\,
            PACKAGEPIN => \ADV_VSYNC_wire\
        );

    \ADV_VSYNC_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23969\,
            PADOUT => \N__23968\,
            PADIN => \N__23967\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__21171\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__23960\,
            DIN => \N__23959\,
            DOUT => \N__23958\,
            PACKAGEPIN => \ADV_B_wire\(5)
        );

    \ADV_B_pad_5_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23960\,
            PADOUT => \N__23959\,
            PADIN => \N__23958\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__14305\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__23951\,
            DIN => \N__23950\,
            DOUT => \N__23949\,
            PACKAGEPIN => DEBUG(7)
        );

    \DEBUG_pad_7_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23951\,
            PADOUT => \N__23950\,
            PADIN => \N__23949\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__23385\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_VIDEO_pad_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__23942\,
            DIN => \N__23941\,
            DOUT => \N__23940\,
            PACKAGEPIN => \TVP_VIDEO_wire\(6)
        );

    \TVP_VIDEO_pad_6_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__23942\,
            PADOUT => \N__23941\,
            PADIN => \N__23940\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_VIDEO_c_6\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__5782\ : InMux
    port map (
            O => \N__23923\,
            I => \N__23920\
        );

    \I__5781\ : LocalMux
    port map (
            O => \N__23920\,
            I => \N__23917\
        );

    \I__5780\ : Span12Mux_h
    port map (
            O => \N__23917\,
            I => \N__23914\
        );

    \I__5779\ : Span12Mux_v
    port map (
            O => \N__23914\,
            I => \N__23911\
        );

    \I__5778\ : Odrv12
    port map (
            O => \N__23911\,
            I => \line_buffer.n548\
        );

    \I__5777\ : InMux
    port map (
            O => \N__23908\,
            I => \N__23905\
        );

    \I__5776\ : LocalMux
    port map (
            O => \N__23905\,
            I => \N__23902\
        );

    \I__5775\ : Span4Mux_h
    port map (
            O => \N__23902\,
            I => \N__23899\
        );

    \I__5774\ : Span4Mux_h
    port map (
            O => \N__23899\,
            I => \N__23896\
        );

    \I__5773\ : Odrv4
    port map (
            O => \N__23896\,
            I => \line_buffer.n556\
        );

    \I__5772\ : CascadeMux
    port map (
            O => \N__23893\,
            I => \N__23890\
        );

    \I__5771\ : InMux
    port map (
            O => \N__23890\,
            I => \N__23887\
        );

    \I__5770\ : LocalMux
    port map (
            O => \N__23887\,
            I => \N__23884\
        );

    \I__5769\ : Odrv12
    port map (
            O => \N__23884\,
            I => \line_buffer.n4077\
        );

    \I__5768\ : InMux
    port map (
            O => \N__23881\,
            I => \N__23878\
        );

    \I__5767\ : LocalMux
    port map (
            O => \N__23878\,
            I => \N__23875\
        );

    \I__5766\ : Span4Mux_v
    port map (
            O => \N__23875\,
            I => \N__23872\
        );

    \I__5765\ : Span4Mux_h
    port map (
            O => \N__23872\,
            I => \N__23869\
        );

    \I__5764\ : Sp12to4
    port map (
            O => \N__23869\,
            I => \N__23866\
        );

    \I__5763\ : Odrv12
    port map (
            O => \N__23866\,
            I => \line_buffer.n674\
        );

    \I__5762\ : InMux
    port map (
            O => \N__23863\,
            I => \N__23860\
        );

    \I__5761\ : LocalMux
    port map (
            O => \N__23860\,
            I => \N__23856\
        );

    \I__5760\ : InMux
    port map (
            O => \N__23859\,
            I => \N__23852\
        );

    \I__5759\ : Span4Mux_v
    port map (
            O => \N__23856\,
            I => \N__23833\
        );

    \I__5758\ : InMux
    port map (
            O => \N__23855\,
            I => \N__23830\
        );

    \I__5757\ : LocalMux
    port map (
            O => \N__23852\,
            I => \N__23825\
        );

    \I__5756\ : InMux
    port map (
            O => \N__23851\,
            I => \N__23822\
        );

    \I__5755\ : InMux
    port map (
            O => \N__23850\,
            I => \N__23819\
        );

    \I__5754\ : InMux
    port map (
            O => \N__23849\,
            I => \N__23813\
        );

    \I__5753\ : InMux
    port map (
            O => \N__23848\,
            I => \N__23813\
        );

    \I__5752\ : InMux
    port map (
            O => \N__23847\,
            I => \N__23808\
        );

    \I__5751\ : InMux
    port map (
            O => \N__23846\,
            I => \N__23808\
        );

    \I__5750\ : InMux
    port map (
            O => \N__23845\,
            I => \N__23803\
        );

    \I__5749\ : InMux
    port map (
            O => \N__23844\,
            I => \N__23800\
        );

    \I__5748\ : InMux
    port map (
            O => \N__23843\,
            I => \N__23795\
        );

    \I__5747\ : InMux
    port map (
            O => \N__23842\,
            I => \N__23795\
        );

    \I__5746\ : InMux
    port map (
            O => \N__23841\,
            I => \N__23790\
        );

    \I__5745\ : InMux
    port map (
            O => \N__23840\,
            I => \N__23790\
        );

    \I__5744\ : InMux
    port map (
            O => \N__23839\,
            I => \N__23783\
        );

    \I__5743\ : InMux
    port map (
            O => \N__23838\,
            I => \N__23783\
        );

    \I__5742\ : InMux
    port map (
            O => \N__23837\,
            I => \N__23783\
        );

    \I__5741\ : InMux
    port map (
            O => \N__23836\,
            I => \N__23780\
        );

    \I__5740\ : Span4Mux_h
    port map (
            O => \N__23833\,
            I => \N__23775\
        );

    \I__5739\ : LocalMux
    port map (
            O => \N__23830\,
            I => \N__23775\
        );

    \I__5738\ : InMux
    port map (
            O => \N__23829\,
            I => \N__23772\
        );

    \I__5737\ : InMux
    port map (
            O => \N__23828\,
            I => \N__23769\
        );

    \I__5736\ : Span4Mux_v
    port map (
            O => \N__23825\,
            I => \N__23762\
        );

    \I__5735\ : LocalMux
    port map (
            O => \N__23822\,
            I => \N__23762\
        );

    \I__5734\ : LocalMux
    port map (
            O => \N__23819\,
            I => \N__23762\
        );

    \I__5733\ : InMux
    port map (
            O => \N__23818\,
            I => \N__23759\
        );

    \I__5732\ : LocalMux
    port map (
            O => \N__23813\,
            I => \N__23756\
        );

    \I__5731\ : LocalMux
    port map (
            O => \N__23808\,
            I => \N__23753\
        );

    \I__5730\ : InMux
    port map (
            O => \N__23807\,
            I => \N__23750\
        );

    \I__5729\ : CascadeMux
    port map (
            O => \N__23806\,
            I => \N__23747\
        );

    \I__5728\ : LocalMux
    port map (
            O => \N__23803\,
            I => \N__23742\
        );

    \I__5727\ : LocalMux
    port map (
            O => \N__23800\,
            I => \N__23742\
        );

    \I__5726\ : LocalMux
    port map (
            O => \N__23795\,
            I => \N__23736\
        );

    \I__5725\ : LocalMux
    port map (
            O => \N__23790\,
            I => \N__23736\
        );

    \I__5724\ : LocalMux
    port map (
            O => \N__23783\,
            I => \N__23731\
        );

    \I__5723\ : LocalMux
    port map (
            O => \N__23780\,
            I => \N__23731\
        );

    \I__5722\ : Span4Mux_h
    port map (
            O => \N__23775\,
            I => \N__23720\
        );

    \I__5721\ : LocalMux
    port map (
            O => \N__23772\,
            I => \N__23720\
        );

    \I__5720\ : LocalMux
    port map (
            O => \N__23769\,
            I => \N__23720\
        );

    \I__5719\ : Span4Mux_v
    port map (
            O => \N__23762\,
            I => \N__23720\
        );

    \I__5718\ : LocalMux
    port map (
            O => \N__23759\,
            I => \N__23720\
        );

    \I__5717\ : Span4Mux_h
    port map (
            O => \N__23756\,
            I => \N__23715\
        );

    \I__5716\ : Span4Mux_h
    port map (
            O => \N__23753\,
            I => \N__23715\
        );

    \I__5715\ : LocalMux
    port map (
            O => \N__23750\,
            I => \N__23712\
        );

    \I__5714\ : InMux
    port map (
            O => \N__23747\,
            I => \N__23709\
        );

    \I__5713\ : Span4Mux_h
    port map (
            O => \N__23742\,
            I => \N__23706\
        );

    \I__5712\ : InMux
    port map (
            O => \N__23741\,
            I => \N__23703\
        );

    \I__5711\ : Span4Mux_h
    port map (
            O => \N__23736\,
            I => \N__23700\
        );

    \I__5710\ : Span12Mux_h
    port map (
            O => \N__23731\,
            I => \N__23697\
        );

    \I__5709\ : Span4Mux_h
    port map (
            O => \N__23720\,
            I => \N__23694\
        );

    \I__5708\ : Span4Mux_v
    port map (
            O => \N__23715\,
            I => \N__23685\
        );

    \I__5707\ : Span4Mux_h
    port map (
            O => \N__23712\,
            I => \N__23685\
        );

    \I__5706\ : LocalMux
    port map (
            O => \N__23709\,
            I => \N__23685\
        );

    \I__5705\ : Span4Mux_h
    port map (
            O => \N__23706\,
            I => \N__23685\
        );

    \I__5704\ : LocalMux
    port map (
            O => \N__23703\,
            I => \TX_ADDR_12\
        );

    \I__5703\ : Odrv4
    port map (
            O => \N__23700\,
            I => \TX_ADDR_12\
        );

    \I__5702\ : Odrv12
    port map (
            O => \N__23697\,
            I => \TX_ADDR_12\
        );

    \I__5701\ : Odrv4
    port map (
            O => \N__23694\,
            I => \TX_ADDR_12\
        );

    \I__5700\ : Odrv4
    port map (
            O => \N__23685\,
            I => \TX_ADDR_12\
        );

    \I__5699\ : CascadeMux
    port map (
            O => \N__23674\,
            I => \N__23671\
        );

    \I__5698\ : InMux
    port map (
            O => \N__23671\,
            I => \N__23668\
        );

    \I__5697\ : LocalMux
    port map (
            O => \N__23668\,
            I => \N__23665\
        );

    \I__5696\ : Span12Mux_h
    port map (
            O => \N__23665\,
            I => \N__23662\
        );

    \I__5695\ : Odrv12
    port map (
            O => \N__23662\,
            I => \line_buffer.n682\
        );

    \I__5694\ : InMux
    port map (
            O => \N__23659\,
            I => \N__23656\
        );

    \I__5693\ : LocalMux
    port map (
            O => \N__23656\,
            I => \line_buffer.n4158\
        );

    \I__5692\ : InMux
    port map (
            O => \N__23653\,
            I => \N__23650\
        );

    \I__5691\ : LocalMux
    port map (
            O => \N__23650\,
            I => \N__23647\
        );

    \I__5690\ : Span4Mux_v
    port map (
            O => \N__23647\,
            I => \N__23644\
        );

    \I__5689\ : Sp12to4
    port map (
            O => \N__23644\,
            I => \N__23641\
        );

    \I__5688\ : Span12Mux_h
    port map (
            O => \N__23641\,
            I => \N__23638\
        );

    \I__5687\ : Odrv12
    port map (
            O => \N__23638\,
            I => \line_buffer.n685\
        );

    \I__5686\ : InMux
    port map (
            O => \N__23635\,
            I => \N__23632\
        );

    \I__5685\ : LocalMux
    port map (
            O => \N__23632\,
            I => \N__23629\
        );

    \I__5684\ : Span4Mux_v
    port map (
            O => \N__23629\,
            I => \N__23626\
        );

    \I__5683\ : Span4Mux_v
    port map (
            O => \N__23626\,
            I => \N__23623\
        );

    \I__5682\ : Span4Mux_v
    port map (
            O => \N__23623\,
            I => \N__23620\
        );

    \I__5681\ : Span4Mux_h
    port map (
            O => \N__23620\,
            I => \N__23617\
        );

    \I__5680\ : Odrv4
    port map (
            O => \N__23617\,
            I => \line_buffer.n677\
        );

    \I__5679\ : InMux
    port map (
            O => \N__23614\,
            I => \N__23608\
        );

    \I__5678\ : CascadeMux
    port map (
            O => \N__23613\,
            I => \N__23605\
        );

    \I__5677\ : InMux
    port map (
            O => \N__23612\,
            I => \N__23595\
        );

    \I__5676\ : InMux
    port map (
            O => \N__23611\,
            I => \N__23592\
        );

    \I__5675\ : LocalMux
    port map (
            O => \N__23608\,
            I => \N__23587\
        );

    \I__5674\ : InMux
    port map (
            O => \N__23605\,
            I => \N__23583\
        );

    \I__5673\ : InMux
    port map (
            O => \N__23604\,
            I => \N__23578\
        );

    \I__5672\ : InMux
    port map (
            O => \N__23603\,
            I => \N__23578\
        );

    \I__5671\ : InMux
    port map (
            O => \N__23602\,
            I => \N__23573\
        );

    \I__5670\ : InMux
    port map (
            O => \N__23601\,
            I => \N__23570\
        );

    \I__5669\ : InMux
    port map (
            O => \N__23600\,
            I => \N__23563\
        );

    \I__5668\ : InMux
    port map (
            O => \N__23599\,
            I => \N__23563\
        );

    \I__5667\ : InMux
    port map (
            O => \N__23598\,
            I => \N__23563\
        );

    \I__5666\ : LocalMux
    port map (
            O => \N__23595\,
            I => \N__23560\
        );

    \I__5665\ : LocalMux
    port map (
            O => \N__23592\,
            I => \N__23557\
        );

    \I__5664\ : InMux
    port map (
            O => \N__23591\,
            I => \N__23554\
        );

    \I__5663\ : InMux
    port map (
            O => \N__23590\,
            I => \N__23550\
        );

    \I__5662\ : Span4Mux_v
    port map (
            O => \N__23587\,
            I => \N__23547\
        );

    \I__5661\ : InMux
    port map (
            O => \N__23586\,
            I => \N__23544\
        );

    \I__5660\ : LocalMux
    port map (
            O => \N__23583\,
            I => \N__23540\
        );

    \I__5659\ : LocalMux
    port map (
            O => \N__23578\,
            I => \N__23537\
        );

    \I__5658\ : InMux
    port map (
            O => \N__23577\,
            I => \N__23532\
        );

    \I__5657\ : InMux
    port map (
            O => \N__23576\,
            I => \N__23529\
        );

    \I__5656\ : LocalMux
    port map (
            O => \N__23573\,
            I => \N__23522\
        );

    \I__5655\ : LocalMux
    port map (
            O => \N__23570\,
            I => \N__23522\
        );

    \I__5654\ : LocalMux
    port map (
            O => \N__23563\,
            I => \N__23522\
        );

    \I__5653\ : Span4Mux_h
    port map (
            O => \N__23560\,
            I => \N__23519\
        );

    \I__5652\ : Span4Mux_h
    port map (
            O => \N__23557\,
            I => \N__23513\
        );

    \I__5651\ : LocalMux
    port map (
            O => \N__23554\,
            I => \N__23513\
        );

    \I__5650\ : InMux
    port map (
            O => \N__23553\,
            I => \N__23510\
        );

    \I__5649\ : LocalMux
    port map (
            O => \N__23550\,
            I => \N__23503\
        );

    \I__5648\ : Span4Mux_v
    port map (
            O => \N__23547\,
            I => \N__23503\
        );

    \I__5647\ : LocalMux
    port map (
            O => \N__23544\,
            I => \N__23503\
        );

    \I__5646\ : InMux
    port map (
            O => \N__23543\,
            I => \N__23500\
        );

    \I__5645\ : Span4Mux_h
    port map (
            O => \N__23540\,
            I => \N__23497\
        );

    \I__5644\ : Span4Mux_h
    port map (
            O => \N__23537\,
            I => \N__23494\
        );

    \I__5643\ : InMux
    port map (
            O => \N__23536\,
            I => \N__23489\
        );

    \I__5642\ : InMux
    port map (
            O => \N__23535\,
            I => \N__23486\
        );

    \I__5641\ : LocalMux
    port map (
            O => \N__23532\,
            I => \N__23482\
        );

    \I__5640\ : LocalMux
    port map (
            O => \N__23529\,
            I => \N__23479\
        );

    \I__5639\ : Span4Mux_v
    port map (
            O => \N__23522\,
            I => \N__23474\
        );

    \I__5638\ : Span4Mux_v
    port map (
            O => \N__23519\,
            I => \N__23474\
        );

    \I__5637\ : InMux
    port map (
            O => \N__23518\,
            I => \N__23471\
        );

    \I__5636\ : Span4Mux_v
    port map (
            O => \N__23513\,
            I => \N__23468\
        );

    \I__5635\ : LocalMux
    port map (
            O => \N__23510\,
            I => \N__23465\
        );

    \I__5634\ : Span4Mux_v
    port map (
            O => \N__23503\,
            I => \N__23462\
        );

    \I__5633\ : LocalMux
    port map (
            O => \N__23500\,
            I => \N__23459\
        );

    \I__5632\ : Span4Mux_v
    port map (
            O => \N__23497\,
            I => \N__23454\
        );

    \I__5631\ : Span4Mux_v
    port map (
            O => \N__23494\,
            I => \N__23454\
        );

    \I__5630\ : InMux
    port map (
            O => \N__23493\,
            I => \N__23449\
        );

    \I__5629\ : InMux
    port map (
            O => \N__23492\,
            I => \N__23449\
        );

    \I__5628\ : LocalMux
    port map (
            O => \N__23489\,
            I => \N__23444\
        );

    \I__5627\ : LocalMux
    port map (
            O => \N__23486\,
            I => \N__23444\
        );

    \I__5626\ : InMux
    port map (
            O => \N__23485\,
            I => \N__23441\
        );

    \I__5625\ : Span12Mux_h
    port map (
            O => \N__23482\,
            I => \N__23438\
        );

    \I__5624\ : Span4Mux_h
    port map (
            O => \N__23479\,
            I => \N__23431\
        );

    \I__5623\ : Span4Mux_h
    port map (
            O => \N__23474\,
            I => \N__23431\
        );

    \I__5622\ : LocalMux
    port map (
            O => \N__23471\,
            I => \N__23431\
        );

    \I__5621\ : Span4Mux_v
    port map (
            O => \N__23468\,
            I => \N__23422\
        );

    \I__5620\ : Span4Mux_v
    port map (
            O => \N__23465\,
            I => \N__23422\
        );

    \I__5619\ : Span4Mux_h
    port map (
            O => \N__23462\,
            I => \N__23422\
        );

    \I__5618\ : Span4Mux_h
    port map (
            O => \N__23459\,
            I => \N__23422\
        );

    \I__5617\ : Span4Mux_h
    port map (
            O => \N__23454\,
            I => \N__23419\
        );

    \I__5616\ : LocalMux
    port map (
            O => \N__23449\,
            I => \N__23414\
        );

    \I__5615\ : Span12Mux_h
    port map (
            O => \N__23444\,
            I => \N__23414\
        );

    \I__5614\ : LocalMux
    port map (
            O => \N__23441\,
            I => \TX_ADDR_11\
        );

    \I__5613\ : Odrv12
    port map (
            O => \N__23438\,
            I => \TX_ADDR_11\
        );

    \I__5612\ : Odrv4
    port map (
            O => \N__23431\,
            I => \TX_ADDR_11\
        );

    \I__5611\ : Odrv4
    port map (
            O => \N__23422\,
            I => \TX_ADDR_11\
        );

    \I__5610\ : Odrv4
    port map (
            O => \N__23419\,
            I => \TX_ADDR_11\
        );

    \I__5609\ : Odrv12
    port map (
            O => \N__23414\,
            I => \TX_ADDR_11\
        );

    \I__5608\ : InMux
    port map (
            O => \N__23401\,
            I => \N__23398\
        );

    \I__5607\ : LocalMux
    port map (
            O => \N__23398\,
            I => \line_buffer.n4063\
        );

    \I__5606\ : SRMux
    port map (
            O => \N__23395\,
            I => \N__23391\
        );

    \I__5605\ : SRMux
    port map (
            O => \N__23394\,
            I => \N__23388\
        );

    \I__5604\ : LocalMux
    port map (
            O => \N__23391\,
            I => \N__23380\
        );

    \I__5603\ : LocalMux
    port map (
            O => \N__23388\,
            I => \N__23380\
        );

    \I__5602\ : SRMux
    port map (
            O => \N__23387\,
            I => \N__23377\
        );

    \I__5601\ : SRMux
    port map (
            O => \N__23386\,
            I => \N__23374\
        );

    \I__5600\ : IoInMux
    port map (
            O => \N__23385\,
            I => \N__23367\
        );

    \I__5599\ : Span4Mux_s3_v
    port map (
            O => \N__23380\,
            I => \N__23360\
        );

    \I__5598\ : LocalMux
    port map (
            O => \N__23377\,
            I => \N__23360\
        );

    \I__5597\ : LocalMux
    port map (
            O => \N__23374\,
            I => \N__23360\
        );

    \I__5596\ : SRMux
    port map (
            O => \N__23373\,
            I => \N__23357\
        );

    \I__5595\ : SRMux
    port map (
            O => \N__23372\,
            I => \N__23354\
        );

    \I__5594\ : SRMux
    port map (
            O => \N__23371\,
            I => \N__23349\
        );

    \I__5593\ : SRMux
    port map (
            O => \N__23370\,
            I => \N__23346\
        );

    \I__5592\ : LocalMux
    port map (
            O => \N__23367\,
            I => \N__23340\
        );

    \I__5591\ : Span4Mux_v
    port map (
            O => \N__23360\,
            I => \N__23333\
        );

    \I__5590\ : LocalMux
    port map (
            O => \N__23357\,
            I => \N__23333\
        );

    \I__5589\ : LocalMux
    port map (
            O => \N__23354\,
            I => \N__23333\
        );

    \I__5588\ : SRMux
    port map (
            O => \N__23353\,
            I => \N__23330\
        );

    \I__5587\ : SRMux
    port map (
            O => \N__23352\,
            I => \N__23327\
        );

    \I__5586\ : LocalMux
    port map (
            O => \N__23349\,
            I => \N__23318\
        );

    \I__5585\ : LocalMux
    port map (
            O => \N__23346\,
            I => \N__23318\
        );

    \I__5584\ : SRMux
    port map (
            O => \N__23345\,
            I => \N__23315\
        );

    \I__5583\ : SRMux
    port map (
            O => \N__23344\,
            I => \N__23312\
        );

    \I__5582\ : SRMux
    port map (
            O => \N__23343\,
            I => \N__23300\
        );

    \I__5581\ : Span4Mux_s0_h
    port map (
            O => \N__23340\,
            I => \N__23296\
        );

    \I__5580\ : Span4Mux_v
    port map (
            O => \N__23333\,
            I => \N__23289\
        );

    \I__5579\ : LocalMux
    port map (
            O => \N__23330\,
            I => \N__23289\
        );

    \I__5578\ : LocalMux
    port map (
            O => \N__23327\,
            I => \N__23289\
        );

    \I__5577\ : SRMux
    port map (
            O => \N__23326\,
            I => \N__23286\
        );

    \I__5576\ : SRMux
    port map (
            O => \N__23325\,
            I => \N__23283\
        );

    \I__5575\ : IoInMux
    port map (
            O => \N__23324\,
            I => \N__23278\
        );

    \I__5574\ : IoInMux
    port map (
            O => \N__23323\,
            I => \N__23275\
        );

    \I__5573\ : Span4Mux_s3_v
    port map (
            O => \N__23318\,
            I => \N__23268\
        );

    \I__5572\ : LocalMux
    port map (
            O => \N__23315\,
            I => \N__23268\
        );

    \I__5571\ : LocalMux
    port map (
            O => \N__23312\,
            I => \N__23268\
        );

    \I__5570\ : SRMux
    port map (
            O => \N__23311\,
            I => \N__23265\
        );

    \I__5569\ : SRMux
    port map (
            O => \N__23310\,
            I => \N__23262\
        );

    \I__5568\ : CascadeMux
    port map (
            O => \N__23309\,
            I => \N__23257\
        );

    \I__5567\ : CascadeMux
    port map (
            O => \N__23308\,
            I => \N__23253\
        );

    \I__5566\ : CascadeMux
    port map (
            O => \N__23307\,
            I => \N__23249\
        );

    \I__5565\ : CascadeMux
    port map (
            O => \N__23306\,
            I => \N__23246\
        );

    \I__5564\ : CascadeMux
    port map (
            O => \N__23305\,
            I => \N__23242\
        );

    \I__5563\ : CascadeMux
    port map (
            O => \N__23304\,
            I => \N__23239\
        );

    \I__5562\ : CascadeMux
    port map (
            O => \N__23303\,
            I => \N__23235\
        );

    \I__5561\ : LocalMux
    port map (
            O => \N__23300\,
            I => \N__23232\
        );

    \I__5560\ : SRMux
    port map (
            O => \N__23299\,
            I => \N__23229\
        );

    \I__5559\ : Span4Mux_h
    port map (
            O => \N__23296\,
            I => \N__23224\
        );

    \I__5558\ : Span4Mux_v
    port map (
            O => \N__23289\,
            I => \N__23217\
        );

    \I__5557\ : LocalMux
    port map (
            O => \N__23286\,
            I => \N__23217\
        );

    \I__5556\ : LocalMux
    port map (
            O => \N__23283\,
            I => \N__23217\
        );

    \I__5555\ : SRMux
    port map (
            O => \N__23282\,
            I => \N__23214\
        );

    \I__5554\ : SRMux
    port map (
            O => \N__23281\,
            I => \N__23211\
        );

    \I__5553\ : LocalMux
    port map (
            O => \N__23278\,
            I => \N__23206\
        );

    \I__5552\ : LocalMux
    port map (
            O => \N__23275\,
            I => \N__23206\
        );

    \I__5551\ : Span4Mux_v
    port map (
            O => \N__23268\,
            I => \N__23199\
        );

    \I__5550\ : LocalMux
    port map (
            O => \N__23265\,
            I => \N__23199\
        );

    \I__5549\ : LocalMux
    port map (
            O => \N__23262\,
            I => \N__23199\
        );

    \I__5548\ : SRMux
    port map (
            O => \N__23261\,
            I => \N__23196\
        );

    \I__5547\ : SRMux
    port map (
            O => \N__23260\,
            I => \N__23193\
        );

    \I__5546\ : InMux
    port map (
            O => \N__23257\,
            I => \N__23178\
        );

    \I__5545\ : InMux
    port map (
            O => \N__23256\,
            I => \N__23178\
        );

    \I__5544\ : InMux
    port map (
            O => \N__23253\,
            I => \N__23178\
        );

    \I__5543\ : InMux
    port map (
            O => \N__23252\,
            I => \N__23178\
        );

    \I__5542\ : InMux
    port map (
            O => \N__23249\,
            I => \N__23178\
        );

    \I__5541\ : InMux
    port map (
            O => \N__23246\,
            I => \N__23175\
        );

    \I__5540\ : InMux
    port map (
            O => \N__23245\,
            I => \N__23164\
        );

    \I__5539\ : InMux
    port map (
            O => \N__23242\,
            I => \N__23164\
        );

    \I__5538\ : InMux
    port map (
            O => \N__23239\,
            I => \N__23164\
        );

    \I__5537\ : InMux
    port map (
            O => \N__23238\,
            I => \N__23164\
        );

    \I__5536\ : InMux
    port map (
            O => \N__23235\,
            I => \N__23164\
        );

    \I__5535\ : Span4Mux_v
    port map (
            O => \N__23232\,
            I => \N__23161\
        );

    \I__5534\ : LocalMux
    port map (
            O => \N__23229\,
            I => \N__23158\
        );

    \I__5533\ : SRMux
    port map (
            O => \N__23228\,
            I => \N__23155\
        );

    \I__5532\ : SRMux
    port map (
            O => \N__23227\,
            I => \N__23152\
        );

    \I__5531\ : Span4Mux_h
    port map (
            O => \N__23224\,
            I => \N__23143\
        );

    \I__5530\ : Span4Mux_v
    port map (
            O => \N__23217\,
            I => \N__23143\
        );

    \I__5529\ : LocalMux
    port map (
            O => \N__23214\,
            I => \N__23143\
        );

    \I__5528\ : LocalMux
    port map (
            O => \N__23211\,
            I => \N__23143\
        );

    \I__5527\ : IoSpan4Mux
    port map (
            O => \N__23206\,
            I => \N__23140\
        );

    \I__5526\ : Span4Mux_v
    port map (
            O => \N__23199\,
            I => \N__23131\
        );

    \I__5525\ : LocalMux
    port map (
            O => \N__23196\,
            I => \N__23131\
        );

    \I__5524\ : LocalMux
    port map (
            O => \N__23193\,
            I => \N__23131\
        );

    \I__5523\ : SRMux
    port map (
            O => \N__23192\,
            I => \N__23128\
        );

    \I__5522\ : SRMux
    port map (
            O => \N__23191\,
            I => \N__23125\
        );

    \I__5521\ : SRMux
    port map (
            O => \N__23190\,
            I => \N__23121\
        );

    \I__5520\ : SRMux
    port map (
            O => \N__23189\,
            I => \N__23118\
        );

    \I__5519\ : LocalMux
    port map (
            O => \N__23178\,
            I => \N__23112\
        );

    \I__5518\ : LocalMux
    port map (
            O => \N__23175\,
            I => \N__23112\
        );

    \I__5517\ : LocalMux
    port map (
            O => \N__23164\,
            I => \N__23109\
        );

    \I__5516\ : Span4Mux_h
    port map (
            O => \N__23161\,
            I => \N__23098\
        );

    \I__5515\ : Span4Mux_v
    port map (
            O => \N__23158\,
            I => \N__23098\
        );

    \I__5514\ : LocalMux
    port map (
            O => \N__23155\,
            I => \N__23098\
        );

    \I__5513\ : LocalMux
    port map (
            O => \N__23152\,
            I => \N__23098\
        );

    \I__5512\ : Span4Mux_v
    port map (
            O => \N__23143\,
            I => \N__23098\
        );

    \I__5511\ : Span4Mux_s0_v
    port map (
            O => \N__23140\,
            I => \N__23095\
        );

    \I__5510\ : SRMux
    port map (
            O => \N__23139\,
            I => \N__23092\
        );

    \I__5509\ : SRMux
    port map (
            O => \N__23138\,
            I => \N__23089\
        );

    \I__5508\ : Span4Mux_v
    port map (
            O => \N__23131\,
            I => \N__23082\
        );

    \I__5507\ : LocalMux
    port map (
            O => \N__23128\,
            I => \N__23082\
        );

    \I__5506\ : LocalMux
    port map (
            O => \N__23125\,
            I => \N__23082\
        );

    \I__5505\ : SRMux
    port map (
            O => \N__23124\,
            I => \N__23079\
        );

    \I__5504\ : LocalMux
    port map (
            O => \N__23121\,
            I => \N__23074\
        );

    \I__5503\ : LocalMux
    port map (
            O => \N__23118\,
            I => \N__23074\
        );

    \I__5502\ : SRMux
    port map (
            O => \N__23117\,
            I => \N__23071\
        );

    \I__5501\ : Sp12to4
    port map (
            O => \N__23112\,
            I => \N__23068\
        );

    \I__5500\ : Span4Mux_v
    port map (
            O => \N__23109\,
            I => \N__23065\
        );

    \I__5499\ : Span4Mux_v
    port map (
            O => \N__23098\,
            I => \N__23062\
        );

    \I__5498\ : Span4Mux_h
    port map (
            O => \N__23095\,
            I => \N__23055\
        );

    \I__5497\ : LocalMux
    port map (
            O => \N__23092\,
            I => \N__23055\
        );

    \I__5496\ : LocalMux
    port map (
            O => \N__23089\,
            I => \N__23055\
        );

    \I__5495\ : Span4Mux_v
    port map (
            O => \N__23082\,
            I => \N__23046\
        );

    \I__5494\ : LocalMux
    port map (
            O => \N__23079\,
            I => \N__23046\
        );

    \I__5493\ : Span4Mux_v
    port map (
            O => \N__23074\,
            I => \N__23046\
        );

    \I__5492\ : LocalMux
    port map (
            O => \N__23071\,
            I => \N__23046\
        );

    \I__5491\ : Span12Mux_v
    port map (
            O => \N__23068\,
            I => \N__23043\
        );

    \I__5490\ : Sp12to4
    port map (
            O => \N__23065\,
            I => \N__23040\
        );

    \I__5489\ : Sp12to4
    port map (
            O => \N__23062\,
            I => \N__23037\
        );

    \I__5488\ : Span4Mux_v
    port map (
            O => \N__23055\,
            I => \N__23032\
        );

    \I__5487\ : Span4Mux_v
    port map (
            O => \N__23046\,
            I => \N__23032\
        );

    \I__5486\ : Span12Mux_h
    port map (
            O => \N__23043\,
            I => \N__23029\
        );

    \I__5485\ : Span12Mux_h
    port map (
            O => \N__23040\,
            I => \N__23026\
        );

    \I__5484\ : Span12Mux_h
    port map (
            O => \N__23037\,
            I => \N__23023\
        );

    \I__5483\ : Span4Mux_v
    port map (
            O => \N__23032\,
            I => \N__23020\
        );

    \I__5482\ : Odrv12
    port map (
            O => \N__23029\,
            I => \CONSTANT_ONE_NET\
        );

    \I__5481\ : Odrv12
    port map (
            O => \N__23026\,
            I => \CONSTANT_ONE_NET\
        );

    \I__5480\ : Odrv12
    port map (
            O => \N__23023\,
            I => \CONSTANT_ONE_NET\
        );

    \I__5479\ : Odrv4
    port map (
            O => \N__23020\,
            I => \CONSTANT_ONE_NET\
        );

    \I__5478\ : InMux
    port map (
            O => \N__23011\,
            I => \N__23008\
        );

    \I__5477\ : LocalMux
    port map (
            O => \N__23008\,
            I => \N__23005\
        );

    \I__5476\ : Span4Mux_v
    port map (
            O => \N__23005\,
            I => \N__23002\
        );

    \I__5475\ : Sp12to4
    port map (
            O => \N__23002\,
            I => \N__22999\
        );

    \I__5474\ : Span12Mux_h
    port map (
            O => \N__22999\,
            I => \N__22996\
        );

    \I__5473\ : Span12Mux_v
    port map (
            O => \N__22996\,
            I => \N__22993\
        );

    \I__5472\ : Odrv12
    port map (
            O => \N__22993\,
            I => \line_buffer.n673\
        );

    \I__5471\ : CascadeMux
    port map (
            O => \N__22990\,
            I => \N__22987\
        );

    \I__5470\ : InMux
    port map (
            O => \N__22987\,
            I => \N__22984\
        );

    \I__5469\ : LocalMux
    port map (
            O => \N__22984\,
            I => \N__22981\
        );

    \I__5468\ : Span4Mux_v
    port map (
            O => \N__22981\,
            I => \N__22978\
        );

    \I__5467\ : Sp12to4
    port map (
            O => \N__22978\,
            I => \N__22975\
        );

    \I__5466\ : Odrv12
    port map (
            O => \N__22975\,
            I => \line_buffer.n681\
        );

    \I__5465\ : InMux
    port map (
            O => \N__22972\,
            I => \N__22969\
        );

    \I__5464\ : LocalMux
    port map (
            O => \N__22969\,
            I => \line_buffer.n4146\
        );

    \I__5463\ : InMux
    port map (
            O => \N__22966\,
            I => \N__22963\
        );

    \I__5462\ : LocalMux
    port map (
            O => \N__22963\,
            I => \line_buffer.n4149\
        );

    \I__5461\ : InMux
    port map (
            O => \N__22960\,
            I => \N__22957\
        );

    \I__5460\ : LocalMux
    port map (
            O => \N__22957\,
            I => \N__22954\
        );

    \I__5459\ : Span4Mux_h
    port map (
            O => \N__22954\,
            I => \N__22951\
        );

    \I__5458\ : Span4Mux_h
    port map (
            O => \N__22951\,
            I => \N__22948\
        );

    \I__5457\ : Odrv4
    port map (
            O => \N__22948\,
            I => \TX_DATA_0\
        );

    \I__5456\ : InMux
    port map (
            O => \N__22945\,
            I => \N__22942\
        );

    \I__5455\ : LocalMux
    port map (
            O => \N__22942\,
            I => \N__22939\
        );

    \I__5454\ : Span12Mux_v
    port map (
            O => \N__22939\,
            I => \N__22936\
        );

    \I__5453\ : Odrv12
    port map (
            O => \N__22936\,
            I => \line_buffer.n621\
        );

    \I__5452\ : InMux
    port map (
            O => \N__22933\,
            I => \N__22930\
        );

    \I__5451\ : LocalMux
    port map (
            O => \N__22930\,
            I => \N__22927\
        );

    \I__5450\ : Span4Mux_v
    port map (
            O => \N__22927\,
            I => \N__22924\
        );

    \I__5449\ : Span4Mux_h
    port map (
            O => \N__22924\,
            I => \N__22921\
        );

    \I__5448\ : Odrv4
    port map (
            O => \N__22921\,
            I => \line_buffer.n613\
        );

    \I__5447\ : InMux
    port map (
            O => \N__22918\,
            I => \N__22915\
        );

    \I__5446\ : LocalMux
    port map (
            O => \N__22915\,
            I => \N__22912\
        );

    \I__5445\ : Span12Mux_v
    port map (
            O => \N__22912\,
            I => \N__22909\
        );

    \I__5444\ : Odrv12
    port map (
            O => \N__22909\,
            I => \line_buffer.n653\
        );

    \I__5443\ : InMux
    port map (
            O => \N__22906\,
            I => \N__22903\
        );

    \I__5442\ : LocalMux
    port map (
            O => \N__22903\,
            I => \N__22900\
        );

    \I__5441\ : Span4Mux_v
    port map (
            O => \N__22900\,
            I => \N__22897\
        );

    \I__5440\ : Span4Mux_h
    port map (
            O => \N__22897\,
            I => \N__22894\
        );

    \I__5439\ : Odrv4
    port map (
            O => \N__22894\,
            I => \line_buffer.n645\
        );

    \I__5438\ : InMux
    port map (
            O => \N__22891\,
            I => \N__22888\
        );

    \I__5437\ : LocalMux
    port map (
            O => \N__22888\,
            I => \N__22885\
        );

    \I__5436\ : Odrv12
    port map (
            O => \N__22885\,
            I => \line_buffer.n4062\
        );

    \I__5435\ : InMux
    port map (
            O => \N__22882\,
            I => \N__22879\
        );

    \I__5434\ : LocalMux
    port map (
            O => \N__22879\,
            I => \N__22876\
        );

    \I__5433\ : Odrv4
    port map (
            O => \N__22876\,
            I => \line_buffer.n4078\
        );

    \I__5432\ : IoInMux
    port map (
            O => \N__22873\,
            I => \N__22870\
        );

    \I__5431\ : LocalMux
    port map (
            O => \N__22870\,
            I => \N__22866\
        );

    \I__5430\ : CascadeMux
    port map (
            O => \N__22869\,
            I => \N__22862\
        );

    \I__5429\ : IoSpan4Mux
    port map (
            O => \N__22866\,
            I => \N__22859\
        );

    \I__5428\ : InMux
    port map (
            O => \N__22865\,
            I => \N__22853\
        );

    \I__5427\ : InMux
    port map (
            O => \N__22862\,
            I => \N__22850\
        );

    \I__5426\ : IoSpan4Mux
    port map (
            O => \N__22859\,
            I => \N__22847\
        );

    \I__5425\ : CascadeMux
    port map (
            O => \N__22858\,
            I => \N__22843\
        );

    \I__5424\ : CascadeMux
    port map (
            O => \N__22857\,
            I => \N__22839\
        );

    \I__5423\ : InMux
    port map (
            O => \N__22856\,
            I => \N__22836\
        );

    \I__5422\ : LocalMux
    port map (
            O => \N__22853\,
            I => \N__22830\
        );

    \I__5421\ : LocalMux
    port map (
            O => \N__22850\,
            I => \N__22830\
        );

    \I__5420\ : Span4Mux_s2_h
    port map (
            O => \N__22847\,
            I => \N__22826\
        );

    \I__5419\ : InMux
    port map (
            O => \N__22846\,
            I => \N__22823\
        );

    \I__5418\ : InMux
    port map (
            O => \N__22843\,
            I => \N__22820\
        );

    \I__5417\ : InMux
    port map (
            O => \N__22842\,
            I => \N__22815\
        );

    \I__5416\ : InMux
    port map (
            O => \N__22839\,
            I => \N__22812\
        );

    \I__5415\ : LocalMux
    port map (
            O => \N__22836\,
            I => \N__22809\
        );

    \I__5414\ : InMux
    port map (
            O => \N__22835\,
            I => \N__22806\
        );

    \I__5413\ : Span4Mux_v
    port map (
            O => \N__22830\,
            I => \N__22803\
        );

    \I__5412\ : InMux
    port map (
            O => \N__22829\,
            I => \N__22799\
        );

    \I__5411\ : Span4Mux_h
    port map (
            O => \N__22826\,
            I => \N__22794\
        );

    \I__5410\ : LocalMux
    port map (
            O => \N__22823\,
            I => \N__22794\
        );

    \I__5409\ : LocalMux
    port map (
            O => \N__22820\,
            I => \N__22790\
        );

    \I__5408\ : InMux
    port map (
            O => \N__22819\,
            I => \N__22787\
        );

    \I__5407\ : InMux
    port map (
            O => \N__22818\,
            I => \N__22784\
        );

    \I__5406\ : LocalMux
    port map (
            O => \N__22815\,
            I => \N__22779\
        );

    \I__5405\ : LocalMux
    port map (
            O => \N__22812\,
            I => \N__22779\
        );

    \I__5404\ : Span4Mux_v
    port map (
            O => \N__22809\,
            I => \N__22776\
        );

    \I__5403\ : LocalMux
    port map (
            O => \N__22806\,
            I => \N__22771\
        );

    \I__5402\ : Span4Mux_v
    port map (
            O => \N__22803\,
            I => \N__22771\
        );

    \I__5401\ : InMux
    port map (
            O => \N__22802\,
            I => \N__22768\
        );

    \I__5400\ : LocalMux
    port map (
            O => \N__22799\,
            I => \N__22765\
        );

    \I__5399\ : Span4Mux_h
    port map (
            O => \N__22794\,
            I => \N__22761\
        );

    \I__5398\ : InMux
    port map (
            O => \N__22793\,
            I => \N__22758\
        );

    \I__5397\ : Span4Mux_v
    port map (
            O => \N__22790\,
            I => \N__22755\
        );

    \I__5396\ : LocalMux
    port map (
            O => \N__22787\,
            I => \N__22748\
        );

    \I__5395\ : LocalMux
    port map (
            O => \N__22784\,
            I => \N__22748\
        );

    \I__5394\ : Span4Mux_v
    port map (
            O => \N__22779\,
            I => \N__22748\
        );

    \I__5393\ : Span4Mux_v
    port map (
            O => \N__22776\,
            I => \N__22741\
        );

    \I__5392\ : Span4Mux_h
    port map (
            O => \N__22771\,
            I => \N__22741\
        );

    \I__5391\ : LocalMux
    port map (
            O => \N__22768\,
            I => \N__22741\
        );

    \I__5390\ : Span4Mux_h
    port map (
            O => \N__22765\,
            I => \N__22738\
        );

    \I__5389\ : InMux
    port map (
            O => \N__22764\,
            I => \N__22735\
        );

    \I__5388\ : Span4Mux_v
    port map (
            O => \N__22761\,
            I => \N__22726\
        );

    \I__5387\ : LocalMux
    port map (
            O => \N__22758\,
            I => \N__22726\
        );

    \I__5386\ : Span4Mux_v
    port map (
            O => \N__22755\,
            I => \N__22726\
        );

    \I__5385\ : Span4Mux_h
    port map (
            O => \N__22748\,
            I => \N__22726\
        );

    \I__5384\ : Span4Mux_h
    port map (
            O => \N__22741\,
            I => \N__22723\
        );

    \I__5383\ : Odrv4
    port map (
            O => \N__22738\,
            I => \DEBUG_c_2\
        );

    \I__5382\ : LocalMux
    port map (
            O => \N__22735\,
            I => \DEBUG_c_2\
        );

    \I__5381\ : Odrv4
    port map (
            O => \N__22726\,
            I => \DEBUG_c_2\
        );

    \I__5380\ : Odrv4
    port map (
            O => \N__22723\,
            I => \DEBUG_c_2\
        );

    \I__5379\ : InMux
    port map (
            O => \N__22714\,
            I => \N__22711\
        );

    \I__5378\ : LocalMux
    port map (
            O => \N__22711\,
            I => \line_buffer.n4140\
        );

    \I__5377\ : InMux
    port map (
            O => \N__22708\,
            I => \N__22705\
        );

    \I__5376\ : LocalMux
    port map (
            O => \N__22705\,
            I => \N__22702\
        );

    \I__5375\ : Span4Mux_h
    port map (
            O => \N__22702\,
            I => \N__22699\
        );

    \I__5374\ : Span4Mux_h
    port map (
            O => \N__22699\,
            I => \N__22696\
        );

    \I__5373\ : Span4Mux_v
    port map (
            O => \N__22696\,
            I => \N__22693\
        );

    \I__5372\ : Odrv4
    port map (
            O => \N__22693\,
            I => \TX_DATA_4\
        );

    \I__5371\ : ClkMux
    port map (
            O => \N__22690\,
            I => \N__22685\
        );

    \I__5370\ : ClkMux
    port map (
            O => \N__22689\,
            I => \N__22681\
        );

    \I__5369\ : ClkMux
    port map (
            O => \N__22688\,
            I => \N__22678\
        );

    \I__5368\ : LocalMux
    port map (
            O => \N__22685\,
            I => \N__22672\
        );

    \I__5367\ : ClkMux
    port map (
            O => \N__22684\,
            I => \N__22669\
        );

    \I__5366\ : LocalMux
    port map (
            O => \N__22681\,
            I => \N__22665\
        );

    \I__5365\ : LocalMux
    port map (
            O => \N__22678\,
            I => \N__22662\
        );

    \I__5364\ : ClkMux
    port map (
            O => \N__22677\,
            I => \N__22659\
        );

    \I__5363\ : ClkMux
    port map (
            O => \N__22676\,
            I => \N__22656\
        );

    \I__5362\ : ClkMux
    port map (
            O => \N__22675\,
            I => \N__22651\
        );

    \I__5361\ : Span4Mux_s2_v
    port map (
            O => \N__22672\,
            I => \N__22644\
        );

    \I__5360\ : LocalMux
    port map (
            O => \N__22669\,
            I => \N__22644\
        );

    \I__5359\ : ClkMux
    port map (
            O => \N__22668\,
            I => \N__22641\
        );

    \I__5358\ : Span4Mux_s2_v
    port map (
            O => \N__22665\,
            I => \N__22633\
        );

    \I__5357\ : Span4Mux_h
    port map (
            O => \N__22662\,
            I => \N__22633\
        );

    \I__5356\ : LocalMux
    port map (
            O => \N__22659\,
            I => \N__22633\
        );

    \I__5355\ : LocalMux
    port map (
            O => \N__22656\,
            I => \N__22630\
        );

    \I__5354\ : ClkMux
    port map (
            O => \N__22655\,
            I => \N__22627\
        );

    \I__5353\ : ClkMux
    port map (
            O => \N__22654\,
            I => \N__22624\
        );

    \I__5352\ : LocalMux
    port map (
            O => \N__22651\,
            I => \N__22616\
        );

    \I__5351\ : ClkMux
    port map (
            O => \N__22650\,
            I => \N__22613\
        );

    \I__5350\ : ClkMux
    port map (
            O => \N__22649\,
            I => \N__22610\
        );

    \I__5349\ : Span4Mux_v
    port map (
            O => \N__22644\,
            I => \N__22604\
        );

    \I__5348\ : LocalMux
    port map (
            O => \N__22641\,
            I => \N__22604\
        );

    \I__5347\ : ClkMux
    port map (
            O => \N__22640\,
            I => \N__22601\
        );

    \I__5346\ : Span4Mux_v
    port map (
            O => \N__22633\,
            I => \N__22593\
        );

    \I__5345\ : Span4Mux_h
    port map (
            O => \N__22630\,
            I => \N__22593\
        );

    \I__5344\ : LocalMux
    port map (
            O => \N__22627\,
            I => \N__22593\
        );

    \I__5343\ : LocalMux
    port map (
            O => \N__22624\,
            I => \N__22590\
        );

    \I__5342\ : ClkMux
    port map (
            O => \N__22623\,
            I => \N__22587\
        );

    \I__5341\ : ClkMux
    port map (
            O => \N__22622\,
            I => \N__22584\
        );

    \I__5340\ : ClkMux
    port map (
            O => \N__22621\,
            I => \N__22575\
        );

    \I__5339\ : ClkMux
    port map (
            O => \N__22620\,
            I => \N__22569\
        );

    \I__5338\ : ClkMux
    port map (
            O => \N__22619\,
            I => \N__22566\
        );

    \I__5337\ : Span4Mux_v
    port map (
            O => \N__22616\,
            I => \N__22555\
        );

    \I__5336\ : LocalMux
    port map (
            O => \N__22613\,
            I => \N__22555\
        );

    \I__5335\ : LocalMux
    port map (
            O => \N__22610\,
            I => \N__22552\
        );

    \I__5334\ : ClkMux
    port map (
            O => \N__22609\,
            I => \N__22549\
        );

    \I__5333\ : Span4Mux_h
    port map (
            O => \N__22604\,
            I => \N__22542\
        );

    \I__5332\ : LocalMux
    port map (
            O => \N__22601\,
            I => \N__22542\
        );

    \I__5331\ : ClkMux
    port map (
            O => \N__22600\,
            I => \N__22539\
        );

    \I__5330\ : Span4Mux_v
    port map (
            O => \N__22593\,
            I => \N__22526\
        );

    \I__5329\ : Span4Mux_h
    port map (
            O => \N__22590\,
            I => \N__22526\
        );

    \I__5328\ : LocalMux
    port map (
            O => \N__22587\,
            I => \N__22526\
        );

    \I__5327\ : LocalMux
    port map (
            O => \N__22584\,
            I => \N__22523\
        );

    \I__5326\ : ClkMux
    port map (
            O => \N__22583\,
            I => \N__22520\
        );

    \I__5325\ : ClkMux
    port map (
            O => \N__22582\,
            I => \N__22517\
        );

    \I__5324\ : ClkMux
    port map (
            O => \N__22581\,
            I => \N__22509\
        );

    \I__5323\ : ClkMux
    port map (
            O => \N__22580\,
            I => \N__22506\
        );

    \I__5322\ : ClkMux
    port map (
            O => \N__22579\,
            I => \N__22503\
        );

    \I__5321\ : ClkMux
    port map (
            O => \N__22578\,
            I => \N__22500\
        );

    \I__5320\ : LocalMux
    port map (
            O => \N__22575\,
            I => \N__22495\
        );

    \I__5319\ : ClkMux
    port map (
            O => \N__22574\,
            I => \N__22492\
        );

    \I__5318\ : ClkMux
    port map (
            O => \N__22573\,
            I => \N__22489\
        );

    \I__5317\ : ClkMux
    port map (
            O => \N__22572\,
            I => \N__22483\
        );

    \I__5316\ : LocalMux
    port map (
            O => \N__22569\,
            I => \N__22478\
        );

    \I__5315\ : LocalMux
    port map (
            O => \N__22566\,
            I => \N__22478\
        );

    \I__5314\ : ClkMux
    port map (
            O => \N__22565\,
            I => \N__22475\
        );

    \I__5313\ : ClkMux
    port map (
            O => \N__22564\,
            I => \N__22471\
        );

    \I__5312\ : ClkMux
    port map (
            O => \N__22563\,
            I => \N__22467\
        );

    \I__5311\ : ClkMux
    port map (
            O => \N__22562\,
            I => \N__22462\
        );

    \I__5310\ : ClkMux
    port map (
            O => \N__22561\,
            I => \N__22459\
        );

    \I__5309\ : ClkMux
    port map (
            O => \N__22560\,
            I => \N__22456\
        );

    \I__5308\ : Span4Mux_h
    port map (
            O => \N__22555\,
            I => \N__22449\
        );

    \I__5307\ : Span4Mux_h
    port map (
            O => \N__22552\,
            I => \N__22449\
        );

    \I__5306\ : LocalMux
    port map (
            O => \N__22549\,
            I => \N__22449\
        );

    \I__5305\ : ClkMux
    port map (
            O => \N__22548\,
            I => \N__22446\
        );

    \I__5304\ : ClkMux
    port map (
            O => \N__22547\,
            I => \N__22441\
        );

    \I__5303\ : Span4Mux_v
    port map (
            O => \N__22542\,
            I => \N__22429\
        );

    \I__5302\ : LocalMux
    port map (
            O => \N__22539\,
            I => \N__22429\
        );

    \I__5301\ : ClkMux
    port map (
            O => \N__22538\,
            I => \N__22426\
        );

    \I__5300\ : ClkMux
    port map (
            O => \N__22537\,
            I => \N__22423\
        );

    \I__5299\ : IoInMux
    port map (
            O => \N__22536\,
            I => \N__22416\
        );

    \I__5298\ : ClkMux
    port map (
            O => \N__22535\,
            I => \N__22413\
        );

    \I__5297\ : ClkMux
    port map (
            O => \N__22534\,
            I => \N__22410\
        );

    \I__5296\ : ClkMux
    port map (
            O => \N__22533\,
            I => \N__22404\
        );

    \I__5295\ : Span4Mux_v
    port map (
            O => \N__22526\,
            I => \N__22397\
        );

    \I__5294\ : Span4Mux_h
    port map (
            O => \N__22523\,
            I => \N__22397\
        );

    \I__5293\ : LocalMux
    port map (
            O => \N__22520\,
            I => \N__22397\
        );

    \I__5292\ : LocalMux
    port map (
            O => \N__22517\,
            I => \N__22394\
        );

    \I__5291\ : ClkMux
    port map (
            O => \N__22516\,
            I => \N__22391\
        );

    \I__5290\ : ClkMux
    port map (
            O => \N__22515\,
            I => \N__22388\
        );

    \I__5289\ : ClkMux
    port map (
            O => \N__22514\,
            I => \N__22383\
        );

    \I__5288\ : ClkMux
    port map (
            O => \N__22513\,
            I => \N__22380\
        );

    \I__5287\ : ClkMux
    port map (
            O => \N__22512\,
            I => \N__22377\
        );

    \I__5286\ : LocalMux
    port map (
            O => \N__22509\,
            I => \N__22374\
        );

    \I__5285\ : LocalMux
    port map (
            O => \N__22506\,
            I => \N__22371\
        );

    \I__5284\ : LocalMux
    port map (
            O => \N__22503\,
            I => \N__22366\
        );

    \I__5283\ : LocalMux
    port map (
            O => \N__22500\,
            I => \N__22366\
        );

    \I__5282\ : ClkMux
    port map (
            O => \N__22499\,
            I => \N__22363\
        );

    \I__5281\ : ClkMux
    port map (
            O => \N__22498\,
            I => \N__22360\
        );

    \I__5280\ : Span4Mux_v
    port map (
            O => \N__22495\,
            I => \N__22353\
        );

    \I__5279\ : LocalMux
    port map (
            O => \N__22492\,
            I => \N__22353\
        );

    \I__5278\ : LocalMux
    port map (
            O => \N__22489\,
            I => \N__22353\
        );

    \I__5277\ : ClkMux
    port map (
            O => \N__22488\,
            I => \N__22349\
        );

    \I__5276\ : ClkMux
    port map (
            O => \N__22487\,
            I => \N__22344\
        );

    \I__5275\ : ClkMux
    port map (
            O => \N__22486\,
            I => \N__22341\
        );

    \I__5274\ : LocalMux
    port map (
            O => \N__22483\,
            I => \N__22337\
        );

    \I__5273\ : Span4Mux_h
    port map (
            O => \N__22478\,
            I => \N__22332\
        );

    \I__5272\ : LocalMux
    port map (
            O => \N__22475\,
            I => \N__22332\
        );

    \I__5271\ : ClkMux
    port map (
            O => \N__22474\,
            I => \N__22329\
        );

    \I__5270\ : LocalMux
    port map (
            O => \N__22471\,
            I => \N__22326\
        );

    \I__5269\ : ClkMux
    port map (
            O => \N__22470\,
            I => \N__22323\
        );

    \I__5268\ : LocalMux
    port map (
            O => \N__22467\,
            I => \N__22319\
        );

    \I__5267\ : ClkMux
    port map (
            O => \N__22466\,
            I => \N__22316\
        );

    \I__5266\ : ClkMux
    port map (
            O => \N__22465\,
            I => \N__22311\
        );

    \I__5265\ : LocalMux
    port map (
            O => \N__22462\,
            I => \N__22308\
        );

    \I__5264\ : LocalMux
    port map (
            O => \N__22459\,
            I => \N__22303\
        );

    \I__5263\ : LocalMux
    port map (
            O => \N__22456\,
            I => \N__22303\
        );

    \I__5262\ : Span4Mux_h
    port map (
            O => \N__22449\,
            I => \N__22298\
        );

    \I__5261\ : LocalMux
    port map (
            O => \N__22446\,
            I => \N__22298\
        );

    \I__5260\ : ClkMux
    port map (
            O => \N__22445\,
            I => \N__22295\
        );

    \I__5259\ : ClkMux
    port map (
            O => \N__22444\,
            I => \N__22292\
        );

    \I__5258\ : LocalMux
    port map (
            O => \N__22441\,
            I => \N__22289\
        );

    \I__5257\ : ClkMux
    port map (
            O => \N__22440\,
            I => \N__22286\
        );

    \I__5256\ : ClkMux
    port map (
            O => \N__22439\,
            I => \N__22283\
        );

    \I__5255\ : ClkMux
    port map (
            O => \N__22438\,
            I => \N__22279\
        );

    \I__5254\ : ClkMux
    port map (
            O => \N__22437\,
            I => \N__22276\
        );

    \I__5253\ : ClkMux
    port map (
            O => \N__22436\,
            I => \N__22273\
        );

    \I__5252\ : ClkMux
    port map (
            O => \N__22435\,
            I => \N__22270\
        );

    \I__5251\ : ClkMux
    port map (
            O => \N__22434\,
            I => \N__22267\
        );

    \I__5250\ : Span4Mux_h
    port map (
            O => \N__22429\,
            I => \N__22263\
        );

    \I__5249\ : LocalMux
    port map (
            O => \N__22426\,
            I => \N__22258\
        );

    \I__5248\ : LocalMux
    port map (
            O => \N__22423\,
            I => \N__22258\
        );

    \I__5247\ : ClkMux
    port map (
            O => \N__22422\,
            I => \N__22255\
        );

    \I__5246\ : ClkMux
    port map (
            O => \N__22421\,
            I => \N__22252\
        );

    \I__5245\ : ClkMux
    port map (
            O => \N__22420\,
            I => \N__22249\
        );

    \I__5244\ : ClkMux
    port map (
            O => \N__22419\,
            I => \N__22244\
        );

    \I__5243\ : LocalMux
    port map (
            O => \N__22416\,
            I => \N__22240\
        );

    \I__5242\ : LocalMux
    port map (
            O => \N__22413\,
            I => \N__22234\
        );

    \I__5241\ : LocalMux
    port map (
            O => \N__22410\,
            I => \N__22234\
        );

    \I__5240\ : ClkMux
    port map (
            O => \N__22409\,
            I => \N__22231\
        );

    \I__5239\ : ClkMux
    port map (
            O => \N__22408\,
            I => \N__22226\
        );

    \I__5238\ : ClkMux
    port map (
            O => \N__22407\,
            I => \N__22222\
        );

    \I__5237\ : LocalMux
    port map (
            O => \N__22404\,
            I => \N__22219\
        );

    \I__5236\ : Span4Mux_v
    port map (
            O => \N__22397\,
            I => \N__22212\
        );

    \I__5235\ : Span4Mux_h
    port map (
            O => \N__22394\,
            I => \N__22212\
        );

    \I__5234\ : LocalMux
    port map (
            O => \N__22391\,
            I => \N__22212\
        );

    \I__5233\ : LocalMux
    port map (
            O => \N__22388\,
            I => \N__22209\
        );

    \I__5232\ : ClkMux
    port map (
            O => \N__22387\,
            I => \N__22206\
        );

    \I__5231\ : ClkMux
    port map (
            O => \N__22386\,
            I => \N__22202\
        );

    \I__5230\ : LocalMux
    port map (
            O => \N__22383\,
            I => \N__22199\
        );

    \I__5229\ : LocalMux
    port map (
            O => \N__22380\,
            I => \N__22196\
        );

    \I__5228\ : LocalMux
    port map (
            O => \N__22377\,
            I => \N__22193\
        );

    \I__5227\ : Span4Mux_h
    port map (
            O => \N__22374\,
            I => \N__22180\
        );

    \I__5226\ : Span4Mux_v
    port map (
            O => \N__22371\,
            I => \N__22180\
        );

    \I__5225\ : Span4Mux_h
    port map (
            O => \N__22366\,
            I => \N__22180\
        );

    \I__5224\ : LocalMux
    port map (
            O => \N__22363\,
            I => \N__22180\
        );

    \I__5223\ : LocalMux
    port map (
            O => \N__22360\,
            I => \N__22180\
        );

    \I__5222\ : Span4Mux_h
    port map (
            O => \N__22353\,
            I => \N__22180\
        );

    \I__5221\ : ClkMux
    port map (
            O => \N__22352\,
            I => \N__22177\
        );

    \I__5220\ : LocalMux
    port map (
            O => \N__22349\,
            I => \N__22174\
        );

    \I__5219\ : ClkMux
    port map (
            O => \N__22348\,
            I => \N__22171\
        );

    \I__5218\ : ClkMux
    port map (
            O => \N__22347\,
            I => \N__22168\
        );

    \I__5217\ : LocalMux
    port map (
            O => \N__22344\,
            I => \N__22165\
        );

    \I__5216\ : LocalMux
    port map (
            O => \N__22341\,
            I => \N__22162\
        );

    \I__5215\ : ClkMux
    port map (
            O => \N__22340\,
            I => \N__22159\
        );

    \I__5214\ : Span4Mux_h
    port map (
            O => \N__22337\,
            I => \N__22154\
        );

    \I__5213\ : Span4Mux_h
    port map (
            O => \N__22332\,
            I => \N__22154\
        );

    \I__5212\ : LocalMux
    port map (
            O => \N__22329\,
            I => \N__22151\
        );

    \I__5211\ : Span4Mux_h
    port map (
            O => \N__22326\,
            I => \N__22146\
        );

    \I__5210\ : LocalMux
    port map (
            O => \N__22323\,
            I => \N__22146\
        );

    \I__5209\ : ClkMux
    port map (
            O => \N__22322\,
            I => \N__22143\
        );

    \I__5208\ : Span4Mux_h
    port map (
            O => \N__22319\,
            I => \N__22140\
        );

    \I__5207\ : LocalMux
    port map (
            O => \N__22316\,
            I => \N__22137\
        );

    \I__5206\ : ClkMux
    port map (
            O => \N__22315\,
            I => \N__22134\
        );

    \I__5205\ : ClkMux
    port map (
            O => \N__22314\,
            I => \N__22131\
        );

    \I__5204\ : LocalMux
    port map (
            O => \N__22311\,
            I => \N__22128\
        );

    \I__5203\ : Span4Mux_h
    port map (
            O => \N__22308\,
            I => \N__22117\
        );

    \I__5202\ : Span4Mux_h
    port map (
            O => \N__22303\,
            I => \N__22117\
        );

    \I__5201\ : Span4Mux_h
    port map (
            O => \N__22298\,
            I => \N__22117\
        );

    \I__5200\ : LocalMux
    port map (
            O => \N__22295\,
            I => \N__22117\
        );

    \I__5199\ : LocalMux
    port map (
            O => \N__22292\,
            I => \N__22117\
        );

    \I__5198\ : Span4Mux_h
    port map (
            O => \N__22289\,
            I => \N__22112\
        );

    \I__5197\ : LocalMux
    port map (
            O => \N__22286\,
            I => \N__22112\
        );

    \I__5196\ : LocalMux
    port map (
            O => \N__22283\,
            I => \N__22109\
        );

    \I__5195\ : ClkMux
    port map (
            O => \N__22282\,
            I => \N__22106\
        );

    \I__5194\ : LocalMux
    port map (
            O => \N__22279\,
            I => \N__22101\
        );

    \I__5193\ : LocalMux
    port map (
            O => \N__22276\,
            I => \N__22101\
        );

    \I__5192\ : LocalMux
    port map (
            O => \N__22273\,
            I => \N__22096\
        );

    \I__5191\ : LocalMux
    port map (
            O => \N__22270\,
            I => \N__22096\
        );

    \I__5190\ : LocalMux
    port map (
            O => \N__22267\,
            I => \N__22093\
        );

    \I__5189\ : ClkMux
    port map (
            O => \N__22266\,
            I => \N__22090\
        );

    \I__5188\ : Span4Mux_v
    port map (
            O => \N__22263\,
            I => \N__22083\
        );

    \I__5187\ : Span4Mux_h
    port map (
            O => \N__22258\,
            I => \N__22083\
        );

    \I__5186\ : LocalMux
    port map (
            O => \N__22255\,
            I => \N__22083\
        );

    \I__5185\ : LocalMux
    port map (
            O => \N__22252\,
            I => \N__22080\
        );

    \I__5184\ : LocalMux
    port map (
            O => \N__22249\,
            I => \N__22077\
        );

    \I__5183\ : ClkMux
    port map (
            O => \N__22248\,
            I => \N__22074\
        );

    \I__5182\ : ClkMux
    port map (
            O => \N__22247\,
            I => \N__22071\
        );

    \I__5181\ : LocalMux
    port map (
            O => \N__22244\,
            I => \N__22066\
        );

    \I__5180\ : ClkMux
    port map (
            O => \N__22243\,
            I => \N__22063\
        );

    \I__5179\ : IoSpan4Mux
    port map (
            O => \N__22240\,
            I => \N__22058\
        );

    \I__5178\ : ClkMux
    port map (
            O => \N__22239\,
            I => \N__22055\
        );

    \I__5177\ : Span4Mux_v
    port map (
            O => \N__22234\,
            I => \N__22050\
        );

    \I__5176\ : LocalMux
    port map (
            O => \N__22231\,
            I => \N__22050\
        );

    \I__5175\ : ClkMux
    port map (
            O => \N__22230\,
            I => \N__22047\
        );

    \I__5174\ : ClkMux
    port map (
            O => \N__22229\,
            I => \N__22044\
        );

    \I__5173\ : LocalMux
    port map (
            O => \N__22226\,
            I => \N__22041\
        );

    \I__5172\ : ClkMux
    port map (
            O => \N__22225\,
            I => \N__22038\
        );

    \I__5171\ : LocalMux
    port map (
            O => \N__22222\,
            I => \N__22034\
        );

    \I__5170\ : Span4Mux_v
    port map (
            O => \N__22219\,
            I => \N__22031\
        );

    \I__5169\ : Span4Mux_v
    port map (
            O => \N__22212\,
            I => \N__22024\
        );

    \I__5168\ : Span4Mux_h
    port map (
            O => \N__22209\,
            I => \N__22024\
        );

    \I__5167\ : LocalMux
    port map (
            O => \N__22206\,
            I => \N__22024\
        );

    \I__5166\ : ClkMux
    port map (
            O => \N__22205\,
            I => \N__22021\
        );

    \I__5165\ : LocalMux
    port map (
            O => \N__22202\,
            I => \N__22017\
        );

    \I__5164\ : Span4Mux_v
    port map (
            O => \N__22199\,
            I => \N__22006\
        );

    \I__5163\ : Span4Mux_v
    port map (
            O => \N__22196\,
            I => \N__22006\
        );

    \I__5162\ : Span4Mux_h
    port map (
            O => \N__22193\,
            I => \N__22006\
        );

    \I__5161\ : Span4Mux_h
    port map (
            O => \N__22180\,
            I => \N__22006\
        );

    \I__5160\ : LocalMux
    port map (
            O => \N__22177\,
            I => \N__22006\
        );

    \I__5159\ : Span4Mux_h
    port map (
            O => \N__22174\,
            I => \N__21999\
        );

    \I__5158\ : LocalMux
    port map (
            O => \N__22171\,
            I => \N__21999\
        );

    \I__5157\ : LocalMux
    port map (
            O => \N__22168\,
            I => \N__21999\
        );

    \I__5156\ : Span4Mux_v
    port map (
            O => \N__22165\,
            I => \N__21992\
        );

    \I__5155\ : Span4Mux_h
    port map (
            O => \N__22162\,
            I => \N__21992\
        );

    \I__5154\ : LocalMux
    port map (
            O => \N__22159\,
            I => \N__21992\
        );

    \I__5153\ : Span4Mux_v
    port map (
            O => \N__22154\,
            I => \N__21985\
        );

    \I__5152\ : Span4Mux_h
    port map (
            O => \N__22151\,
            I => \N__21985\
        );

    \I__5151\ : Span4Mux_h
    port map (
            O => \N__22146\,
            I => \N__21985\
        );

    \I__5150\ : LocalMux
    port map (
            O => \N__22143\,
            I => \N__21982\
        );

    \I__5149\ : Span4Mux_h
    port map (
            O => \N__22140\,
            I => \N__21977\
        );

    \I__5148\ : Span4Mux_h
    port map (
            O => \N__22137\,
            I => \N__21977\
        );

    \I__5147\ : LocalMux
    port map (
            O => \N__22134\,
            I => \N__21972\
        );

    \I__5146\ : LocalMux
    port map (
            O => \N__22131\,
            I => \N__21972\
        );

    \I__5145\ : Span4Mux_h
    port map (
            O => \N__22128\,
            I => \N__21965\
        );

    \I__5144\ : Span4Mux_v
    port map (
            O => \N__22117\,
            I => \N__21965\
        );

    \I__5143\ : Span4Mux_h
    port map (
            O => \N__22112\,
            I => \N__21965\
        );

    \I__5142\ : Span4Mux_v
    port map (
            O => \N__22109\,
            I => \N__21960\
        );

    \I__5141\ : LocalMux
    port map (
            O => \N__22106\,
            I => \N__21960\
        );

    \I__5140\ : Span4Mux_v
    port map (
            O => \N__22101\,
            I => \N__21949\
        );

    \I__5139\ : Span4Mux_h
    port map (
            O => \N__22096\,
            I => \N__21949\
        );

    \I__5138\ : Span4Mux_h
    port map (
            O => \N__22093\,
            I => \N__21949\
        );

    \I__5137\ : LocalMux
    port map (
            O => \N__22090\,
            I => \N__21949\
        );

    \I__5136\ : Span4Mux_h
    port map (
            O => \N__22083\,
            I => \N__21938\
        );

    \I__5135\ : Span4Mux_v
    port map (
            O => \N__22080\,
            I => \N__21938\
        );

    \I__5134\ : Span4Mux_h
    port map (
            O => \N__22077\,
            I => \N__21938\
        );

    \I__5133\ : LocalMux
    port map (
            O => \N__22074\,
            I => \N__21938\
        );

    \I__5132\ : LocalMux
    port map (
            O => \N__22071\,
            I => \N__21938\
        );

    \I__5131\ : ClkMux
    port map (
            O => \N__22070\,
            I => \N__21935\
        );

    \I__5130\ : ClkMux
    port map (
            O => \N__22069\,
            I => \N__21932\
        );

    \I__5129\ : Span4Mux_h
    port map (
            O => \N__22066\,
            I => \N__21927\
        );

    \I__5128\ : LocalMux
    port map (
            O => \N__22063\,
            I => \N__21927\
        );

    \I__5127\ : ClkMux
    port map (
            O => \N__22062\,
            I => \N__21924\
        );

    \I__5126\ : ClkMux
    port map (
            O => \N__22061\,
            I => \N__21921\
        );

    \I__5125\ : Span4Mux_s1_v
    port map (
            O => \N__22058\,
            I => \N__21918\
        );

    \I__5124\ : LocalMux
    port map (
            O => \N__22055\,
            I => \N__21915\
        );

    \I__5123\ : Span4Mux_h
    port map (
            O => \N__22050\,
            I => \N__21908\
        );

    \I__5122\ : LocalMux
    port map (
            O => \N__22047\,
            I => \N__21908\
        );

    \I__5121\ : LocalMux
    port map (
            O => \N__22044\,
            I => \N__21908\
        );

    \I__5120\ : Span4Mux_v
    port map (
            O => \N__22041\,
            I => \N__21903\
        );

    \I__5119\ : LocalMux
    port map (
            O => \N__22038\,
            I => \N__21903\
        );

    \I__5118\ : ClkMux
    port map (
            O => \N__22037\,
            I => \N__21900\
        );

    \I__5117\ : Span12Mux_h
    port map (
            O => \N__22034\,
            I => \N__21897\
        );

    \I__5116\ : Sp12to4
    port map (
            O => \N__22031\,
            I => \N__21894\
        );

    \I__5115\ : Span4Mux_v
    port map (
            O => \N__22024\,
            I => \N__21891\
        );

    \I__5114\ : LocalMux
    port map (
            O => \N__22021\,
            I => \N__21888\
        );

    \I__5113\ : ClkMux
    port map (
            O => \N__22020\,
            I => \N__21885\
        );

    \I__5112\ : Span4Mux_h
    port map (
            O => \N__22017\,
            I => \N__21882\
        );

    \I__5111\ : Span4Mux_v
    port map (
            O => \N__22006\,
            I => \N__21875\
        );

    \I__5110\ : Span4Mux_h
    port map (
            O => \N__21999\,
            I => \N__21875\
        );

    \I__5109\ : Span4Mux_h
    port map (
            O => \N__21992\,
            I => \N__21875\
        );

    \I__5108\ : Span4Mux_v
    port map (
            O => \N__21985\,
            I => \N__21870\
        );

    \I__5107\ : Span4Mux_h
    port map (
            O => \N__21982\,
            I => \N__21870\
        );

    \I__5106\ : Span4Mux_v
    port map (
            O => \N__21977\,
            I => \N__21865\
        );

    \I__5105\ : Span4Mux_h
    port map (
            O => \N__21972\,
            I => \N__21865\
        );

    \I__5104\ : Span4Mux_v
    port map (
            O => \N__21965\,
            I => \N__21860\
        );

    \I__5103\ : Span4Mux_h
    port map (
            O => \N__21960\,
            I => \N__21860\
        );

    \I__5102\ : ClkMux
    port map (
            O => \N__21959\,
            I => \N__21857\
        );

    \I__5101\ : ClkMux
    port map (
            O => \N__21958\,
            I => \N__21854\
        );

    \I__5100\ : Span4Mux_h
    port map (
            O => \N__21949\,
            I => \N__21845\
        );

    \I__5099\ : Span4Mux_v
    port map (
            O => \N__21938\,
            I => \N__21845\
        );

    \I__5098\ : LocalMux
    port map (
            O => \N__21935\,
            I => \N__21845\
        );

    \I__5097\ : LocalMux
    port map (
            O => \N__21932\,
            I => \N__21845\
        );

    \I__5096\ : Span4Mux_v
    port map (
            O => \N__21927\,
            I => \N__21838\
        );

    \I__5095\ : LocalMux
    port map (
            O => \N__21924\,
            I => \N__21838\
        );

    \I__5094\ : LocalMux
    port map (
            O => \N__21921\,
            I => \N__21838\
        );

    \I__5093\ : Span4Mux_h
    port map (
            O => \N__21918\,
            I => \N__21833\
        );

    \I__5092\ : Span4Mux_h
    port map (
            O => \N__21915\,
            I => \N__21833\
        );

    \I__5091\ : Span4Mux_v
    port map (
            O => \N__21908\,
            I => \N__21830\
        );

    \I__5090\ : Span4Mux_v
    port map (
            O => \N__21903\,
            I => \N__21825\
        );

    \I__5089\ : LocalMux
    port map (
            O => \N__21900\,
            I => \N__21825\
        );

    \I__5088\ : Span12Mux_v
    port map (
            O => \N__21897\,
            I => \N__21820\
        );

    \I__5087\ : Span12Mux_h
    port map (
            O => \N__21894\,
            I => \N__21820\
        );

    \I__5086\ : Sp12to4
    port map (
            O => \N__21891\,
            I => \N__21815\
        );

    \I__5085\ : Sp12to4
    port map (
            O => \N__21888\,
            I => \N__21815\
        );

    \I__5084\ : LocalMux
    port map (
            O => \N__21885\,
            I => \N__21812\
        );

    \I__5083\ : Span4Mux_h
    port map (
            O => \N__21882\,
            I => \N__21809\
        );

    \I__5082\ : Span4Mux_v
    port map (
            O => \N__21875\,
            I => \N__21806\
        );

    \I__5081\ : Span4Mux_v
    port map (
            O => \N__21870\,
            I => \N__21801\
        );

    \I__5080\ : Span4Mux_v
    port map (
            O => \N__21865\,
            I => \N__21801\
        );

    \I__5079\ : Span4Mux_v
    port map (
            O => \N__21860\,
            I => \N__21798\
        );

    \I__5078\ : LocalMux
    port map (
            O => \N__21857\,
            I => \N__21793\
        );

    \I__5077\ : LocalMux
    port map (
            O => \N__21854\,
            I => \N__21793\
        );

    \I__5076\ : Span4Mux_v
    port map (
            O => \N__21845\,
            I => \N__21788\
        );

    \I__5075\ : Span4Mux_v
    port map (
            O => \N__21838\,
            I => \N__21788\
        );

    \I__5074\ : Span4Mux_h
    port map (
            O => \N__21833\,
            I => \N__21785\
        );

    \I__5073\ : Span4Mux_v
    port map (
            O => \N__21830\,
            I => \N__21780\
        );

    \I__5072\ : Span4Mux_h
    port map (
            O => \N__21825\,
            I => \N__21780\
        );

    \I__5071\ : Span12Mux_v
    port map (
            O => \N__21820\,
            I => \N__21773\
        );

    \I__5070\ : Span12Mux_h
    port map (
            O => \N__21815\,
            I => \N__21773\
        );

    \I__5069\ : Span12Mux_h
    port map (
            O => \N__21812\,
            I => \N__21773\
        );

    \I__5068\ : Span4Mux_h
    port map (
            O => \N__21809\,
            I => \N__21768\
        );

    \I__5067\ : Span4Mux_v
    port map (
            O => \N__21806\,
            I => \N__21768\
        );

    \I__5066\ : Span4Mux_v
    port map (
            O => \N__21801\,
            I => \N__21765\
        );

    \I__5065\ : Span4Mux_v
    port map (
            O => \N__21798\,
            I => \N__21762\
        );

    \I__5064\ : Span12Mux_h
    port map (
            O => \N__21793\,
            I => \N__21757\
        );

    \I__5063\ : Sp12to4
    port map (
            O => \N__21788\,
            I => \N__21757\
        );

    \I__5062\ : Span4Mux_h
    port map (
            O => \N__21785\,
            I => \N__21752\
        );

    \I__5061\ : Span4Mux_h
    port map (
            O => \N__21780\,
            I => \N__21752\
        );

    \I__5060\ : Odrv12
    port map (
            O => \N__21773\,
            I => \ADV_CLK_c\
        );

    \I__5059\ : Odrv4
    port map (
            O => \N__21768\,
            I => \ADV_CLK_c\
        );

    \I__5058\ : Odrv4
    port map (
            O => \N__21765\,
            I => \ADV_CLK_c\
        );

    \I__5057\ : Odrv4
    port map (
            O => \N__21762\,
            I => \ADV_CLK_c\
        );

    \I__5056\ : Odrv12
    port map (
            O => \N__21757\,
            I => \ADV_CLK_c\
        );

    \I__5055\ : Odrv4
    port map (
            O => \N__21752\,
            I => \ADV_CLK_c\
        );

    \I__5054\ : InMux
    port map (
            O => \N__21739\,
            I => \N__21736\
        );

    \I__5053\ : LocalMux
    port map (
            O => \N__21736\,
            I => \N__21733\
        );

    \I__5052\ : Span4Mux_h
    port map (
            O => \N__21733\,
            I => \N__21730\
        );

    \I__5051\ : Span4Mux_h
    port map (
            O => \N__21730\,
            I => \N__21727\
        );

    \I__5050\ : Odrv4
    port map (
            O => \N__21727\,
            I => \line_buffer.n641\
        );

    \I__5049\ : CascadeMux
    port map (
            O => \N__21724\,
            I => \N__21721\
        );

    \I__5048\ : InMux
    port map (
            O => \N__21721\,
            I => \N__21718\
        );

    \I__5047\ : LocalMux
    port map (
            O => \N__21718\,
            I => \N__21715\
        );

    \I__5046\ : Span12Mux_v
    port map (
            O => \N__21715\,
            I => \N__21712\
        );

    \I__5045\ : Odrv12
    port map (
            O => \N__21712\,
            I => \line_buffer.n649\
        );

    \I__5044\ : InMux
    port map (
            O => \N__21709\,
            I => \N__21706\
        );

    \I__5043\ : LocalMux
    port map (
            O => \N__21706\,
            I => \N__21703\
        );

    \I__5042\ : Span4Mux_v
    port map (
            O => \N__21703\,
            I => \N__21700\
        );

    \I__5041\ : Span4Mux_h
    port map (
            O => \N__21700\,
            I => \N__21697\
        );

    \I__5040\ : Odrv4
    port map (
            O => \N__21697\,
            I => \line_buffer.n552\
        );

    \I__5039\ : InMux
    port map (
            O => \N__21694\,
            I => \N__21691\
        );

    \I__5038\ : LocalMux
    port map (
            O => \N__21691\,
            I => \line_buffer.n4116\
        );

    \I__5037\ : CascadeMux
    port map (
            O => \N__21688\,
            I => \N__21685\
        );

    \I__5036\ : InMux
    port map (
            O => \N__21685\,
            I => \N__21682\
        );

    \I__5035\ : LocalMux
    port map (
            O => \N__21682\,
            I => \N__21679\
        );

    \I__5034\ : Span12Mux_h
    port map (
            O => \N__21679\,
            I => \N__21676\
        );

    \I__5033\ : Span12Mux_v
    port map (
            O => \N__21676\,
            I => \N__21673\
        );

    \I__5032\ : Odrv12
    port map (
            O => \N__21673\,
            I => \line_buffer.n544\
        );

    \I__5031\ : InMux
    port map (
            O => \N__21670\,
            I => \N__21667\
        );

    \I__5030\ : LocalMux
    port map (
            O => \N__21667\,
            I => \line_buffer.n4119\
        );

    \I__5029\ : InMux
    port map (
            O => \N__21664\,
            I => \N__21661\
        );

    \I__5028\ : LocalMux
    port map (
            O => \N__21661\,
            I => \N__21658\
        );

    \I__5027\ : Span4Mux_h
    port map (
            O => \N__21658\,
            I => \N__21655\
        );

    \I__5026\ : Span4Mux_h
    port map (
            O => \N__21655\,
            I => \N__21652\
        );

    \I__5025\ : Span4Mux_h
    port map (
            O => \N__21652\,
            I => \N__21649\
        );

    \I__5024\ : Odrv4
    port map (
            O => \N__21649\,
            I => \line_buffer.n684\
        );

    \I__5023\ : InMux
    port map (
            O => \N__21646\,
            I => \N__21643\
        );

    \I__5022\ : LocalMux
    port map (
            O => \N__21643\,
            I => \N__21640\
        );

    \I__5021\ : Span4Mux_v
    port map (
            O => \N__21640\,
            I => \N__21637\
        );

    \I__5020\ : Sp12to4
    port map (
            O => \N__21637\,
            I => \N__21634\
        );

    \I__5019\ : Span12Mux_h
    port map (
            O => \N__21634\,
            I => \N__21631\
        );

    \I__5018\ : Odrv12
    port map (
            O => \N__21631\,
            I => \line_buffer.n676\
        );

    \I__5017\ : InMux
    port map (
            O => \N__21628\,
            I => \N__21625\
        );

    \I__5016\ : LocalMux
    port map (
            O => \N__21625\,
            I => \line_buffer.n4066\
        );

    \I__5015\ : InMux
    port map (
            O => \N__21622\,
            I => \N__21619\
        );

    \I__5014\ : LocalMux
    port map (
            O => \N__21619\,
            I => \N__21616\
        );

    \I__5013\ : Span4Mux_h
    port map (
            O => \N__21616\,
            I => \N__21613\
        );

    \I__5012\ : Span4Mux_h
    port map (
            O => \N__21613\,
            I => \N__21610\
        );

    \I__5011\ : Odrv4
    port map (
            O => \N__21610\,
            I => \line_buffer.n555\
        );

    \I__5010\ : InMux
    port map (
            O => \N__21607\,
            I => \N__21604\
        );

    \I__5009\ : LocalMux
    port map (
            O => \N__21604\,
            I => \N__21601\
        );

    \I__5008\ : Span4Mux_v
    port map (
            O => \N__21601\,
            I => \N__21598\
        );

    \I__5007\ : Sp12to4
    port map (
            O => \N__21598\,
            I => \N__21595\
        );

    \I__5006\ : Span12Mux_h
    port map (
            O => \N__21595\,
            I => \N__21592\
        );

    \I__5005\ : Odrv12
    port map (
            O => \N__21592\,
            I => \line_buffer.n547\
        );

    \I__5004\ : CascadeMux
    port map (
            O => \N__21589\,
            I => \line_buffer.n4074_cascade_\
        );

    \I__5003\ : InMux
    port map (
            O => \N__21586\,
            I => \N__21583\
        );

    \I__5002\ : LocalMux
    port map (
            O => \N__21583\,
            I => \line_buffer.n4128\
        );

    \I__5001\ : InMux
    port map (
            O => \N__21580\,
            I => \N__21577\
        );

    \I__5000\ : LocalMux
    port map (
            O => \N__21577\,
            I => \N__21574\
        );

    \I__4999\ : Odrv12
    port map (
            O => \N__21574\,
            I => \TX_DATA_3\
        );

    \I__4998\ : InMux
    port map (
            O => \N__21571\,
            I => \N__21568\
        );

    \I__4997\ : LocalMux
    port map (
            O => \N__21568\,
            I => \N__21565\
        );

    \I__4996\ : Span4Mux_h
    port map (
            O => \N__21565\,
            I => \N__21562\
        );

    \I__4995\ : Span4Mux_h
    port map (
            O => \N__21562\,
            I => \N__21559\
        );

    \I__4994\ : Span4Mux_h
    port map (
            O => \N__21559\,
            I => \N__21556\
        );

    \I__4993\ : Span4Mux_v
    port map (
            O => \N__21556\,
            I => \N__21553\
        );

    \I__4992\ : Span4Mux_v
    port map (
            O => \N__21553\,
            I => \N__21550\
        );

    \I__4991\ : Odrv4
    port map (
            O => \N__21550\,
            I => \line_buffer.n652\
        );

    \I__4990\ : InMux
    port map (
            O => \N__21547\,
            I => \N__21544\
        );

    \I__4989\ : LocalMux
    port map (
            O => \N__21544\,
            I => \N__21541\
        );

    \I__4988\ : Span4Mux_v
    port map (
            O => \N__21541\,
            I => \N__21538\
        );

    \I__4987\ : Span4Mux_h
    port map (
            O => \N__21538\,
            I => \N__21535\
        );

    \I__4986\ : Span4Mux_h
    port map (
            O => \N__21535\,
            I => \N__21532\
        );

    \I__4985\ : Odrv4
    port map (
            O => \N__21532\,
            I => \line_buffer.n644\
        );

    \I__4984\ : InMux
    port map (
            O => \N__21529\,
            I => \N__21526\
        );

    \I__4983\ : LocalMux
    port map (
            O => \N__21526\,
            I => \line_buffer.n4075\
        );

    \I__4982\ : InMux
    port map (
            O => \N__21523\,
            I => \N__21520\
        );

    \I__4981\ : LocalMux
    port map (
            O => \N__21520\,
            I => \N__21517\
        );

    \I__4980\ : Span4Mux_v
    port map (
            O => \N__21517\,
            I => \N__21514\
        );

    \I__4979\ : Odrv4
    port map (
            O => \N__21514\,
            I => \transmit_module.Y_DELTA_PATTERN_33\
        );

    \I__4978\ : InMux
    port map (
            O => \N__21511\,
            I => \N__21508\
        );

    \I__4977\ : LocalMux
    port map (
            O => \N__21508\,
            I => \N__21505\
        );

    \I__4976\ : Span4Mux_v
    port map (
            O => \N__21505\,
            I => \N__21502\
        );

    \I__4975\ : Odrv4
    port map (
            O => \N__21502\,
            I => \transmit_module.Y_DELTA_PATTERN_35\
        );

    \I__4974\ : InMux
    port map (
            O => \N__21499\,
            I => \N__21496\
        );

    \I__4973\ : LocalMux
    port map (
            O => \N__21496\,
            I => \transmit_module.Y_DELTA_PATTERN_34\
        );

    \I__4972\ : CEMux
    port map (
            O => \N__21493\,
            I => \N__21490\
        );

    \I__4971\ : LocalMux
    port map (
            O => \N__21490\,
            I => \N__21484\
        );

    \I__4970\ : CEMux
    port map (
            O => \N__21489\,
            I => \N__21481\
        );

    \I__4969\ : CEMux
    port map (
            O => \N__21488\,
            I => \N__21477\
        );

    \I__4968\ : CEMux
    port map (
            O => \N__21487\,
            I => \N__21474\
        );

    \I__4967\ : Span4Mux_h
    port map (
            O => \N__21484\,
            I => \N__21468\
        );

    \I__4966\ : LocalMux
    port map (
            O => \N__21481\,
            I => \N__21468\
        );

    \I__4965\ : CEMux
    port map (
            O => \N__21480\,
            I => \N__21465\
        );

    \I__4964\ : LocalMux
    port map (
            O => \N__21477\,
            I => \N__21460\
        );

    \I__4963\ : LocalMux
    port map (
            O => \N__21474\,
            I => \N__21453\
        );

    \I__4962\ : CEMux
    port map (
            O => \N__21473\,
            I => \N__21450\
        );

    \I__4961\ : Span4Mux_v
    port map (
            O => \N__21468\,
            I => \N__21447\
        );

    \I__4960\ : LocalMux
    port map (
            O => \N__21465\,
            I => \N__21444\
        );

    \I__4959\ : CEMux
    port map (
            O => \N__21464\,
            I => \N__21441\
        );

    \I__4958\ : CEMux
    port map (
            O => \N__21463\,
            I => \N__21438\
        );

    \I__4957\ : Span4Mux_h
    port map (
            O => \N__21460\,
            I => \N__21433\
        );

    \I__4956\ : CEMux
    port map (
            O => \N__21459\,
            I => \N__21430\
        );

    \I__4955\ : CEMux
    port map (
            O => \N__21458\,
            I => \N__21427\
        );

    \I__4954\ : CEMux
    port map (
            O => \N__21457\,
            I => \N__21424\
        );

    \I__4953\ : CEMux
    port map (
            O => \N__21456\,
            I => \N__21421\
        );

    \I__4952\ : Span4Mux_v
    port map (
            O => \N__21453\,
            I => \N__21416\
        );

    \I__4951\ : LocalMux
    port map (
            O => \N__21450\,
            I => \N__21416\
        );

    \I__4950\ : Span4Mux_h
    port map (
            O => \N__21447\,
            I => \N__21409\
        );

    \I__4949\ : Span4Mux_h
    port map (
            O => \N__21444\,
            I => \N__21409\
        );

    \I__4948\ : LocalMux
    port map (
            O => \N__21441\,
            I => \N__21409\
        );

    \I__4947\ : LocalMux
    port map (
            O => \N__21438\,
            I => \N__21406\
        );

    \I__4946\ : CEMux
    port map (
            O => \N__21437\,
            I => \N__21403\
        );

    \I__4945\ : CEMux
    port map (
            O => \N__21436\,
            I => \N__21400\
        );

    \I__4944\ : Span4Mux_v
    port map (
            O => \N__21433\,
            I => \N__21395\
        );

    \I__4943\ : LocalMux
    port map (
            O => \N__21430\,
            I => \N__21395\
        );

    \I__4942\ : LocalMux
    port map (
            O => \N__21427\,
            I => \N__21392\
        );

    \I__4941\ : LocalMux
    port map (
            O => \N__21424\,
            I => \N__21389\
        );

    \I__4940\ : LocalMux
    port map (
            O => \N__21421\,
            I => \N__21386\
        );

    \I__4939\ : Span4Mux_v
    port map (
            O => \N__21416\,
            I => \N__21379\
        );

    \I__4938\ : Span4Mux_v
    port map (
            O => \N__21409\,
            I => \N__21379\
        );

    \I__4937\ : Span4Mux_h
    port map (
            O => \N__21406\,
            I => \N__21379\
        );

    \I__4936\ : LocalMux
    port map (
            O => \N__21403\,
            I => \N__21374\
        );

    \I__4935\ : LocalMux
    port map (
            O => \N__21400\,
            I => \N__21374\
        );

    \I__4934\ : Span4Mux_h
    port map (
            O => \N__21395\,
            I => \N__21371\
        );

    \I__4933\ : Span12Mux_v
    port map (
            O => \N__21392\,
            I => \N__21368\
        );

    \I__4932\ : Span4Mux_h
    port map (
            O => \N__21389\,
            I => \N__21365\
        );

    \I__4931\ : Span4Mux_v
    port map (
            O => \N__21386\,
            I => \N__21360\
        );

    \I__4930\ : Span4Mux_h
    port map (
            O => \N__21379\,
            I => \N__21360\
        );

    \I__4929\ : Span4Mux_v
    port map (
            O => \N__21374\,
            I => \N__21357\
        );

    \I__4928\ : Odrv4
    port map (
            O => \N__21371\,
            I => \transmit_module.n4225\
        );

    \I__4927\ : Odrv12
    port map (
            O => \N__21368\,
            I => \transmit_module.n4225\
        );

    \I__4926\ : Odrv4
    port map (
            O => \N__21365\,
            I => \transmit_module.n4225\
        );

    \I__4925\ : Odrv4
    port map (
            O => \N__21360\,
            I => \transmit_module.n4225\
        );

    \I__4924\ : Odrv4
    port map (
            O => \N__21357\,
            I => \transmit_module.n4225\
        );

    \I__4923\ : CascadeMux
    port map (
            O => \N__21346\,
            I => \N__21332\
        );

    \I__4922\ : SRMux
    port map (
            O => \N__21345\,
            I => \N__21329\
        );

    \I__4921\ : SRMux
    port map (
            O => \N__21344\,
            I => \N__21326\
        );

    \I__4920\ : SRMux
    port map (
            O => \N__21343\,
            I => \N__21318\
        );

    \I__4919\ : SRMux
    port map (
            O => \N__21342\,
            I => \N__21314\
        );

    \I__4918\ : SRMux
    port map (
            O => \N__21341\,
            I => \N__21311\
        );

    \I__4917\ : SRMux
    port map (
            O => \N__21340\,
            I => \N__21308\
        );

    \I__4916\ : SRMux
    port map (
            O => \N__21339\,
            I => \N__21303\
        );

    \I__4915\ : SRMux
    port map (
            O => \N__21338\,
            I => \N__21300\
        );

    \I__4914\ : SRMux
    port map (
            O => \N__21337\,
            I => \N__21297\
        );

    \I__4913\ : CascadeMux
    port map (
            O => \N__21336\,
            I => \N__21289\
        );

    \I__4912\ : CascadeMux
    port map (
            O => \N__21335\,
            I => \N__21285\
        );

    \I__4911\ : InMux
    port map (
            O => \N__21332\,
            I => \N__21282\
        );

    \I__4910\ : LocalMux
    port map (
            O => \N__21329\,
            I => \N__21273\
        );

    \I__4909\ : LocalMux
    port map (
            O => \N__21326\,
            I => \N__21273\
        );

    \I__4908\ : SRMux
    port map (
            O => \N__21325\,
            I => \N__21270\
        );

    \I__4907\ : SRMux
    port map (
            O => \N__21324\,
            I => \N__21263\
        );

    \I__4906\ : SRMux
    port map (
            O => \N__21323\,
            I => \N__21256\
        );

    \I__4905\ : SRMux
    port map (
            O => \N__21322\,
            I => \N__21253\
        );

    \I__4904\ : SRMux
    port map (
            O => \N__21321\,
            I => \N__21248\
        );

    \I__4903\ : LocalMux
    port map (
            O => \N__21318\,
            I => \N__21245\
        );

    \I__4902\ : SRMux
    port map (
            O => \N__21317\,
            I => \N__21242\
        );

    \I__4901\ : LocalMux
    port map (
            O => \N__21314\,
            I => \N__21237\
        );

    \I__4900\ : LocalMux
    port map (
            O => \N__21311\,
            I => \N__21237\
        );

    \I__4899\ : LocalMux
    port map (
            O => \N__21308\,
            I => \N__21234\
        );

    \I__4898\ : SRMux
    port map (
            O => \N__21307\,
            I => \N__21231\
        );

    \I__4897\ : SRMux
    port map (
            O => \N__21306\,
            I => \N__21228\
        );

    \I__4896\ : LocalMux
    port map (
            O => \N__21303\,
            I => \N__21225\
        );

    \I__4895\ : LocalMux
    port map (
            O => \N__21300\,
            I => \N__21220\
        );

    \I__4894\ : LocalMux
    port map (
            O => \N__21297\,
            I => \N__21220\
        );

    \I__4893\ : SRMux
    port map (
            O => \N__21296\,
            I => \N__21214\
        );

    \I__4892\ : SRMux
    port map (
            O => \N__21295\,
            I => \N__21211\
        );

    \I__4891\ : CascadeMux
    port map (
            O => \N__21294\,
            I => \N__21206\
        );

    \I__4890\ : CascadeMux
    port map (
            O => \N__21293\,
            I => \N__21203\
        );

    \I__4889\ : CascadeMux
    port map (
            O => \N__21292\,
            I => \N__21200\
        );

    \I__4888\ : InMux
    port map (
            O => \N__21289\,
            I => \N__21191\
        );

    \I__4887\ : SRMux
    port map (
            O => \N__21288\,
            I => \N__21188\
        );

    \I__4886\ : InMux
    port map (
            O => \N__21285\,
            I => \N__21185\
        );

    \I__4885\ : LocalMux
    port map (
            O => \N__21282\,
            I => \N__21182\
        );

    \I__4884\ : CascadeMux
    port map (
            O => \N__21281\,
            I => \N__21176\
        );

    \I__4883\ : CascadeMux
    port map (
            O => \N__21280\,
            I => \N__21173\
        );

    \I__4882\ : SRMux
    port map (
            O => \N__21279\,
            I => \N__21168\
        );

    \I__4881\ : SRMux
    port map (
            O => \N__21278\,
            I => \N__21163\
        );

    \I__4880\ : Span4Mux_v
    port map (
            O => \N__21273\,
            I => \N__21158\
        );

    \I__4879\ : LocalMux
    port map (
            O => \N__21270\,
            I => \N__21158\
        );

    \I__4878\ : SRMux
    port map (
            O => \N__21269\,
            I => \N__21155\
        );

    \I__4877\ : InMux
    port map (
            O => \N__21268\,
            I => \N__21152\
        );

    \I__4876\ : SRMux
    port map (
            O => \N__21267\,
            I => \N__21148\
        );

    \I__4875\ : SRMux
    port map (
            O => \N__21266\,
            I => \N__21144\
        );

    \I__4874\ : LocalMux
    port map (
            O => \N__21263\,
            I => \N__21141\
        );

    \I__4873\ : SRMux
    port map (
            O => \N__21262\,
            I => \N__21138\
        );

    \I__4872\ : SRMux
    port map (
            O => \N__21261\,
            I => \N__21135\
        );

    \I__4871\ : SRMux
    port map (
            O => \N__21260\,
            I => \N__21132\
        );

    \I__4870\ : CascadeMux
    port map (
            O => \N__21259\,
            I => \N__21129\
        );

    \I__4869\ : LocalMux
    port map (
            O => \N__21256\,
            I => \N__21124\
        );

    \I__4868\ : LocalMux
    port map (
            O => \N__21253\,
            I => \N__21124\
        );

    \I__4867\ : SRMux
    port map (
            O => \N__21252\,
            I => \N__21121\
        );

    \I__4866\ : SRMux
    port map (
            O => \N__21251\,
            I => \N__21118\
        );

    \I__4865\ : LocalMux
    port map (
            O => \N__21248\,
            I => \N__21115\
        );

    \I__4864\ : Span4Mux_h
    port map (
            O => \N__21245\,
            I => \N__21108\
        );

    \I__4863\ : LocalMux
    port map (
            O => \N__21242\,
            I => \N__21108\
        );

    \I__4862\ : Span4Mux_h
    port map (
            O => \N__21237\,
            I => \N__21108\
        );

    \I__4861\ : Span4Mux_v
    port map (
            O => \N__21234\,
            I => \N__21097\
        );

    \I__4860\ : LocalMux
    port map (
            O => \N__21231\,
            I => \N__21097\
        );

    \I__4859\ : LocalMux
    port map (
            O => \N__21228\,
            I => \N__21097\
        );

    \I__4858\ : Span4Mux_h
    port map (
            O => \N__21225\,
            I => \N__21097\
        );

    \I__4857\ : Span4Mux_h
    port map (
            O => \N__21220\,
            I => \N__21097\
        );

    \I__4856\ : CascadeMux
    port map (
            O => \N__21219\,
            I => \N__21094\
        );

    \I__4855\ : InMux
    port map (
            O => \N__21218\,
            I => \N__21087\
        );

    \I__4854\ : InMux
    port map (
            O => \N__21217\,
            I => \N__21087\
        );

    \I__4853\ : LocalMux
    port map (
            O => \N__21214\,
            I => \N__21084\
        );

    \I__4852\ : LocalMux
    port map (
            O => \N__21211\,
            I => \N__21081\
        );

    \I__4851\ : SRMux
    port map (
            O => \N__21210\,
            I => \N__21078\
        );

    \I__4850\ : InMux
    port map (
            O => \N__21209\,
            I => \N__21063\
        );

    \I__4849\ : InMux
    port map (
            O => \N__21206\,
            I => \N__21063\
        );

    \I__4848\ : InMux
    port map (
            O => \N__21203\,
            I => \N__21063\
        );

    \I__4847\ : InMux
    port map (
            O => \N__21200\,
            I => \N__21063\
        );

    \I__4846\ : InMux
    port map (
            O => \N__21199\,
            I => \N__21063\
        );

    \I__4845\ : InMux
    port map (
            O => \N__21198\,
            I => \N__21063\
        );

    \I__4844\ : InMux
    port map (
            O => \N__21197\,
            I => \N__21063\
        );

    \I__4843\ : CascadeMux
    port map (
            O => \N__21196\,
            I => \N__21060\
        );

    \I__4842\ : CascadeMux
    port map (
            O => \N__21195\,
            I => \N__21057\
        );

    \I__4841\ : CascadeMux
    port map (
            O => \N__21194\,
            I => \N__21052\
        );

    \I__4840\ : LocalMux
    port map (
            O => \N__21191\,
            I => \N__21049\
        );

    \I__4839\ : LocalMux
    port map (
            O => \N__21188\,
            I => \N__21046\
        );

    \I__4838\ : LocalMux
    port map (
            O => \N__21185\,
            I => \N__21041\
        );

    \I__4837\ : Span4Mux_h
    port map (
            O => \N__21182\,
            I => \N__21041\
        );

    \I__4836\ : SRMux
    port map (
            O => \N__21181\,
            I => \N__21038\
        );

    \I__4835\ : CascadeMux
    port map (
            O => \N__21180\,
            I => \N__21030\
        );

    \I__4834\ : InMux
    port map (
            O => \N__21179\,
            I => \N__21027\
        );

    \I__4833\ : InMux
    port map (
            O => \N__21176\,
            I => \N__21024\
        );

    \I__4832\ : InMux
    port map (
            O => \N__21173\,
            I => \N__21019\
        );

    \I__4831\ : InMux
    port map (
            O => \N__21172\,
            I => \N__21019\
        );

    \I__4830\ : IoInMux
    port map (
            O => \N__21171\,
            I => \N__21016\
        );

    \I__4829\ : LocalMux
    port map (
            O => \N__21168\,
            I => \N__21013\
        );

    \I__4828\ : SRMux
    port map (
            O => \N__21167\,
            I => \N__21010\
        );

    \I__4827\ : SRMux
    port map (
            O => \N__21166\,
            I => \N__21007\
        );

    \I__4826\ : LocalMux
    port map (
            O => \N__21163\,
            I => \N__21000\
        );

    \I__4825\ : Span4Mux_h
    port map (
            O => \N__21158\,
            I => \N__21000\
        );

    \I__4824\ : LocalMux
    port map (
            O => \N__21155\,
            I => \N__21000\
        );

    \I__4823\ : LocalMux
    port map (
            O => \N__21152\,
            I => \N__20997\
        );

    \I__4822\ : SRMux
    port map (
            O => \N__21151\,
            I => \N__20994\
        );

    \I__4821\ : LocalMux
    port map (
            O => \N__21148\,
            I => \N__20991\
        );

    \I__4820\ : SRMux
    port map (
            O => \N__21147\,
            I => \N__20988\
        );

    \I__4819\ : LocalMux
    port map (
            O => \N__21144\,
            I => \N__20985\
        );

    \I__4818\ : Span4Mux_h
    port map (
            O => \N__21141\,
            I => \N__20976\
        );

    \I__4817\ : LocalMux
    port map (
            O => \N__21138\,
            I => \N__20976\
        );

    \I__4816\ : LocalMux
    port map (
            O => \N__21135\,
            I => \N__20976\
        );

    \I__4815\ : LocalMux
    port map (
            O => \N__21132\,
            I => \N__20976\
        );

    \I__4814\ : InMux
    port map (
            O => \N__21129\,
            I => \N__20973\
        );

    \I__4813\ : Span4Mux_v
    port map (
            O => \N__21124\,
            I => \N__20970\
        );

    \I__4812\ : LocalMux
    port map (
            O => \N__21121\,
            I => \N__20959\
        );

    \I__4811\ : LocalMux
    port map (
            O => \N__21118\,
            I => \N__20959\
        );

    \I__4810\ : Span4Mux_h
    port map (
            O => \N__21115\,
            I => \N__20959\
        );

    \I__4809\ : Span4Mux_h
    port map (
            O => \N__21108\,
            I => \N__20959\
        );

    \I__4808\ : Span4Mux_h
    port map (
            O => \N__21097\,
            I => \N__20959\
        );

    \I__4807\ : InMux
    port map (
            O => \N__21094\,
            I => \N__20956\
        );

    \I__4806\ : SRMux
    port map (
            O => \N__21093\,
            I => \N__20952\
        );

    \I__4805\ : SRMux
    port map (
            O => \N__21092\,
            I => \N__20949\
        );

    \I__4804\ : LocalMux
    port map (
            O => \N__21087\,
            I => \N__20946\
        );

    \I__4803\ : Span4Mux_h
    port map (
            O => \N__21084\,
            I => \N__20937\
        );

    \I__4802\ : Span4Mux_h
    port map (
            O => \N__21081\,
            I => \N__20937\
        );

    \I__4801\ : LocalMux
    port map (
            O => \N__21078\,
            I => \N__20937\
        );

    \I__4800\ : LocalMux
    port map (
            O => \N__21063\,
            I => \N__20937\
        );

    \I__4799\ : InMux
    port map (
            O => \N__21060\,
            I => \N__20932\
        );

    \I__4798\ : InMux
    port map (
            O => \N__21057\,
            I => \N__20932\
        );

    \I__4797\ : SRMux
    port map (
            O => \N__21056\,
            I => \N__20929\
        );

    \I__4796\ : SRMux
    port map (
            O => \N__21055\,
            I => \N__20926\
        );

    \I__4795\ : InMux
    port map (
            O => \N__21052\,
            I => \N__20923\
        );

    \I__4794\ : Span4Mux_v
    port map (
            O => \N__21049\,
            I => \N__20920\
        );

    \I__4793\ : Span4Mux_h
    port map (
            O => \N__21046\,
            I => \N__20915\
        );

    \I__4792\ : Span4Mux_v
    port map (
            O => \N__21041\,
            I => \N__20915\
        );

    \I__4791\ : LocalMux
    port map (
            O => \N__21038\,
            I => \N__20912\
        );

    \I__4790\ : InMux
    port map (
            O => \N__21037\,
            I => \N__20909\
        );

    \I__4789\ : InMux
    port map (
            O => \N__21036\,
            I => \N__20906\
        );

    \I__4788\ : InMux
    port map (
            O => \N__21035\,
            I => \N__20903\
        );

    \I__4787\ : InMux
    port map (
            O => \N__21034\,
            I => \N__20896\
        );

    \I__4786\ : InMux
    port map (
            O => \N__21033\,
            I => \N__20896\
        );

    \I__4785\ : InMux
    port map (
            O => \N__21030\,
            I => \N__20896\
        );

    \I__4784\ : LocalMux
    port map (
            O => \N__21027\,
            I => \N__20889\
        );

    \I__4783\ : LocalMux
    port map (
            O => \N__21024\,
            I => \N__20889\
        );

    \I__4782\ : LocalMux
    port map (
            O => \N__21019\,
            I => \N__20889\
        );

    \I__4781\ : LocalMux
    port map (
            O => \N__21016\,
            I => \N__20886\
        );

    \I__4780\ : Span4Mux_h
    port map (
            O => \N__21013\,
            I => \N__20881\
        );

    \I__4779\ : LocalMux
    port map (
            O => \N__21010\,
            I => \N__20881\
        );

    \I__4778\ : LocalMux
    port map (
            O => \N__21007\,
            I => \N__20874\
        );

    \I__4777\ : Sp12to4
    port map (
            O => \N__21000\,
            I => \N__20874\
        );

    \I__4776\ : Sp12to4
    port map (
            O => \N__20997\,
            I => \N__20874\
        );

    \I__4775\ : LocalMux
    port map (
            O => \N__20994\,
            I => \N__20871\
        );

    \I__4774\ : Span4Mux_h
    port map (
            O => \N__20991\,
            I => \N__20862\
        );

    \I__4773\ : LocalMux
    port map (
            O => \N__20988\,
            I => \N__20862\
        );

    \I__4772\ : Span4Mux_v
    port map (
            O => \N__20985\,
            I => \N__20862\
        );

    \I__4771\ : Span4Mux_v
    port map (
            O => \N__20976\,
            I => \N__20862\
        );

    \I__4770\ : LocalMux
    port map (
            O => \N__20973\,
            I => \N__20853\
        );

    \I__4769\ : Span4Mux_h
    port map (
            O => \N__20970\,
            I => \N__20853\
        );

    \I__4768\ : Span4Mux_v
    port map (
            O => \N__20959\,
            I => \N__20853\
        );

    \I__4767\ : LocalMux
    port map (
            O => \N__20956\,
            I => \N__20853\
        );

    \I__4766\ : SRMux
    port map (
            O => \N__20955\,
            I => \N__20850\
        );

    \I__4765\ : LocalMux
    port map (
            O => \N__20952\,
            I => \N__20845\
        );

    \I__4764\ : LocalMux
    port map (
            O => \N__20949\,
            I => \N__20845\
        );

    \I__4763\ : Span4Mux_h
    port map (
            O => \N__20946\,
            I => \N__20838\
        );

    \I__4762\ : Span4Mux_v
    port map (
            O => \N__20937\,
            I => \N__20838\
        );

    \I__4761\ : LocalMux
    port map (
            O => \N__20932\,
            I => \N__20838\
        );

    \I__4760\ : LocalMux
    port map (
            O => \N__20929\,
            I => \N__20835\
        );

    \I__4759\ : LocalMux
    port map (
            O => \N__20926\,
            I => \N__20832\
        );

    \I__4758\ : LocalMux
    port map (
            O => \N__20923\,
            I => \N__20829\
        );

    \I__4757\ : Span4Mux_h
    port map (
            O => \N__20920\,
            I => \N__20824\
        );

    \I__4756\ : Span4Mux_v
    port map (
            O => \N__20915\,
            I => \N__20824\
        );

    \I__4755\ : Span4Mux_v
    port map (
            O => \N__20912\,
            I => \N__20811\
        );

    \I__4754\ : LocalMux
    port map (
            O => \N__20909\,
            I => \N__20811\
        );

    \I__4753\ : LocalMux
    port map (
            O => \N__20906\,
            I => \N__20811\
        );

    \I__4752\ : LocalMux
    port map (
            O => \N__20903\,
            I => \N__20811\
        );

    \I__4751\ : LocalMux
    port map (
            O => \N__20896\,
            I => \N__20811\
        );

    \I__4750\ : Span4Mux_h
    port map (
            O => \N__20889\,
            I => \N__20811\
        );

    \I__4749\ : Span12Mux_s10_h
    port map (
            O => \N__20886\,
            I => \N__20808\
        );

    \I__4748\ : Span4Mux_v
    port map (
            O => \N__20881\,
            I => \N__20805\
        );

    \I__4747\ : Span12Mux_v
    port map (
            O => \N__20874\,
            I => \N__20802\
        );

    \I__4746\ : Span4Mux_v
    port map (
            O => \N__20871\,
            I => \N__20797\
        );

    \I__4745\ : Span4Mux_h
    port map (
            O => \N__20862\,
            I => \N__20797\
        );

    \I__4744\ : Span4Mux_h
    port map (
            O => \N__20853\,
            I => \N__20794\
        );

    \I__4743\ : LocalMux
    port map (
            O => \N__20850\,
            I => \N__20787\
        );

    \I__4742\ : Span4Mux_v
    port map (
            O => \N__20845\,
            I => \N__20787\
        );

    \I__4741\ : Span4Mux_h
    port map (
            O => \N__20838\,
            I => \N__20787\
        );

    \I__4740\ : Span4Mux_h
    port map (
            O => \N__20835\,
            I => \N__20776\
        );

    \I__4739\ : Span4Mux_h
    port map (
            O => \N__20832\,
            I => \N__20776\
        );

    \I__4738\ : Span4Mux_h
    port map (
            O => \N__20829\,
            I => \N__20776\
        );

    \I__4737\ : Span4Mux_v
    port map (
            O => \N__20824\,
            I => \N__20776\
        );

    \I__4736\ : Span4Mux_h
    port map (
            O => \N__20811\,
            I => \N__20776\
        );

    \I__4735\ : Odrv12
    port map (
            O => \N__20808\,
            I => \ADV_VSYNC_c\
        );

    \I__4734\ : Odrv4
    port map (
            O => \N__20805\,
            I => \ADV_VSYNC_c\
        );

    \I__4733\ : Odrv12
    port map (
            O => \N__20802\,
            I => \ADV_VSYNC_c\
        );

    \I__4732\ : Odrv4
    port map (
            O => \N__20797\,
            I => \ADV_VSYNC_c\
        );

    \I__4731\ : Odrv4
    port map (
            O => \N__20794\,
            I => \ADV_VSYNC_c\
        );

    \I__4730\ : Odrv4
    port map (
            O => \N__20787\,
            I => \ADV_VSYNC_c\
        );

    \I__4729\ : Odrv4
    port map (
            O => \N__20776\,
            I => \ADV_VSYNC_c\
        );

    \I__4728\ : InMux
    port map (
            O => \N__20761\,
            I => \N__20758\
        );

    \I__4727\ : LocalMux
    port map (
            O => \N__20758\,
            I => \N__20755\
        );

    \I__4726\ : Span12Mux_h
    port map (
            O => \N__20755\,
            I => \N__20752\
        );

    \I__4725\ : Span12Mux_v
    port map (
            O => \N__20752\,
            I => \N__20749\
        );

    \I__4724\ : Odrv12
    port map (
            O => \N__20749\,
            I => \line_buffer.n617\
        );

    \I__4723\ : CascadeMux
    port map (
            O => \N__20746\,
            I => \N__20743\
        );

    \I__4722\ : InMux
    port map (
            O => \N__20743\,
            I => \N__20740\
        );

    \I__4721\ : LocalMux
    port map (
            O => \N__20740\,
            I => \N__20737\
        );

    \I__4720\ : Span4Mux_h
    port map (
            O => \N__20737\,
            I => \N__20734\
        );

    \I__4719\ : Span4Mux_h
    port map (
            O => \N__20734\,
            I => \N__20731\
        );

    \I__4718\ : Span4Mux_v
    port map (
            O => \N__20731\,
            I => \N__20728\
        );

    \I__4717\ : Odrv4
    port map (
            O => \N__20728\,
            I => \line_buffer.n609\
        );

    \I__4716\ : InMux
    port map (
            O => \N__20725\,
            I => \N__20722\
        );

    \I__4715\ : LocalMux
    port map (
            O => \N__20722\,
            I => \N__20719\
        );

    \I__4714\ : Span4Mux_h
    port map (
            O => \N__20719\,
            I => \N__20716\
        );

    \I__4713\ : Span4Mux_h
    port map (
            O => \N__20716\,
            I => \N__20713\
        );

    \I__4712\ : Span4Mux_v
    port map (
            O => \N__20713\,
            I => \N__20710\
        );

    \I__4711\ : Odrv4
    port map (
            O => \N__20710\,
            I => \line_buffer.n610\
        );

    \I__4710\ : CascadeMux
    port map (
            O => \N__20707\,
            I => \N__20704\
        );

    \I__4709\ : InMux
    port map (
            O => \N__20704\,
            I => \N__20701\
        );

    \I__4708\ : LocalMux
    port map (
            O => \N__20701\,
            I => \N__20698\
        );

    \I__4707\ : Span4Mux_v
    port map (
            O => \N__20698\,
            I => \N__20695\
        );

    \I__4706\ : Sp12to4
    port map (
            O => \N__20695\,
            I => \N__20692\
        );

    \I__4705\ : Span12Mux_h
    port map (
            O => \N__20692\,
            I => \N__20689\
        );

    \I__4704\ : Span12Mux_v
    port map (
            O => \N__20689\,
            I => \N__20686\
        );

    \I__4703\ : Odrv12
    port map (
            O => \N__20686\,
            I => \line_buffer.n618\
        );

    \I__4702\ : InMux
    port map (
            O => \N__20683\,
            I => \N__20680\
        );

    \I__4701\ : LocalMux
    port map (
            O => \N__20680\,
            I => \line_buffer.n4161\
        );

    \I__4700\ : InMux
    port map (
            O => \N__20677\,
            I => \N__20674\
        );

    \I__4699\ : LocalMux
    port map (
            O => \N__20674\,
            I => \N__20671\
        );

    \I__4698\ : Odrv4
    port map (
            O => \N__20671\,
            I => \transmit_module.Y_DELTA_PATTERN_17\
        );

    \I__4697\ : InMux
    port map (
            O => \N__20668\,
            I => \N__20665\
        );

    \I__4696\ : LocalMux
    port map (
            O => \N__20665\,
            I => \transmit_module.Y_DELTA_PATTERN_16\
        );

    \I__4695\ : InMux
    port map (
            O => \N__20662\,
            I => \N__20659\
        );

    \I__4694\ : LocalMux
    port map (
            O => \N__20659\,
            I => \transmit_module.Y_DELTA_PATTERN_3\
        );

    \I__4693\ : InMux
    port map (
            O => \N__20656\,
            I => \N__20653\
        );

    \I__4692\ : LocalMux
    port map (
            O => \N__20653\,
            I => \N__20650\
        );

    \I__4691\ : Odrv4
    port map (
            O => \N__20650\,
            I => \transmit_module.Y_DELTA_PATTERN_2\
        );

    \I__4690\ : InMux
    port map (
            O => \N__20647\,
            I => \N__20644\
        );

    \I__4689\ : LocalMux
    port map (
            O => \N__20644\,
            I => \N__20641\
        );

    \I__4688\ : Span4Mux_h
    port map (
            O => \N__20641\,
            I => \N__20638\
        );

    \I__4687\ : Odrv4
    port map (
            O => \N__20638\,
            I => \transmit_module.Y_DELTA_PATTERN_22\
        );

    \I__4686\ : InMux
    port map (
            O => \N__20635\,
            I => \N__20632\
        );

    \I__4685\ : LocalMux
    port map (
            O => \N__20632\,
            I => \transmit_module.Y_DELTA_PATTERN_24\
        );

    \I__4684\ : InMux
    port map (
            O => \N__20629\,
            I => \N__20626\
        );

    \I__4683\ : LocalMux
    port map (
            O => \N__20626\,
            I => \transmit_module.Y_DELTA_PATTERN_23\
        );

    \I__4682\ : CEMux
    port map (
            O => \N__20623\,
            I => \N__20619\
        );

    \I__4681\ : CEMux
    port map (
            O => \N__20622\,
            I => \N__20615\
        );

    \I__4680\ : LocalMux
    port map (
            O => \N__20619\,
            I => \N__20611\
        );

    \I__4679\ : CEMux
    port map (
            O => \N__20618\,
            I => \N__20608\
        );

    \I__4678\ : LocalMux
    port map (
            O => \N__20615\,
            I => \N__20603\
        );

    \I__4677\ : CEMux
    port map (
            O => \N__20614\,
            I => \N__20600\
        );

    \I__4676\ : Span4Mux_v
    port map (
            O => \N__20611\,
            I => \N__20591\
        );

    \I__4675\ : LocalMux
    port map (
            O => \N__20608\,
            I => \N__20591\
        );

    \I__4674\ : CEMux
    port map (
            O => \N__20607\,
            I => \N__20588\
        );

    \I__4673\ : CEMux
    port map (
            O => \N__20606\,
            I => \N__20584\
        );

    \I__4672\ : Span4Mux_h
    port map (
            O => \N__20603\,
            I => \N__20578\
        );

    \I__4671\ : LocalMux
    port map (
            O => \N__20600\,
            I => \N__20578\
        );

    \I__4670\ : CEMux
    port map (
            O => \N__20599\,
            I => \N__20575\
        );

    \I__4669\ : CEMux
    port map (
            O => \N__20598\,
            I => \N__20572\
        );

    \I__4668\ : CEMux
    port map (
            O => \N__20597\,
            I => \N__20569\
        );

    \I__4667\ : CEMux
    port map (
            O => \N__20596\,
            I => \N__20566\
        );

    \I__4666\ : Span4Mux_h
    port map (
            O => \N__20591\,
            I => \N__20560\
        );

    \I__4665\ : LocalMux
    port map (
            O => \N__20588\,
            I => \N__20560\
        );

    \I__4664\ : SRMux
    port map (
            O => \N__20587\,
            I => \N__20557\
        );

    \I__4663\ : LocalMux
    port map (
            O => \N__20584\,
            I => \N__20554\
        );

    \I__4662\ : SRMux
    port map (
            O => \N__20583\,
            I => \N__20551\
        );

    \I__4661\ : Span4Mux_v
    port map (
            O => \N__20578\,
            I => \N__20547\
        );

    \I__4660\ : LocalMux
    port map (
            O => \N__20575\,
            I => \N__20542\
        );

    \I__4659\ : LocalMux
    port map (
            O => \N__20572\,
            I => \N__20542\
        );

    \I__4658\ : LocalMux
    port map (
            O => \N__20569\,
            I => \N__20539\
        );

    \I__4657\ : LocalMux
    port map (
            O => \N__20566\,
            I => \N__20536\
        );

    \I__4656\ : SRMux
    port map (
            O => \N__20565\,
            I => \N__20533\
        );

    \I__4655\ : Span4Mux_v
    port map (
            O => \N__20560\,
            I => \N__20530\
        );

    \I__4654\ : LocalMux
    port map (
            O => \N__20557\,
            I => \N__20527\
        );

    \I__4653\ : Span4Mux_v
    port map (
            O => \N__20554\,
            I => \N__20522\
        );

    \I__4652\ : LocalMux
    port map (
            O => \N__20551\,
            I => \N__20522\
        );

    \I__4651\ : SRMux
    port map (
            O => \N__20550\,
            I => \N__20519\
        );

    \I__4650\ : Span4Mux_h
    port map (
            O => \N__20547\,
            I => \N__20514\
        );

    \I__4649\ : Span4Mux_v
    port map (
            O => \N__20542\,
            I => \N__20514\
        );

    \I__4648\ : Span4Mux_v
    port map (
            O => \N__20539\,
            I => \N__20511\
        );

    \I__4647\ : Sp12to4
    port map (
            O => \N__20536\,
            I => \N__20508\
        );

    \I__4646\ : LocalMux
    port map (
            O => \N__20533\,
            I => \N__20505\
        );

    \I__4645\ : Span4Mux_h
    port map (
            O => \N__20530\,
            I => \N__20496\
        );

    \I__4644\ : Span4Mux_v
    port map (
            O => \N__20527\,
            I => \N__20496\
        );

    \I__4643\ : Span4Mux_h
    port map (
            O => \N__20522\,
            I => \N__20496\
        );

    \I__4642\ : LocalMux
    port map (
            O => \N__20519\,
            I => \N__20496\
        );

    \I__4641\ : Odrv4
    port map (
            O => \N__20514\,
            I => \transmit_module.n4224\
        );

    \I__4640\ : Odrv4
    port map (
            O => \N__20511\,
            I => \transmit_module.n4224\
        );

    \I__4639\ : Odrv12
    port map (
            O => \N__20508\,
            I => \transmit_module.n4224\
        );

    \I__4638\ : Odrv12
    port map (
            O => \N__20505\,
            I => \transmit_module.n4224\
        );

    \I__4637\ : Odrv4
    port map (
            O => \N__20496\,
            I => \transmit_module.n4224\
        );

    \I__4636\ : InMux
    port map (
            O => \N__20485\,
            I => \N__20482\
        );

    \I__4635\ : LocalMux
    port map (
            O => \N__20482\,
            I => \N__20479\
        );

    \I__4634\ : Span4Mux_v
    port map (
            O => \N__20479\,
            I => \N__20476\
        );

    \I__4633\ : Span4Mux_h
    port map (
            O => \N__20476\,
            I => \N__20473\
        );

    \I__4632\ : Odrv4
    port map (
            O => \N__20473\,
            I => \line_buffer.n642\
        );

    \I__4631\ : CascadeMux
    port map (
            O => \N__20470\,
            I => \N__20467\
        );

    \I__4630\ : InMux
    port map (
            O => \N__20467\,
            I => \N__20464\
        );

    \I__4629\ : LocalMux
    port map (
            O => \N__20464\,
            I => \N__20461\
        );

    \I__4628\ : Span4Mux_v
    port map (
            O => \N__20461\,
            I => \N__20458\
        );

    \I__4627\ : Span4Mux_v
    port map (
            O => \N__20458\,
            I => \N__20455\
        );

    \I__4626\ : Sp12to4
    port map (
            O => \N__20455\,
            I => \N__20452\
        );

    \I__4625\ : Odrv12
    port map (
            O => \N__20452\,
            I => \line_buffer.n650\
        );

    \I__4624\ : InMux
    port map (
            O => \N__20449\,
            I => \N__20446\
        );

    \I__4623\ : LocalMux
    port map (
            O => \N__20446\,
            I => \N__20443\
        );

    \I__4622\ : Span4Mux_v
    port map (
            O => \N__20443\,
            I => \N__20440\
        );

    \I__4621\ : Sp12to4
    port map (
            O => \N__20440\,
            I => \N__20437\
        );

    \I__4620\ : Span12Mux_h
    port map (
            O => \N__20437\,
            I => \N__20434\
        );

    \I__4619\ : Span12Mux_v
    port map (
            O => \N__20434\,
            I => \N__20431\
        );

    \I__4618\ : Odrv12
    port map (
            O => \N__20431\,
            I => \line_buffer.n545\
        );

    \I__4617\ : CascadeMux
    port map (
            O => \N__20428\,
            I => \line_buffer.n4164_cascade_\
        );

    \I__4616\ : InMux
    port map (
            O => \N__20425\,
            I => \N__20422\
        );

    \I__4615\ : LocalMux
    port map (
            O => \N__20422\,
            I => \N__20419\
        );

    \I__4614\ : Span4Mux_h
    port map (
            O => \N__20419\,
            I => \N__20416\
        );

    \I__4613\ : Span4Mux_v
    port map (
            O => \N__20416\,
            I => \N__20413\
        );

    \I__4612\ : Span4Mux_h
    port map (
            O => \N__20413\,
            I => \N__20410\
        );

    \I__4611\ : Odrv4
    port map (
            O => \N__20410\,
            I => \line_buffer.n553\
        );

    \I__4610\ : CascadeMux
    port map (
            O => \N__20407\,
            I => \line_buffer.n4167_cascade_\
        );

    \I__4609\ : InMux
    port map (
            O => \N__20404\,
            I => \N__20401\
        );

    \I__4608\ : LocalMux
    port map (
            O => \N__20401\,
            I => \N__20398\
        );

    \I__4607\ : Span4Mux_h
    port map (
            O => \N__20398\,
            I => \N__20395\
        );

    \I__4606\ : Span4Mux_h
    port map (
            O => \N__20395\,
            I => \N__20392\
        );

    \I__4605\ : Odrv4
    port map (
            O => \N__20392\,
            I => \TX_DATA_1\
        );

    \I__4604\ : InMux
    port map (
            O => \N__20389\,
            I => \N__20386\
        );

    \I__4603\ : LocalMux
    port map (
            O => \N__20386\,
            I => \N__20383\
        );

    \I__4602\ : Span12Mux_v
    port map (
            O => \N__20383\,
            I => \N__20380\
        );

    \I__4601\ : Odrv12
    port map (
            O => \N__20380\,
            I => \line_buffer.n4065\
        );

    \I__4600\ : InMux
    port map (
            O => \N__20377\,
            I => \N__20374\
        );

    \I__4599\ : LocalMux
    port map (
            O => \N__20374\,
            I => \N__20371\
        );

    \I__4598\ : Span4Mux_v
    port map (
            O => \N__20371\,
            I => \N__20368\
        );

    \I__4597\ : Span4Mux_v
    port map (
            O => \N__20368\,
            I => \N__20365\
        );

    \I__4596\ : Sp12to4
    port map (
            O => \N__20365\,
            I => \N__20362\
        );

    \I__4595\ : Odrv12
    port map (
            O => \N__20362\,
            I => \line_buffer.n620\
        );

    \I__4594\ : InMux
    port map (
            O => \N__20359\,
            I => \N__20356\
        );

    \I__4593\ : LocalMux
    port map (
            O => \N__20356\,
            I => \N__20353\
        );

    \I__4592\ : Odrv12
    port map (
            O => \N__20353\,
            I => \line_buffer.n612\
        );

    \I__4591\ : InMux
    port map (
            O => \N__20350\,
            I => \N__20347\
        );

    \I__4590\ : LocalMux
    port map (
            O => \N__20347\,
            I => \transmit_module.Y_DELTA_PATTERN_6\
        );

    \I__4589\ : InMux
    port map (
            O => \N__20344\,
            I => \N__20341\
        );

    \I__4588\ : LocalMux
    port map (
            O => \N__20341\,
            I => \transmit_module.Y_DELTA_PATTERN_5\
        );

    \I__4587\ : InMux
    port map (
            O => \N__20338\,
            I => \N__20335\
        );

    \I__4586\ : LocalMux
    port map (
            O => \N__20335\,
            I => \transmit_module.Y_DELTA_PATTERN_7\
        );

    \I__4585\ : InMux
    port map (
            O => \N__20332\,
            I => \N__20329\
        );

    \I__4584\ : LocalMux
    port map (
            O => \N__20329\,
            I => \transmit_module.Y_DELTA_PATTERN_11\
        );

    \I__4583\ : InMux
    port map (
            O => \N__20326\,
            I => \N__20323\
        );

    \I__4582\ : LocalMux
    port map (
            O => \N__20323\,
            I => \transmit_module.Y_DELTA_PATTERN_10\
        );

    \I__4581\ : InMux
    port map (
            O => \N__20320\,
            I => \N__20317\
        );

    \I__4580\ : LocalMux
    port map (
            O => \N__20317\,
            I => \transmit_module.Y_DELTA_PATTERN_9\
        );

    \I__4579\ : InMux
    port map (
            O => \N__20314\,
            I => \N__20311\
        );

    \I__4578\ : LocalMux
    port map (
            O => \N__20311\,
            I => \transmit_module.Y_DELTA_PATTERN_8\
        );

    \I__4577\ : InMux
    port map (
            O => \N__20308\,
            I => \N__20305\
        );

    \I__4576\ : LocalMux
    port map (
            O => \N__20305\,
            I => \transmit_module.Y_DELTA_PATTERN_15\
        );

    \I__4575\ : InMux
    port map (
            O => \N__20302\,
            I => \N__20299\
        );

    \I__4574\ : LocalMux
    port map (
            O => \N__20299\,
            I => \N__20296\
        );

    \I__4573\ : Odrv4
    port map (
            O => \N__20296\,
            I => \transmit_module.Y_DELTA_PATTERN_4\
        );

    \I__4572\ : InMux
    port map (
            O => \N__20293\,
            I => \N__20290\
        );

    \I__4571\ : LocalMux
    port map (
            O => \N__20290\,
            I => \transmit_module.Y_DELTA_PATTERN_37\
        );

    \I__4570\ : InMux
    port map (
            O => \N__20287\,
            I => \N__20284\
        );

    \I__4569\ : LocalMux
    port map (
            O => \N__20284\,
            I => \transmit_module.Y_DELTA_PATTERN_36\
        );

    \I__4568\ : InMux
    port map (
            O => \N__20281\,
            I => \N__20278\
        );

    \I__4567\ : LocalMux
    port map (
            O => \N__20278\,
            I => \transmit_module.Y_DELTA_PATTERN_38\
        );

    \I__4566\ : InMux
    port map (
            O => \N__20275\,
            I => \N__20271\
        );

    \I__4565\ : InMux
    port map (
            O => \N__20274\,
            I => \N__20268\
        );

    \I__4564\ : LocalMux
    port map (
            O => \N__20271\,
            I => \N__20265\
        );

    \I__4563\ : LocalMux
    port map (
            O => \N__20268\,
            I => \transmit_module.n185\
        );

    \I__4562\ : Odrv4
    port map (
            O => \N__20265\,
            I => \transmit_module.n185\
        );

    \I__4561\ : InMux
    port map (
            O => \N__20260\,
            I => \N__20256\
        );

    \I__4560\ : InMux
    port map (
            O => \N__20259\,
            I => \N__20253\
        );

    \I__4559\ : LocalMux
    port map (
            O => \N__20256\,
            I => \N__20250\
        );

    \I__4558\ : LocalMux
    port map (
            O => \N__20253\,
            I => \transmit_module.n216\
        );

    \I__4557\ : Odrv12
    port map (
            O => \N__20250\,
            I => \transmit_module.n216\
        );

    \I__4556\ : InMux
    port map (
            O => \N__20245\,
            I => \N__20242\
        );

    \I__4555\ : LocalMux
    port map (
            O => \N__20242\,
            I => \N__20236\
        );

    \I__4554\ : InMux
    port map (
            O => \N__20241\,
            I => \N__20233\
        );

    \I__4553\ : InMux
    port map (
            O => \N__20240\,
            I => \N__20230\
        );

    \I__4552\ : InMux
    port map (
            O => \N__20239\,
            I => \N__20225\
        );

    \I__4551\ : Span4Mux_h
    port map (
            O => \N__20236\,
            I => \N__20220\
        );

    \I__4550\ : LocalMux
    port map (
            O => \N__20233\,
            I => \N__20220\
        );

    \I__4549\ : LocalMux
    port map (
            O => \N__20230\,
            I => \N__20217\
        );

    \I__4548\ : InMux
    port map (
            O => \N__20229\,
            I => \N__20210\
        );

    \I__4547\ : InMux
    port map (
            O => \N__20228\,
            I => \N__20210\
        );

    \I__4546\ : LocalMux
    port map (
            O => \N__20225\,
            I => \N__20202\
        );

    \I__4545\ : Span4Mux_v
    port map (
            O => \N__20220\,
            I => \N__20202\
        );

    \I__4544\ : Span4Mux_h
    port map (
            O => \N__20217\,
            I => \N__20202\
        );

    \I__4543\ : InMux
    port map (
            O => \N__20216\,
            I => \N__20199\
        );

    \I__4542\ : InMux
    port map (
            O => \N__20215\,
            I => \N__20188\
        );

    \I__4541\ : LocalMux
    port map (
            O => \N__20210\,
            I => \N__20185\
        );

    \I__4540\ : InMux
    port map (
            O => \N__20209\,
            I => \N__20182\
        );

    \I__4539\ : Span4Mux_v
    port map (
            O => \N__20202\,
            I => \N__20179\
        );

    \I__4538\ : LocalMux
    port map (
            O => \N__20199\,
            I => \N__20176\
        );

    \I__4537\ : InMux
    port map (
            O => \N__20198\,
            I => \N__20171\
        );

    \I__4536\ : InMux
    port map (
            O => \N__20197\,
            I => \N__20171\
        );

    \I__4535\ : InMux
    port map (
            O => \N__20196\,
            I => \N__20153\
        );

    \I__4534\ : InMux
    port map (
            O => \N__20195\,
            I => \N__20153\
        );

    \I__4533\ : InMux
    port map (
            O => \N__20194\,
            I => \N__20153\
        );

    \I__4532\ : InMux
    port map (
            O => \N__20193\,
            I => \N__20153\
        );

    \I__4531\ : InMux
    port map (
            O => \N__20192\,
            I => \N__20153\
        );

    \I__4530\ : InMux
    port map (
            O => \N__20191\,
            I => \N__20153\
        );

    \I__4529\ : LocalMux
    port map (
            O => \N__20188\,
            I => \N__20150\
        );

    \I__4528\ : Span4Mux_v
    port map (
            O => \N__20185\,
            I => \N__20139\
        );

    \I__4527\ : LocalMux
    port map (
            O => \N__20182\,
            I => \N__20139\
        );

    \I__4526\ : Span4Mux_v
    port map (
            O => \N__20179\,
            I => \N__20139\
        );

    \I__4525\ : Span4Mux_h
    port map (
            O => \N__20176\,
            I => \N__20139\
        );

    \I__4524\ : LocalMux
    port map (
            O => \N__20171\,
            I => \N__20139\
        );

    \I__4523\ : InMux
    port map (
            O => \N__20170\,
            I => \N__20132\
        );

    \I__4522\ : InMux
    port map (
            O => \N__20169\,
            I => \N__20132\
        );

    \I__4521\ : InMux
    port map (
            O => \N__20168\,
            I => \N__20132\
        );

    \I__4520\ : InMux
    port map (
            O => \N__20167\,
            I => \N__20127\
        );

    \I__4519\ : InMux
    port map (
            O => \N__20166\,
            I => \N__20127\
        );

    \I__4518\ : LocalMux
    port map (
            O => \N__20153\,
            I => \transmit_module.n4211\
        );

    \I__4517\ : Odrv4
    port map (
            O => \N__20150\,
            I => \transmit_module.n4211\
        );

    \I__4516\ : Odrv4
    port map (
            O => \N__20139\,
            I => \transmit_module.n4211\
        );

    \I__4515\ : LocalMux
    port map (
            O => \N__20132\,
            I => \transmit_module.n4211\
        );

    \I__4514\ : LocalMux
    port map (
            O => \N__20127\,
            I => \transmit_module.n4211\
        );

    \I__4513\ : CascadeMux
    port map (
            O => \N__20116\,
            I => \N__20112\
        );

    \I__4512\ : CascadeMux
    port map (
            O => \N__20115\,
            I => \N__20109\
        );

    \I__4511\ : CascadeBuf
    port map (
            O => \N__20112\,
            I => \N__20106\
        );

    \I__4510\ : CascadeBuf
    port map (
            O => \N__20109\,
            I => \N__20103\
        );

    \I__4509\ : CascadeMux
    port map (
            O => \N__20106\,
            I => \N__20100\
        );

    \I__4508\ : CascadeMux
    port map (
            O => \N__20103\,
            I => \N__20097\
        );

    \I__4507\ : CascadeBuf
    port map (
            O => \N__20100\,
            I => \N__20094\
        );

    \I__4506\ : CascadeBuf
    port map (
            O => \N__20097\,
            I => \N__20091\
        );

    \I__4505\ : CascadeMux
    port map (
            O => \N__20094\,
            I => \N__20088\
        );

    \I__4504\ : CascadeMux
    port map (
            O => \N__20091\,
            I => \N__20085\
        );

    \I__4503\ : CascadeBuf
    port map (
            O => \N__20088\,
            I => \N__20082\
        );

    \I__4502\ : CascadeBuf
    port map (
            O => \N__20085\,
            I => \N__20079\
        );

    \I__4501\ : CascadeMux
    port map (
            O => \N__20082\,
            I => \N__20076\
        );

    \I__4500\ : CascadeMux
    port map (
            O => \N__20079\,
            I => \N__20073\
        );

    \I__4499\ : CascadeBuf
    port map (
            O => \N__20076\,
            I => \N__20070\
        );

    \I__4498\ : CascadeBuf
    port map (
            O => \N__20073\,
            I => \N__20067\
        );

    \I__4497\ : CascadeMux
    port map (
            O => \N__20070\,
            I => \N__20064\
        );

    \I__4496\ : CascadeMux
    port map (
            O => \N__20067\,
            I => \N__20061\
        );

    \I__4495\ : CascadeBuf
    port map (
            O => \N__20064\,
            I => \N__20058\
        );

    \I__4494\ : CascadeBuf
    port map (
            O => \N__20061\,
            I => \N__20055\
        );

    \I__4493\ : CascadeMux
    port map (
            O => \N__20058\,
            I => \N__20052\
        );

    \I__4492\ : CascadeMux
    port map (
            O => \N__20055\,
            I => \N__20049\
        );

    \I__4491\ : CascadeBuf
    port map (
            O => \N__20052\,
            I => \N__20046\
        );

    \I__4490\ : CascadeBuf
    port map (
            O => \N__20049\,
            I => \N__20043\
        );

    \I__4489\ : CascadeMux
    port map (
            O => \N__20046\,
            I => \N__20040\
        );

    \I__4488\ : CascadeMux
    port map (
            O => \N__20043\,
            I => \N__20037\
        );

    \I__4487\ : CascadeBuf
    port map (
            O => \N__20040\,
            I => \N__20034\
        );

    \I__4486\ : CascadeBuf
    port map (
            O => \N__20037\,
            I => \N__20031\
        );

    \I__4485\ : CascadeMux
    port map (
            O => \N__20034\,
            I => \N__20028\
        );

    \I__4484\ : CascadeMux
    port map (
            O => \N__20031\,
            I => \N__20025\
        );

    \I__4483\ : CascadeBuf
    port map (
            O => \N__20028\,
            I => \N__20022\
        );

    \I__4482\ : CascadeBuf
    port map (
            O => \N__20025\,
            I => \N__20019\
        );

    \I__4481\ : CascadeMux
    port map (
            O => \N__20022\,
            I => \N__20016\
        );

    \I__4480\ : CascadeMux
    port map (
            O => \N__20019\,
            I => \N__20013\
        );

    \I__4479\ : CascadeBuf
    port map (
            O => \N__20016\,
            I => \N__20010\
        );

    \I__4478\ : CascadeBuf
    port map (
            O => \N__20013\,
            I => \N__20007\
        );

    \I__4477\ : CascadeMux
    port map (
            O => \N__20010\,
            I => \N__20004\
        );

    \I__4476\ : CascadeMux
    port map (
            O => \N__20007\,
            I => \N__20001\
        );

    \I__4475\ : CascadeBuf
    port map (
            O => \N__20004\,
            I => \N__19998\
        );

    \I__4474\ : CascadeBuf
    port map (
            O => \N__20001\,
            I => \N__19995\
        );

    \I__4473\ : CascadeMux
    port map (
            O => \N__19998\,
            I => \N__19992\
        );

    \I__4472\ : CascadeMux
    port map (
            O => \N__19995\,
            I => \N__19989\
        );

    \I__4471\ : CascadeBuf
    port map (
            O => \N__19992\,
            I => \N__19986\
        );

    \I__4470\ : CascadeBuf
    port map (
            O => \N__19989\,
            I => \N__19983\
        );

    \I__4469\ : CascadeMux
    port map (
            O => \N__19986\,
            I => \N__19980\
        );

    \I__4468\ : CascadeMux
    port map (
            O => \N__19983\,
            I => \N__19977\
        );

    \I__4467\ : CascadeBuf
    port map (
            O => \N__19980\,
            I => \N__19974\
        );

    \I__4466\ : CascadeBuf
    port map (
            O => \N__19977\,
            I => \N__19971\
        );

    \I__4465\ : CascadeMux
    port map (
            O => \N__19974\,
            I => \N__19968\
        );

    \I__4464\ : CascadeMux
    port map (
            O => \N__19971\,
            I => \N__19965\
        );

    \I__4463\ : CascadeBuf
    port map (
            O => \N__19968\,
            I => \N__19962\
        );

    \I__4462\ : CascadeBuf
    port map (
            O => \N__19965\,
            I => \N__19959\
        );

    \I__4461\ : CascadeMux
    port map (
            O => \N__19962\,
            I => \N__19956\
        );

    \I__4460\ : CascadeMux
    port map (
            O => \N__19959\,
            I => \N__19953\
        );

    \I__4459\ : CascadeBuf
    port map (
            O => \N__19956\,
            I => \N__19950\
        );

    \I__4458\ : CascadeBuf
    port map (
            O => \N__19953\,
            I => \N__19947\
        );

    \I__4457\ : CascadeMux
    port map (
            O => \N__19950\,
            I => \N__19944\
        );

    \I__4456\ : CascadeMux
    port map (
            O => \N__19947\,
            I => \N__19941\
        );

    \I__4455\ : CascadeBuf
    port map (
            O => \N__19944\,
            I => \N__19938\
        );

    \I__4454\ : CascadeBuf
    port map (
            O => \N__19941\,
            I => \N__19935\
        );

    \I__4453\ : CascadeMux
    port map (
            O => \N__19938\,
            I => \N__19932\
        );

    \I__4452\ : CascadeMux
    port map (
            O => \N__19935\,
            I => \N__19929\
        );

    \I__4451\ : InMux
    port map (
            O => \N__19932\,
            I => \N__19926\
        );

    \I__4450\ : InMux
    port map (
            O => \N__19929\,
            I => \N__19923\
        );

    \I__4449\ : LocalMux
    port map (
            O => \N__19926\,
            I => \N__19920\
        );

    \I__4448\ : LocalMux
    port map (
            O => \N__19923\,
            I => \N__19917\
        );

    \I__4447\ : Span12Mux_h
    port map (
            O => \N__19920\,
            I => \N__19912\
        );

    \I__4446\ : Span12Mux_h
    port map (
            O => \N__19917\,
            I => \N__19912\
        );

    \I__4445\ : Span12Mux_v
    port map (
            O => \N__19912\,
            I => \N__19909\
        );

    \I__4444\ : Odrv12
    port map (
            O => \N__19909\,
            I => n25
        );

    \I__4443\ : CascadeMux
    port map (
            O => \N__19906\,
            I => \N__19903\
        );

    \I__4442\ : InMux
    port map (
            O => \N__19903\,
            I => \N__19900\
        );

    \I__4441\ : LocalMux
    port map (
            O => \N__19900\,
            I => \transmit_module.ADDR_Y_COMPONENT_12\
        );

    \I__4440\ : CascadeMux
    port map (
            O => \N__19897\,
            I => \N__19894\
        );

    \I__4439\ : InMux
    port map (
            O => \N__19894\,
            I => \N__19891\
        );

    \I__4438\ : LocalMux
    port map (
            O => \N__19891\,
            I => \N__19888\
        );

    \I__4437\ : Span4Mux_v
    port map (
            O => \N__19888\,
            I => \N__19885\
        );

    \I__4436\ : Odrv4
    port map (
            O => \N__19885\,
            I => \transmit_module.ADDR_Y_COMPONENT_13\
        );

    \I__4435\ : CEMux
    port map (
            O => \N__19882\,
            I => \N__19878\
        );

    \I__4434\ : CEMux
    port map (
            O => \N__19881\,
            I => \N__19871\
        );

    \I__4433\ : LocalMux
    port map (
            O => \N__19878\,
            I => \N__19866\
        );

    \I__4432\ : CEMux
    port map (
            O => \N__19877\,
            I => \N__19863\
        );

    \I__4431\ : CEMux
    port map (
            O => \N__19876\,
            I => \N__19860\
        );

    \I__4430\ : CEMux
    port map (
            O => \N__19875\,
            I => \N__19857\
        );

    \I__4429\ : CEMux
    port map (
            O => \N__19874\,
            I => \N__19854\
        );

    \I__4428\ : LocalMux
    port map (
            O => \N__19871\,
            I => \N__19850\
        );

    \I__4427\ : CEMux
    port map (
            O => \N__19870\,
            I => \N__19847\
        );

    \I__4426\ : CEMux
    port map (
            O => \N__19869\,
            I => \N__19844\
        );

    \I__4425\ : Span4Mux_v
    port map (
            O => \N__19866\,
            I => \N__19841\
        );

    \I__4424\ : LocalMux
    port map (
            O => \N__19863\,
            I => \N__19836\
        );

    \I__4423\ : LocalMux
    port map (
            O => \N__19860\,
            I => \N__19836\
        );

    \I__4422\ : LocalMux
    port map (
            O => \N__19857\,
            I => \N__19831\
        );

    \I__4421\ : LocalMux
    port map (
            O => \N__19854\,
            I => \N__19831\
        );

    \I__4420\ : CEMux
    port map (
            O => \N__19853\,
            I => \N__19828\
        );

    \I__4419\ : Span4Mux_h
    port map (
            O => \N__19850\,
            I => \N__19825\
        );

    \I__4418\ : LocalMux
    port map (
            O => \N__19847\,
            I => \N__19822\
        );

    \I__4417\ : LocalMux
    port map (
            O => \N__19844\,
            I => \N__19819\
        );

    \I__4416\ : Span4Mux_v
    port map (
            O => \N__19841\,
            I => \N__19814\
        );

    \I__4415\ : Span4Mux_h
    port map (
            O => \N__19836\,
            I => \N__19814\
        );

    \I__4414\ : Span4Mux_v
    port map (
            O => \N__19831\,
            I => \N__19809\
        );

    \I__4413\ : LocalMux
    port map (
            O => \N__19828\,
            I => \N__19809\
        );

    \I__4412\ : Span4Mux_v
    port map (
            O => \N__19825\,
            I => \N__19804\
        );

    \I__4411\ : Span4Mux_h
    port map (
            O => \N__19822\,
            I => \N__19804\
        );

    \I__4410\ : Span4Mux_h
    port map (
            O => \N__19819\,
            I => \N__19799\
        );

    \I__4409\ : Span4Mux_h
    port map (
            O => \N__19814\,
            I => \N__19799\
        );

    \I__4408\ : Span4Mux_h
    port map (
            O => \N__19809\,
            I => \N__19796\
        );

    \I__4407\ : Odrv4
    port map (
            O => \N__19804\,
            I => \transmit_module.n2305\
        );

    \I__4406\ : Odrv4
    port map (
            O => \N__19799\,
            I => \transmit_module.n2305\
        );

    \I__4405\ : Odrv4
    port map (
            O => \N__19796\,
            I => \transmit_module.n2305\
        );

    \I__4404\ : InMux
    port map (
            O => \N__19789\,
            I => \N__19786\
        );

    \I__4403\ : LocalMux
    port map (
            O => \N__19786\,
            I => \N__19783\
        );

    \I__4402\ : Odrv4
    port map (
            O => \N__19783\,
            I => \transmit_module.Y_DELTA_PATTERN_39\
        );

    \I__4401\ : InMux
    port map (
            O => \N__19780\,
            I => \N__19777\
        );

    \I__4400\ : LocalMux
    port map (
            O => \N__19777\,
            I => \transmit_module.Y_DELTA_PATTERN_41\
        );

    \I__4399\ : InMux
    port map (
            O => \N__19774\,
            I => \N__19771\
        );

    \I__4398\ : LocalMux
    port map (
            O => \N__19771\,
            I => \transmit_module.Y_DELTA_PATTERN_40\
        );

    \I__4397\ : InMux
    port map (
            O => \N__19768\,
            I => \N__19765\
        );

    \I__4396\ : LocalMux
    port map (
            O => \N__19765\,
            I => \transmit_module.Y_DELTA_PATTERN_12\
        );

    \I__4395\ : InMux
    port map (
            O => \N__19762\,
            I => \N__19759\
        );

    \I__4394\ : LocalMux
    port map (
            O => \N__19759\,
            I => \transmit_module.Y_DELTA_PATTERN_32\
        );

    \I__4393\ : InMux
    port map (
            O => \N__19756\,
            I => \N__19753\
        );

    \I__4392\ : LocalMux
    port map (
            O => \N__19753\,
            I => \transmit_module.Y_DELTA_PATTERN_13\
        );

    \I__4391\ : InMux
    port map (
            O => \N__19750\,
            I => \N__19747\
        );

    \I__4390\ : LocalMux
    port map (
            O => \N__19747\,
            I => \transmit_module.Y_DELTA_PATTERN_14\
        );

    \I__4389\ : InMux
    port map (
            O => \N__19744\,
            I => \N__19741\
        );

    \I__4388\ : LocalMux
    port map (
            O => \N__19741\,
            I => \transmit_module.Y_DELTA_PATTERN_26\
        );

    \I__4387\ : InMux
    port map (
            O => \N__19738\,
            I => \N__19735\
        );

    \I__4386\ : LocalMux
    port map (
            O => \N__19735\,
            I => \transmit_module.Y_DELTA_PATTERN_25\
        );

    \I__4385\ : InMux
    port map (
            O => \N__19732\,
            I => \N__19729\
        );

    \I__4384\ : LocalMux
    port map (
            O => \N__19729\,
            I => \N__19726\
        );

    \I__4383\ : Odrv4
    port map (
            O => \N__19726\,
            I => \transmit_module.Y_DELTA_PATTERN_28\
        );

    \I__4382\ : InMux
    port map (
            O => \N__19723\,
            I => \N__19720\
        );

    \I__4381\ : LocalMux
    port map (
            O => \N__19720\,
            I => \transmit_module.Y_DELTA_PATTERN_27\
        );

    \I__4380\ : InMux
    port map (
            O => \N__19717\,
            I => \N__19710\
        );

    \I__4379\ : InMux
    port map (
            O => \N__19716\,
            I => \N__19707\
        );

    \I__4378\ : InMux
    port map (
            O => \N__19715\,
            I => \N__19702\
        );

    \I__4377\ : InMux
    port map (
            O => \N__19714\,
            I => \N__19702\
        );

    \I__4376\ : InMux
    port map (
            O => \N__19713\,
            I => \N__19698\
        );

    \I__4375\ : LocalMux
    port map (
            O => \N__19710\,
            I => \N__19694\
        );

    \I__4374\ : LocalMux
    port map (
            O => \N__19707\,
            I => \N__19686\
        );

    \I__4373\ : LocalMux
    port map (
            O => \N__19702\,
            I => \N__19686\
        );

    \I__4372\ : InMux
    port map (
            O => \N__19701\,
            I => \N__19683\
        );

    \I__4371\ : LocalMux
    port map (
            O => \N__19698\,
            I => \N__19680\
        );

    \I__4370\ : InMux
    port map (
            O => \N__19697\,
            I => \N__19677\
        );

    \I__4369\ : Span4Mux_v
    port map (
            O => \N__19694\,
            I => \N__19674\
        );

    \I__4368\ : InMux
    port map (
            O => \N__19693\,
            I => \N__19671\
        );

    \I__4367\ : InMux
    port map (
            O => \N__19692\,
            I => \N__19667\
        );

    \I__4366\ : InMux
    port map (
            O => \N__19691\,
            I => \N__19664\
        );

    \I__4365\ : Span4Mux_v
    port map (
            O => \N__19686\,
            I => \N__19658\
        );

    \I__4364\ : LocalMux
    port map (
            O => \N__19683\,
            I => \N__19651\
        );

    \I__4363\ : Span4Mux_v
    port map (
            O => \N__19680\,
            I => \N__19651\
        );

    \I__4362\ : LocalMux
    port map (
            O => \N__19677\,
            I => \N__19651\
        );

    \I__4361\ : Span4Mux_h
    port map (
            O => \N__19674\,
            I => \N__19646\
        );

    \I__4360\ : LocalMux
    port map (
            O => \N__19671\,
            I => \N__19646\
        );

    \I__4359\ : InMux
    port map (
            O => \N__19670\,
            I => \N__19643\
        );

    \I__4358\ : LocalMux
    port map (
            O => \N__19667\,
            I => \N__19638\
        );

    \I__4357\ : LocalMux
    port map (
            O => \N__19664\,
            I => \N__19638\
        );

    \I__4356\ : InMux
    port map (
            O => \N__19663\,
            I => \N__19635\
        );

    \I__4355\ : InMux
    port map (
            O => \N__19662\,
            I => \N__19632\
        );

    \I__4354\ : InMux
    port map (
            O => \N__19661\,
            I => \N__19629\
        );

    \I__4353\ : Span4Mux_h
    port map (
            O => \N__19658\,
            I => \N__19626\
        );

    \I__4352\ : Span4Mux_v
    port map (
            O => \N__19651\,
            I => \N__19623\
        );

    \I__4351\ : Span4Mux_v
    port map (
            O => \N__19646\,
            I => \N__19612\
        );

    \I__4350\ : LocalMux
    port map (
            O => \N__19643\,
            I => \N__19612\
        );

    \I__4349\ : Span4Mux_h
    port map (
            O => \N__19638\,
            I => \N__19612\
        );

    \I__4348\ : LocalMux
    port map (
            O => \N__19635\,
            I => \N__19612\
        );

    \I__4347\ : LocalMux
    port map (
            O => \N__19632\,
            I => \N__19612\
        );

    \I__4346\ : LocalMux
    port map (
            O => \N__19629\,
            I => \transmit_module.Y_DELTA_PATTERN_0\
        );

    \I__4345\ : Odrv4
    port map (
            O => \N__19626\,
            I => \transmit_module.Y_DELTA_PATTERN_0\
        );

    \I__4344\ : Odrv4
    port map (
            O => \N__19623\,
            I => \transmit_module.Y_DELTA_PATTERN_0\
        );

    \I__4343\ : Odrv4
    port map (
            O => \N__19612\,
            I => \transmit_module.Y_DELTA_PATTERN_0\
        );

    \I__4342\ : InMux
    port map (
            O => \N__19603\,
            I => \N__19600\
        );

    \I__4341\ : LocalMux
    port map (
            O => \N__19600\,
            I => \N__19597\
        );

    \I__4340\ : Span4Mux_h
    port map (
            O => \N__19597\,
            I => \N__19594\
        );

    \I__4339\ : Span4Mux_h
    port map (
            O => \N__19594\,
            I => \N__19591\
        );

    \I__4338\ : Odrv4
    port map (
            O => \N__19591\,
            I => \transmit_module.Y_DELTA_PATTERN_99\
        );

    \I__4337\ : InMux
    port map (
            O => \N__19588\,
            I => \N__19584\
        );

    \I__4336\ : InMux
    port map (
            O => \N__19587\,
            I => \N__19579\
        );

    \I__4335\ : LocalMux
    port map (
            O => \N__19584\,
            I => \N__19576\
        );

    \I__4334\ : InMux
    port map (
            O => \N__19583\,
            I => \N__19573\
        );

    \I__4333\ : InMux
    port map (
            O => \N__19582\,
            I => \N__19569\
        );

    \I__4332\ : LocalMux
    port map (
            O => \N__19579\,
            I => \N__19566\
        );

    \I__4331\ : Span4Mux_h
    port map (
            O => \N__19576\,
            I => \N__19563\
        );

    \I__4330\ : LocalMux
    port map (
            O => \N__19573\,
            I => \N__19560\
        );

    \I__4329\ : InMux
    port map (
            O => \N__19572\,
            I => \N__19557\
        );

    \I__4328\ : LocalMux
    port map (
            O => \N__19569\,
            I => \N__19552\
        );

    \I__4327\ : Span4Mux_h
    port map (
            O => \N__19566\,
            I => \N__19552\
        );

    \I__4326\ : Odrv4
    port map (
            O => \N__19563\,
            I => \transmit_module.n4220\
        );

    \I__4325\ : Odrv12
    port map (
            O => \N__19560\,
            I => \transmit_module.n4220\
        );

    \I__4324\ : LocalMux
    port map (
            O => \N__19557\,
            I => \transmit_module.n4220\
        );

    \I__4323\ : Odrv4
    port map (
            O => \N__19552\,
            I => \transmit_module.n4220\
        );

    \I__4322\ : InMux
    port map (
            O => \N__19543\,
            I => \N__19540\
        );

    \I__4321\ : LocalMux
    port map (
            O => \N__19540\,
            I => \N__19537\
        );

    \I__4320\ : Odrv4
    port map (
            O => \N__19537\,
            I => \transmit_module.n192\
        );

    \I__4319\ : InMux
    port map (
            O => \N__19534\,
            I => \N__19529\
        );

    \I__4318\ : CascadeMux
    port map (
            O => \N__19533\,
            I => \N__19526\
        );

    \I__4317\ : InMux
    port map (
            O => \N__19532\,
            I => \N__19522\
        );

    \I__4316\ : LocalMux
    port map (
            O => \N__19529\,
            I => \N__19517\
        );

    \I__4315\ : InMux
    port map (
            O => \N__19526\,
            I => \N__19514\
        );

    \I__4314\ : InMux
    port map (
            O => \N__19525\,
            I => \N__19508\
        );

    \I__4313\ : LocalMux
    port map (
            O => \N__19522\,
            I => \N__19505\
        );

    \I__4312\ : InMux
    port map (
            O => \N__19521\,
            I => \N__19502\
        );

    \I__4311\ : InMux
    port map (
            O => \N__19520\,
            I => \N__19497\
        );

    \I__4310\ : Span4Mux_v
    port map (
            O => \N__19517\,
            I => \N__19487\
        );

    \I__4309\ : LocalMux
    port map (
            O => \N__19514\,
            I => \N__19487\
        );

    \I__4308\ : InMux
    port map (
            O => \N__19513\,
            I => \N__19480\
        );

    \I__4307\ : InMux
    port map (
            O => \N__19512\,
            I => \N__19480\
        );

    \I__4306\ : InMux
    port map (
            O => \N__19511\,
            I => \N__19480\
        );

    \I__4305\ : LocalMux
    port map (
            O => \N__19508\,
            I => \N__19477\
        );

    \I__4304\ : Span4Mux_v
    port map (
            O => \N__19505\,
            I => \N__19472\
        );

    \I__4303\ : LocalMux
    port map (
            O => \N__19502\,
            I => \N__19472\
        );

    \I__4302\ : InMux
    port map (
            O => \N__19501\,
            I => \N__19462\
        );

    \I__4301\ : InMux
    port map (
            O => \N__19500\,
            I => \N__19462\
        );

    \I__4300\ : LocalMux
    port map (
            O => \N__19497\,
            I => \N__19459\
        );

    \I__4299\ : InMux
    port map (
            O => \N__19496\,
            I => \N__19448\
        );

    \I__4298\ : InMux
    port map (
            O => \N__19495\,
            I => \N__19448\
        );

    \I__4297\ : InMux
    port map (
            O => \N__19494\,
            I => \N__19448\
        );

    \I__4296\ : InMux
    port map (
            O => \N__19493\,
            I => \N__19448\
        );

    \I__4295\ : InMux
    port map (
            O => \N__19492\,
            I => \N__19448\
        );

    \I__4294\ : Sp12to4
    port map (
            O => \N__19487\,
            I => \N__19443\
        );

    \I__4293\ : LocalMux
    port map (
            O => \N__19480\,
            I => \N__19443\
        );

    \I__4292\ : Span4Mux_h
    port map (
            O => \N__19477\,
            I => \N__19438\
        );

    \I__4291\ : Span4Mux_h
    port map (
            O => \N__19472\,
            I => \N__19438\
        );

    \I__4290\ : InMux
    port map (
            O => \N__19471\,
            I => \N__19433\
        );

    \I__4289\ : InMux
    port map (
            O => \N__19470\,
            I => \N__19433\
        );

    \I__4288\ : InMux
    port map (
            O => \N__19469\,
            I => \N__19426\
        );

    \I__4287\ : InMux
    port map (
            O => \N__19468\,
            I => \N__19426\
        );

    \I__4286\ : InMux
    port map (
            O => \N__19467\,
            I => \N__19426\
        );

    \I__4285\ : LocalMux
    port map (
            O => \N__19462\,
            I => \transmit_module.n3926\
        );

    \I__4284\ : Odrv12
    port map (
            O => \N__19459\,
            I => \transmit_module.n3926\
        );

    \I__4283\ : LocalMux
    port map (
            O => \N__19448\,
            I => \transmit_module.n3926\
        );

    \I__4282\ : Odrv12
    port map (
            O => \N__19443\,
            I => \transmit_module.n3926\
        );

    \I__4281\ : Odrv4
    port map (
            O => \N__19438\,
            I => \transmit_module.n3926\
        );

    \I__4280\ : LocalMux
    port map (
            O => \N__19433\,
            I => \transmit_module.n3926\
        );

    \I__4279\ : LocalMux
    port map (
            O => \N__19426\,
            I => \transmit_module.n3926\
        );

    \I__4278\ : CEMux
    port map (
            O => \N__19411\,
            I => \N__19407\
        );

    \I__4277\ : CEMux
    port map (
            O => \N__19410\,
            I => \N__19404\
        );

    \I__4276\ : LocalMux
    port map (
            O => \N__19407\,
            I => \N__19401\
        );

    \I__4275\ : LocalMux
    port map (
            O => \N__19404\,
            I => \N__19398\
        );

    \I__4274\ : Span4Mux_h
    port map (
            O => \N__19401\,
            I => \N__19394\
        );

    \I__4273\ : Span4Mux_h
    port map (
            O => \N__19398\,
            I => \N__19391\
        );

    \I__4272\ : InMux
    port map (
            O => \N__19397\,
            I => \N__19388\
        );

    \I__4271\ : Odrv4
    port map (
            O => \N__19394\,
            I => \transmit_module.n2277\
        );

    \I__4270\ : Odrv4
    port map (
            O => \N__19391\,
            I => \transmit_module.n2277\
        );

    \I__4269\ : LocalMux
    port map (
            O => \N__19388\,
            I => \transmit_module.n2277\
        );

    \I__4268\ : InMux
    port map (
            O => \N__19381\,
            I => \N__19378\
        );

    \I__4267\ : LocalMux
    port map (
            O => \N__19378\,
            I => \N__19375\
        );

    \I__4266\ : Odrv4
    port map (
            O => \N__19375\,
            I => \transmit_module.Y_DELTA_PATTERN_42\
        );

    \I__4265\ : InMux
    port map (
            O => \N__19372\,
            I => \N__19369\
        );

    \I__4264\ : LocalMux
    port map (
            O => \N__19369\,
            I => \N__19356\
        );

    \I__4263\ : ClkMux
    port map (
            O => \N__19368\,
            I => \N__19228\
        );

    \I__4262\ : ClkMux
    port map (
            O => \N__19367\,
            I => \N__19228\
        );

    \I__4261\ : ClkMux
    port map (
            O => \N__19366\,
            I => \N__19228\
        );

    \I__4260\ : ClkMux
    port map (
            O => \N__19365\,
            I => \N__19228\
        );

    \I__4259\ : ClkMux
    port map (
            O => \N__19364\,
            I => \N__19228\
        );

    \I__4258\ : ClkMux
    port map (
            O => \N__19363\,
            I => \N__19228\
        );

    \I__4257\ : ClkMux
    port map (
            O => \N__19362\,
            I => \N__19228\
        );

    \I__4256\ : ClkMux
    port map (
            O => \N__19361\,
            I => \N__19228\
        );

    \I__4255\ : ClkMux
    port map (
            O => \N__19360\,
            I => \N__19228\
        );

    \I__4254\ : ClkMux
    port map (
            O => \N__19359\,
            I => \N__19228\
        );

    \I__4253\ : Glb2LocalMux
    port map (
            O => \N__19356\,
            I => \N__19228\
        );

    \I__4252\ : ClkMux
    port map (
            O => \N__19355\,
            I => \N__19228\
        );

    \I__4251\ : ClkMux
    port map (
            O => \N__19354\,
            I => \N__19228\
        );

    \I__4250\ : ClkMux
    port map (
            O => \N__19353\,
            I => \N__19228\
        );

    \I__4249\ : ClkMux
    port map (
            O => \N__19352\,
            I => \N__19228\
        );

    \I__4248\ : ClkMux
    port map (
            O => \N__19351\,
            I => \N__19228\
        );

    \I__4247\ : ClkMux
    port map (
            O => \N__19350\,
            I => \N__19228\
        );

    \I__4246\ : ClkMux
    port map (
            O => \N__19349\,
            I => \N__19228\
        );

    \I__4245\ : ClkMux
    port map (
            O => \N__19348\,
            I => \N__19228\
        );

    \I__4244\ : ClkMux
    port map (
            O => \N__19347\,
            I => \N__19228\
        );

    \I__4243\ : ClkMux
    port map (
            O => \N__19346\,
            I => \N__19228\
        );

    \I__4242\ : ClkMux
    port map (
            O => \N__19345\,
            I => \N__19228\
        );

    \I__4241\ : ClkMux
    port map (
            O => \N__19344\,
            I => \N__19228\
        );

    \I__4240\ : ClkMux
    port map (
            O => \N__19343\,
            I => \N__19228\
        );

    \I__4239\ : ClkMux
    port map (
            O => \N__19342\,
            I => \N__19228\
        );

    \I__4238\ : ClkMux
    port map (
            O => \N__19341\,
            I => \N__19228\
        );

    \I__4237\ : ClkMux
    port map (
            O => \N__19340\,
            I => \N__19228\
        );

    \I__4236\ : ClkMux
    port map (
            O => \N__19339\,
            I => \N__19228\
        );

    \I__4235\ : ClkMux
    port map (
            O => \N__19338\,
            I => \N__19228\
        );

    \I__4234\ : ClkMux
    port map (
            O => \N__19337\,
            I => \N__19228\
        );

    \I__4233\ : ClkMux
    port map (
            O => \N__19336\,
            I => \N__19228\
        );

    \I__4232\ : ClkMux
    port map (
            O => \N__19335\,
            I => \N__19228\
        );

    \I__4231\ : ClkMux
    port map (
            O => \N__19334\,
            I => \N__19228\
        );

    \I__4230\ : ClkMux
    port map (
            O => \N__19333\,
            I => \N__19228\
        );

    \I__4229\ : ClkMux
    port map (
            O => \N__19332\,
            I => \N__19228\
        );

    \I__4228\ : ClkMux
    port map (
            O => \N__19331\,
            I => \N__19228\
        );

    \I__4227\ : ClkMux
    port map (
            O => \N__19330\,
            I => \N__19228\
        );

    \I__4226\ : ClkMux
    port map (
            O => \N__19329\,
            I => \N__19228\
        );

    \I__4225\ : ClkMux
    port map (
            O => \N__19328\,
            I => \N__19228\
        );

    \I__4224\ : ClkMux
    port map (
            O => \N__19327\,
            I => \N__19228\
        );

    \I__4223\ : ClkMux
    port map (
            O => \N__19326\,
            I => \N__19228\
        );

    \I__4222\ : ClkMux
    port map (
            O => \N__19325\,
            I => \N__19228\
        );

    \I__4221\ : ClkMux
    port map (
            O => \N__19324\,
            I => \N__19228\
        );

    \I__4220\ : ClkMux
    port map (
            O => \N__19323\,
            I => \N__19228\
        );

    \I__4219\ : ClkMux
    port map (
            O => \N__19322\,
            I => \N__19228\
        );

    \I__4218\ : ClkMux
    port map (
            O => \N__19321\,
            I => \N__19228\
        );

    \I__4217\ : GlobalMux
    port map (
            O => \N__19228\,
            I => \N__19225\
        );

    \I__4216\ : gio2CtrlBuf
    port map (
            O => \N__19225\,
            I => \DEBUG_c_1_c\
        );

    \I__4215\ : IoInMux
    port map (
            O => \N__19222\,
            I => \N__19219\
        );

    \I__4214\ : LocalMux
    port map (
            O => \N__19219\,
            I => \N__19216\
        );

    \I__4213\ : Span12Mux_s6_h
    port map (
            O => \N__19216\,
            I => \N__19212\
        );

    \I__4212\ : IoInMux
    port map (
            O => \N__19215\,
            I => \N__19209\
        );

    \I__4211\ : Span12Mux_v
    port map (
            O => \N__19212\,
            I => \N__19206\
        );

    \I__4210\ : LocalMux
    port map (
            O => \N__19209\,
            I => \N__19203\
        );

    \I__4209\ : Span12Mux_v
    port map (
            O => \N__19206\,
            I => \N__19200\
        );

    \I__4208\ : IoSpan4Mux
    port map (
            O => \N__19203\,
            I => \N__19197\
        );

    \I__4207\ : Odrv12
    port map (
            O => \N__19200\,
            I => \GB_BUFFER_DEBUG_c_1_c_THRU_CO\
        );

    \I__4206\ : Odrv4
    port map (
            O => \N__19197\,
            I => \GB_BUFFER_DEBUG_c_1_c_THRU_CO\
        );

    \I__4205\ : InMux
    port map (
            O => \N__19192\,
            I => \N__19189\
        );

    \I__4204\ : LocalMux
    port map (
            O => \N__19189\,
            I => \transmit_module.Y_DELTA_PATTERN_29\
        );

    \I__4203\ : InMux
    port map (
            O => \N__19186\,
            I => \N__19183\
        );

    \I__4202\ : LocalMux
    port map (
            O => \N__19183\,
            I => \transmit_module.Y_DELTA_PATTERN_31\
        );

    \I__4201\ : InMux
    port map (
            O => \N__19180\,
            I => \N__19177\
        );

    \I__4200\ : LocalMux
    port map (
            O => \N__19177\,
            I => \transmit_module.Y_DELTA_PATTERN_30\
        );

    \I__4199\ : CascadeMux
    port map (
            O => \N__19174\,
            I => \N__19171\
        );

    \I__4198\ : InMux
    port map (
            O => \N__19171\,
            I => \N__19168\
        );

    \I__4197\ : LocalMux
    port map (
            O => \N__19168\,
            I => \transmit_module.n200\
        );

    \I__4196\ : CascadeMux
    port map (
            O => \N__19165\,
            I => \transmit_module.n215_cascade_\
        );

    \I__4195\ : InMux
    port map (
            O => \N__19162\,
            I => \N__19159\
        );

    \I__4194\ : LocalMux
    port map (
            O => \N__19159\,
            I => \transmit_module.ADDR_Y_COMPONENT_5\
        );

    \I__4193\ : InMux
    port map (
            O => \N__19156\,
            I => \N__19153\
        );

    \I__4192\ : LocalMux
    port map (
            O => \N__19153\,
            I => \transmit_module.n191\
        );

    \I__4191\ : InMux
    port map (
            O => \N__19150\,
            I => \N__19147\
        );

    \I__4190\ : LocalMux
    port map (
            O => \N__19147\,
            I => \N__19144\
        );

    \I__4189\ : Span4Mux_v
    port map (
            O => \N__19144\,
            I => \N__19141\
        );

    \I__4188\ : Odrv4
    port map (
            O => \N__19141\,
            I => \transmit_module.BRAM_ADDR_13_N_258_13\
        );

    \I__4187\ : InMux
    port map (
            O => \N__19138\,
            I => \N__19135\
        );

    \I__4186\ : LocalMux
    port map (
            O => \N__19135\,
            I => \N__19132\
        );

    \I__4185\ : Odrv4
    port map (
            O => \N__19132\,
            I => \transmit_module.n199\
        );

    \I__4184\ : InMux
    port map (
            O => \N__19129\,
            I => \N__19123\
        );

    \I__4183\ : InMux
    port map (
            O => \N__19128\,
            I => \N__19117\
        );

    \I__4182\ : InMux
    port map (
            O => \N__19127\,
            I => \N__19114\
        );

    \I__4181\ : InMux
    port map (
            O => \N__19126\,
            I => \N__19111\
        );

    \I__4180\ : LocalMux
    port map (
            O => \N__19123\,
            I => \N__19108\
        );

    \I__4179\ : InMux
    port map (
            O => \N__19122\,
            I => \N__19105\
        );

    \I__4178\ : CascadeMux
    port map (
            O => \N__19121\,
            I => \N__19096\
        );

    \I__4177\ : InMux
    port map (
            O => \N__19120\,
            I => \N__19092\
        );

    \I__4176\ : LocalMux
    port map (
            O => \N__19117\,
            I => \N__19089\
        );

    \I__4175\ : LocalMux
    port map (
            O => \N__19114\,
            I => \N__19084\
        );

    \I__4174\ : LocalMux
    port map (
            O => \N__19111\,
            I => \N__19084\
        );

    \I__4173\ : Span4Mux_v
    port map (
            O => \N__19108\,
            I => \N__19079\
        );

    \I__4172\ : LocalMux
    port map (
            O => \N__19105\,
            I => \N__19079\
        );

    \I__4171\ : InMux
    port map (
            O => \N__19104\,
            I => \N__19076\
        );

    \I__4170\ : InMux
    port map (
            O => \N__19103\,
            I => \N__19071\
        );

    \I__4169\ : InMux
    port map (
            O => \N__19102\,
            I => \N__19071\
        );

    \I__4168\ : InMux
    port map (
            O => \N__19101\,
            I => \N__19068\
        );

    \I__4167\ : InMux
    port map (
            O => \N__19100\,
            I => \N__19065\
        );

    \I__4166\ : InMux
    port map (
            O => \N__19099\,
            I => \N__19058\
        );

    \I__4165\ : InMux
    port map (
            O => \N__19096\,
            I => \N__19058\
        );

    \I__4164\ : InMux
    port map (
            O => \N__19095\,
            I => \N__19058\
        );

    \I__4163\ : LocalMux
    port map (
            O => \N__19092\,
            I => \N__19053\
        );

    \I__4162\ : Span4Mux_v
    port map (
            O => \N__19089\,
            I => \N__19053\
        );

    \I__4161\ : Span4Mux_h
    port map (
            O => \N__19084\,
            I => \N__19042\
        );

    \I__4160\ : Span4Mux_v
    port map (
            O => \N__19079\,
            I => \N__19042\
        );

    \I__4159\ : LocalMux
    port map (
            O => \N__19076\,
            I => \N__19042\
        );

    \I__4158\ : LocalMux
    port map (
            O => \N__19071\,
            I => \N__19042\
        );

    \I__4157\ : LocalMux
    port map (
            O => \N__19068\,
            I => \N__19042\
        );

    \I__4156\ : LocalMux
    port map (
            O => \N__19065\,
            I => \N__19037\
        );

    \I__4155\ : LocalMux
    port map (
            O => \N__19058\,
            I => \N__19037\
        );

    \I__4154\ : Odrv4
    port map (
            O => \N__19053\,
            I => \transmit_module.n3910\
        );

    \I__4153\ : Odrv4
    port map (
            O => \N__19042\,
            I => \transmit_module.n3910\
        );

    \I__4152\ : Odrv12
    port map (
            O => \N__19037\,
            I => \transmit_module.n3910\
        );

    \I__4151\ : CascadeMux
    port map (
            O => \N__19030\,
            I => \transmit_module.n214_cascade_\
        );

    \I__4150\ : CascadeMux
    port map (
            O => \N__19027\,
            I => \N__19023\
        );

    \I__4149\ : InMux
    port map (
            O => \N__19026\,
            I => \N__19018\
        );

    \I__4148\ : InMux
    port map (
            O => \N__19023\,
            I => \N__19013\
        );

    \I__4147\ : InMux
    port map (
            O => \N__19022\,
            I => \N__19013\
        );

    \I__4146\ : InMux
    port map (
            O => \N__19021\,
            I => \N__19010\
        );

    \I__4145\ : LocalMux
    port map (
            O => \N__19018\,
            I => \transmit_module.TX_ADDR_5\
        );

    \I__4144\ : LocalMux
    port map (
            O => \N__19013\,
            I => \transmit_module.TX_ADDR_5\
        );

    \I__4143\ : LocalMux
    port map (
            O => \N__19010\,
            I => \transmit_module.TX_ADDR_5\
        );

    \I__4142\ : InMux
    port map (
            O => \N__19003\,
            I => \N__19000\
        );

    \I__4141\ : LocalMux
    port map (
            O => \N__19000\,
            I => \N__18997\
        );

    \I__4140\ : Span4Mux_h
    port map (
            O => \N__18997\,
            I => \N__18994\
        );

    \I__4139\ : Odrv4
    port map (
            O => \N__18994\,
            I => \transmit_module.ADDR_Y_COMPONENT_4\
        );

    \I__4138\ : InMux
    port map (
            O => \N__18991\,
            I => \N__18988\
        );

    \I__4137\ : LocalMux
    port map (
            O => \N__18988\,
            I => \N__18984\
        );

    \I__4136\ : CascadeMux
    port map (
            O => \N__18987\,
            I => \N__18979\
        );

    \I__4135\ : Span4Mux_v
    port map (
            O => \N__18984\,
            I => \N__18976\
        );

    \I__4134\ : InMux
    port map (
            O => \N__18983\,
            I => \N__18971\
        );

    \I__4133\ : InMux
    port map (
            O => \N__18982\,
            I => \N__18971\
        );

    \I__4132\ : InMux
    port map (
            O => \N__18979\,
            I => \N__18968\
        );

    \I__4131\ : Odrv4
    port map (
            O => \N__18976\,
            I => \transmit_module.TX_ADDR_4\
        );

    \I__4130\ : LocalMux
    port map (
            O => \N__18971\,
            I => \transmit_module.TX_ADDR_4\
        );

    \I__4129\ : LocalMux
    port map (
            O => \N__18968\,
            I => \transmit_module.TX_ADDR_4\
        );

    \I__4128\ : InMux
    port map (
            O => \N__18961\,
            I => \N__18957\
        );

    \I__4127\ : InMux
    port map (
            O => \N__18960\,
            I => \N__18954\
        );

    \I__4126\ : LocalMux
    port map (
            O => \N__18957\,
            I => \transmit_module.n184\
        );

    \I__4125\ : LocalMux
    port map (
            O => \N__18954\,
            I => \transmit_module.n184\
        );

    \I__4124\ : InMux
    port map (
            O => \N__18949\,
            I => \N__18946\
        );

    \I__4123\ : LocalMux
    port map (
            O => \N__18946\,
            I => \transmit_module.n215\
        );

    \I__4122\ : CascadeMux
    port map (
            O => \N__18943\,
            I => \N__18939\
        );

    \I__4121\ : CascadeMux
    port map (
            O => \N__18942\,
            I => \N__18936\
        );

    \I__4120\ : CascadeBuf
    port map (
            O => \N__18939\,
            I => \N__18933\
        );

    \I__4119\ : CascadeBuf
    port map (
            O => \N__18936\,
            I => \N__18930\
        );

    \I__4118\ : CascadeMux
    port map (
            O => \N__18933\,
            I => \N__18927\
        );

    \I__4117\ : CascadeMux
    port map (
            O => \N__18930\,
            I => \N__18924\
        );

    \I__4116\ : CascadeBuf
    port map (
            O => \N__18927\,
            I => \N__18921\
        );

    \I__4115\ : CascadeBuf
    port map (
            O => \N__18924\,
            I => \N__18918\
        );

    \I__4114\ : CascadeMux
    port map (
            O => \N__18921\,
            I => \N__18915\
        );

    \I__4113\ : CascadeMux
    port map (
            O => \N__18918\,
            I => \N__18912\
        );

    \I__4112\ : CascadeBuf
    port map (
            O => \N__18915\,
            I => \N__18909\
        );

    \I__4111\ : CascadeBuf
    port map (
            O => \N__18912\,
            I => \N__18906\
        );

    \I__4110\ : CascadeMux
    port map (
            O => \N__18909\,
            I => \N__18903\
        );

    \I__4109\ : CascadeMux
    port map (
            O => \N__18906\,
            I => \N__18900\
        );

    \I__4108\ : CascadeBuf
    port map (
            O => \N__18903\,
            I => \N__18897\
        );

    \I__4107\ : CascadeBuf
    port map (
            O => \N__18900\,
            I => \N__18894\
        );

    \I__4106\ : CascadeMux
    port map (
            O => \N__18897\,
            I => \N__18891\
        );

    \I__4105\ : CascadeMux
    port map (
            O => \N__18894\,
            I => \N__18888\
        );

    \I__4104\ : CascadeBuf
    port map (
            O => \N__18891\,
            I => \N__18885\
        );

    \I__4103\ : CascadeBuf
    port map (
            O => \N__18888\,
            I => \N__18882\
        );

    \I__4102\ : CascadeMux
    port map (
            O => \N__18885\,
            I => \N__18879\
        );

    \I__4101\ : CascadeMux
    port map (
            O => \N__18882\,
            I => \N__18876\
        );

    \I__4100\ : CascadeBuf
    port map (
            O => \N__18879\,
            I => \N__18873\
        );

    \I__4099\ : CascadeBuf
    port map (
            O => \N__18876\,
            I => \N__18870\
        );

    \I__4098\ : CascadeMux
    port map (
            O => \N__18873\,
            I => \N__18867\
        );

    \I__4097\ : CascadeMux
    port map (
            O => \N__18870\,
            I => \N__18864\
        );

    \I__4096\ : CascadeBuf
    port map (
            O => \N__18867\,
            I => \N__18861\
        );

    \I__4095\ : CascadeBuf
    port map (
            O => \N__18864\,
            I => \N__18858\
        );

    \I__4094\ : CascadeMux
    port map (
            O => \N__18861\,
            I => \N__18855\
        );

    \I__4093\ : CascadeMux
    port map (
            O => \N__18858\,
            I => \N__18852\
        );

    \I__4092\ : CascadeBuf
    port map (
            O => \N__18855\,
            I => \N__18849\
        );

    \I__4091\ : CascadeBuf
    port map (
            O => \N__18852\,
            I => \N__18846\
        );

    \I__4090\ : CascadeMux
    port map (
            O => \N__18849\,
            I => \N__18843\
        );

    \I__4089\ : CascadeMux
    port map (
            O => \N__18846\,
            I => \N__18840\
        );

    \I__4088\ : CascadeBuf
    port map (
            O => \N__18843\,
            I => \N__18837\
        );

    \I__4087\ : CascadeBuf
    port map (
            O => \N__18840\,
            I => \N__18834\
        );

    \I__4086\ : CascadeMux
    port map (
            O => \N__18837\,
            I => \N__18831\
        );

    \I__4085\ : CascadeMux
    port map (
            O => \N__18834\,
            I => \N__18828\
        );

    \I__4084\ : CascadeBuf
    port map (
            O => \N__18831\,
            I => \N__18825\
        );

    \I__4083\ : CascadeBuf
    port map (
            O => \N__18828\,
            I => \N__18822\
        );

    \I__4082\ : CascadeMux
    port map (
            O => \N__18825\,
            I => \N__18819\
        );

    \I__4081\ : CascadeMux
    port map (
            O => \N__18822\,
            I => \N__18816\
        );

    \I__4080\ : CascadeBuf
    port map (
            O => \N__18819\,
            I => \N__18813\
        );

    \I__4079\ : CascadeBuf
    port map (
            O => \N__18816\,
            I => \N__18810\
        );

    \I__4078\ : CascadeMux
    port map (
            O => \N__18813\,
            I => \N__18807\
        );

    \I__4077\ : CascadeMux
    port map (
            O => \N__18810\,
            I => \N__18804\
        );

    \I__4076\ : CascadeBuf
    port map (
            O => \N__18807\,
            I => \N__18801\
        );

    \I__4075\ : CascadeBuf
    port map (
            O => \N__18804\,
            I => \N__18798\
        );

    \I__4074\ : CascadeMux
    port map (
            O => \N__18801\,
            I => \N__18795\
        );

    \I__4073\ : CascadeMux
    port map (
            O => \N__18798\,
            I => \N__18792\
        );

    \I__4072\ : CascadeBuf
    port map (
            O => \N__18795\,
            I => \N__18789\
        );

    \I__4071\ : CascadeBuf
    port map (
            O => \N__18792\,
            I => \N__18786\
        );

    \I__4070\ : CascadeMux
    port map (
            O => \N__18789\,
            I => \N__18783\
        );

    \I__4069\ : CascadeMux
    port map (
            O => \N__18786\,
            I => \N__18780\
        );

    \I__4068\ : CascadeBuf
    port map (
            O => \N__18783\,
            I => \N__18777\
        );

    \I__4067\ : CascadeBuf
    port map (
            O => \N__18780\,
            I => \N__18774\
        );

    \I__4066\ : CascadeMux
    port map (
            O => \N__18777\,
            I => \N__18771\
        );

    \I__4065\ : CascadeMux
    port map (
            O => \N__18774\,
            I => \N__18768\
        );

    \I__4064\ : CascadeBuf
    port map (
            O => \N__18771\,
            I => \N__18765\
        );

    \I__4063\ : CascadeBuf
    port map (
            O => \N__18768\,
            I => \N__18762\
        );

    \I__4062\ : CascadeMux
    port map (
            O => \N__18765\,
            I => \N__18759\
        );

    \I__4061\ : CascadeMux
    port map (
            O => \N__18762\,
            I => \N__18756\
        );

    \I__4060\ : InMux
    port map (
            O => \N__18759\,
            I => \N__18753\
        );

    \I__4059\ : InMux
    port map (
            O => \N__18756\,
            I => \N__18750\
        );

    \I__4058\ : LocalMux
    port map (
            O => \N__18753\,
            I => \N__18747\
        );

    \I__4057\ : LocalMux
    port map (
            O => \N__18750\,
            I => \N__18744\
        );

    \I__4056\ : Span12Mux_h
    port map (
            O => \N__18747\,
            I => \N__18739\
        );

    \I__4055\ : Span12Mux_h
    port map (
            O => \N__18744\,
            I => \N__18739\
        );

    \I__4054\ : Span12Mux_v
    port map (
            O => \N__18739\,
            I => \N__18736\
        );

    \I__4053\ : Odrv12
    port map (
            O => \N__18736\,
            I => n24
        );

    \I__4052\ : CascadeMux
    port map (
            O => \N__18733\,
            I => \N__18729\
        );

    \I__4051\ : InMux
    port map (
            O => \N__18732\,
            I => \N__18726\
        );

    \I__4050\ : InMux
    port map (
            O => \N__18729\,
            I => \N__18723\
        );

    \I__4049\ : LocalMux
    port map (
            O => \N__18726\,
            I => \transmit_module.n183\
        );

    \I__4048\ : LocalMux
    port map (
            O => \N__18723\,
            I => \transmit_module.n183\
        );

    \I__4047\ : InMux
    port map (
            O => \N__18718\,
            I => \N__18715\
        );

    \I__4046\ : LocalMux
    port map (
            O => \N__18715\,
            I => \transmit_module.n214\
        );

    \I__4045\ : CascadeMux
    port map (
            O => \N__18712\,
            I => \N__18708\
        );

    \I__4044\ : CascadeMux
    port map (
            O => \N__18711\,
            I => \N__18705\
        );

    \I__4043\ : CascadeBuf
    port map (
            O => \N__18708\,
            I => \N__18702\
        );

    \I__4042\ : CascadeBuf
    port map (
            O => \N__18705\,
            I => \N__18699\
        );

    \I__4041\ : CascadeMux
    port map (
            O => \N__18702\,
            I => \N__18696\
        );

    \I__4040\ : CascadeMux
    port map (
            O => \N__18699\,
            I => \N__18693\
        );

    \I__4039\ : CascadeBuf
    port map (
            O => \N__18696\,
            I => \N__18690\
        );

    \I__4038\ : CascadeBuf
    port map (
            O => \N__18693\,
            I => \N__18687\
        );

    \I__4037\ : CascadeMux
    port map (
            O => \N__18690\,
            I => \N__18684\
        );

    \I__4036\ : CascadeMux
    port map (
            O => \N__18687\,
            I => \N__18681\
        );

    \I__4035\ : CascadeBuf
    port map (
            O => \N__18684\,
            I => \N__18678\
        );

    \I__4034\ : CascadeBuf
    port map (
            O => \N__18681\,
            I => \N__18675\
        );

    \I__4033\ : CascadeMux
    port map (
            O => \N__18678\,
            I => \N__18672\
        );

    \I__4032\ : CascadeMux
    port map (
            O => \N__18675\,
            I => \N__18669\
        );

    \I__4031\ : CascadeBuf
    port map (
            O => \N__18672\,
            I => \N__18666\
        );

    \I__4030\ : CascadeBuf
    port map (
            O => \N__18669\,
            I => \N__18663\
        );

    \I__4029\ : CascadeMux
    port map (
            O => \N__18666\,
            I => \N__18660\
        );

    \I__4028\ : CascadeMux
    port map (
            O => \N__18663\,
            I => \N__18657\
        );

    \I__4027\ : CascadeBuf
    port map (
            O => \N__18660\,
            I => \N__18654\
        );

    \I__4026\ : CascadeBuf
    port map (
            O => \N__18657\,
            I => \N__18651\
        );

    \I__4025\ : CascadeMux
    port map (
            O => \N__18654\,
            I => \N__18648\
        );

    \I__4024\ : CascadeMux
    port map (
            O => \N__18651\,
            I => \N__18645\
        );

    \I__4023\ : CascadeBuf
    port map (
            O => \N__18648\,
            I => \N__18642\
        );

    \I__4022\ : CascadeBuf
    port map (
            O => \N__18645\,
            I => \N__18639\
        );

    \I__4021\ : CascadeMux
    port map (
            O => \N__18642\,
            I => \N__18636\
        );

    \I__4020\ : CascadeMux
    port map (
            O => \N__18639\,
            I => \N__18633\
        );

    \I__4019\ : CascadeBuf
    port map (
            O => \N__18636\,
            I => \N__18630\
        );

    \I__4018\ : CascadeBuf
    port map (
            O => \N__18633\,
            I => \N__18627\
        );

    \I__4017\ : CascadeMux
    port map (
            O => \N__18630\,
            I => \N__18624\
        );

    \I__4016\ : CascadeMux
    port map (
            O => \N__18627\,
            I => \N__18621\
        );

    \I__4015\ : CascadeBuf
    port map (
            O => \N__18624\,
            I => \N__18618\
        );

    \I__4014\ : CascadeBuf
    port map (
            O => \N__18621\,
            I => \N__18615\
        );

    \I__4013\ : CascadeMux
    port map (
            O => \N__18618\,
            I => \N__18612\
        );

    \I__4012\ : CascadeMux
    port map (
            O => \N__18615\,
            I => \N__18609\
        );

    \I__4011\ : CascadeBuf
    port map (
            O => \N__18612\,
            I => \N__18606\
        );

    \I__4010\ : CascadeBuf
    port map (
            O => \N__18609\,
            I => \N__18603\
        );

    \I__4009\ : CascadeMux
    port map (
            O => \N__18606\,
            I => \N__18600\
        );

    \I__4008\ : CascadeMux
    port map (
            O => \N__18603\,
            I => \N__18597\
        );

    \I__4007\ : CascadeBuf
    port map (
            O => \N__18600\,
            I => \N__18594\
        );

    \I__4006\ : CascadeBuf
    port map (
            O => \N__18597\,
            I => \N__18591\
        );

    \I__4005\ : CascadeMux
    port map (
            O => \N__18594\,
            I => \N__18588\
        );

    \I__4004\ : CascadeMux
    port map (
            O => \N__18591\,
            I => \N__18585\
        );

    \I__4003\ : CascadeBuf
    port map (
            O => \N__18588\,
            I => \N__18582\
        );

    \I__4002\ : CascadeBuf
    port map (
            O => \N__18585\,
            I => \N__18579\
        );

    \I__4001\ : CascadeMux
    port map (
            O => \N__18582\,
            I => \N__18576\
        );

    \I__4000\ : CascadeMux
    port map (
            O => \N__18579\,
            I => \N__18573\
        );

    \I__3999\ : CascadeBuf
    port map (
            O => \N__18576\,
            I => \N__18570\
        );

    \I__3998\ : CascadeBuf
    port map (
            O => \N__18573\,
            I => \N__18567\
        );

    \I__3997\ : CascadeMux
    port map (
            O => \N__18570\,
            I => \N__18564\
        );

    \I__3996\ : CascadeMux
    port map (
            O => \N__18567\,
            I => \N__18561\
        );

    \I__3995\ : CascadeBuf
    port map (
            O => \N__18564\,
            I => \N__18558\
        );

    \I__3994\ : CascadeBuf
    port map (
            O => \N__18561\,
            I => \N__18555\
        );

    \I__3993\ : CascadeMux
    port map (
            O => \N__18558\,
            I => \N__18552\
        );

    \I__3992\ : CascadeMux
    port map (
            O => \N__18555\,
            I => \N__18549\
        );

    \I__3991\ : CascadeBuf
    port map (
            O => \N__18552\,
            I => \N__18546\
        );

    \I__3990\ : CascadeBuf
    port map (
            O => \N__18549\,
            I => \N__18543\
        );

    \I__3989\ : CascadeMux
    port map (
            O => \N__18546\,
            I => \N__18540\
        );

    \I__3988\ : CascadeMux
    port map (
            O => \N__18543\,
            I => \N__18537\
        );

    \I__3987\ : CascadeBuf
    port map (
            O => \N__18540\,
            I => \N__18534\
        );

    \I__3986\ : CascadeBuf
    port map (
            O => \N__18537\,
            I => \N__18531\
        );

    \I__3985\ : CascadeMux
    port map (
            O => \N__18534\,
            I => \N__18528\
        );

    \I__3984\ : CascadeMux
    port map (
            O => \N__18531\,
            I => \N__18525\
        );

    \I__3983\ : InMux
    port map (
            O => \N__18528\,
            I => \N__18522\
        );

    \I__3982\ : InMux
    port map (
            O => \N__18525\,
            I => \N__18519\
        );

    \I__3981\ : LocalMux
    port map (
            O => \N__18522\,
            I => \N__18516\
        );

    \I__3980\ : LocalMux
    port map (
            O => \N__18519\,
            I => \N__18513\
        );

    \I__3979\ : Span12Mux_h
    port map (
            O => \N__18516\,
            I => \N__18510\
        );

    \I__3978\ : Span12Mux_v
    port map (
            O => \N__18513\,
            I => \N__18507\
        );

    \I__3977\ : Span12Mux_v
    port map (
            O => \N__18510\,
            I => \N__18504\
        );

    \I__3976\ : Odrv12
    port map (
            O => \N__18507\,
            I => n23
        );

    \I__3975\ : Odrv12
    port map (
            O => \N__18504\,
            I => n23
        );

    \I__3974\ : InMux
    port map (
            O => \N__18499\,
            I => \N__18496\
        );

    \I__3973\ : LocalMux
    port map (
            O => \N__18496\,
            I => \transmit_module.Y_DELTA_PATTERN_18\
        );

    \I__3972\ : InMux
    port map (
            O => \N__18493\,
            I => \N__18490\
        );

    \I__3971\ : LocalMux
    port map (
            O => \N__18490\,
            I => \transmit_module.Y_DELTA_PATTERN_21\
        );

    \I__3970\ : InMux
    port map (
            O => \N__18487\,
            I => \N__18484\
        );

    \I__3969\ : LocalMux
    port map (
            O => \N__18484\,
            I => \transmit_module.Y_DELTA_PATTERN_20\
        );

    \I__3968\ : InMux
    port map (
            O => \N__18481\,
            I => \N__18478\
        );

    \I__3967\ : LocalMux
    port map (
            O => \N__18478\,
            I => \transmit_module.Y_DELTA_PATTERN_19\
        );

    \I__3966\ : InMux
    port map (
            O => \N__18475\,
            I => \N__18472\
        );

    \I__3965\ : LocalMux
    port map (
            O => \N__18472\,
            I => \transmit_module.Y_DELTA_PATTERN_1\
        );

    \I__3964\ : InMux
    port map (
            O => \N__18469\,
            I => \N__18466\
        );

    \I__3963\ : LocalMux
    port map (
            O => \N__18466\,
            I => \N__18461\
        );

    \I__3962\ : CascadeMux
    port map (
            O => \N__18465\,
            I => \N__18458\
        );

    \I__3961\ : CascadeMux
    port map (
            O => \N__18464\,
            I => \N__18454\
        );

    \I__3960\ : Span4Mux_h
    port map (
            O => \N__18461\,
            I => \N__18451\
        );

    \I__3959\ : InMux
    port map (
            O => \N__18458\,
            I => \N__18448\
        );

    \I__3958\ : InMux
    port map (
            O => \N__18457\,
            I => \N__18445\
        );

    \I__3957\ : InMux
    port map (
            O => \N__18454\,
            I => \N__18442\
        );

    \I__3956\ : Odrv4
    port map (
            O => \N__18451\,
            I => \transmit_module.TX_ADDR_9\
        );

    \I__3955\ : LocalMux
    port map (
            O => \N__18448\,
            I => \transmit_module.TX_ADDR_9\
        );

    \I__3954\ : LocalMux
    port map (
            O => \N__18445\,
            I => \transmit_module.TX_ADDR_9\
        );

    \I__3953\ : LocalMux
    port map (
            O => \N__18442\,
            I => \transmit_module.TX_ADDR_9\
        );

    \I__3952\ : InMux
    port map (
            O => \N__18433\,
            I => \N__18430\
        );

    \I__3951\ : LocalMux
    port map (
            O => \N__18430\,
            I => \N__18427\
        );

    \I__3950\ : Span4Mux_h
    port map (
            O => \N__18427\,
            I => \N__18424\
        );

    \I__3949\ : Odrv4
    port map (
            O => \N__18424\,
            I => \transmit_module.ADDR_Y_COMPONENT_9\
        );

    \I__3948\ : InMux
    port map (
            O => \N__18421\,
            I => \N__18417\
        );

    \I__3947\ : InMux
    port map (
            O => \N__18420\,
            I => \N__18414\
        );

    \I__3946\ : LocalMux
    port map (
            O => \N__18417\,
            I => \N__18411\
        );

    \I__3945\ : LocalMux
    port map (
            O => \N__18414\,
            I => \N__18408\
        );

    \I__3944\ : Span4Mux_v
    port map (
            O => \N__18411\,
            I => \N__18403\
        );

    \I__3943\ : Span4Mux_h
    port map (
            O => \N__18408\,
            I => \N__18400\
        );

    \I__3942\ : InMux
    port map (
            O => \N__18407\,
            I => \N__18397\
        );

    \I__3941\ : InMux
    port map (
            O => \N__18406\,
            I => \N__18394\
        );

    \I__3940\ : Odrv4
    port map (
            O => \N__18403\,
            I => \transmit_module.TX_ADDR_0\
        );

    \I__3939\ : Odrv4
    port map (
            O => \N__18400\,
            I => \transmit_module.TX_ADDR_0\
        );

    \I__3938\ : LocalMux
    port map (
            O => \N__18397\,
            I => \transmit_module.TX_ADDR_0\
        );

    \I__3937\ : LocalMux
    port map (
            O => \N__18394\,
            I => \transmit_module.TX_ADDR_0\
        );

    \I__3936\ : InMux
    port map (
            O => \N__18385\,
            I => \N__18382\
        );

    \I__3935\ : LocalMux
    port map (
            O => \N__18382\,
            I => \transmit_module.ADDR_Y_COMPONENT_0\
        );

    \I__3934\ : InMux
    port map (
            O => \N__18379\,
            I => \N__18376\
        );

    \I__3933\ : LocalMux
    port map (
            O => \N__18376\,
            I => \N__18370\
        );

    \I__3932\ : InMux
    port map (
            O => \N__18375\,
            I => \N__18367\
        );

    \I__3931\ : InMux
    port map (
            O => \N__18374\,
            I => \N__18364\
        );

    \I__3930\ : InMux
    port map (
            O => \N__18373\,
            I => \N__18361\
        );

    \I__3929\ : Odrv4
    port map (
            O => \N__18370\,
            I => \transmit_module.TX_ADDR_3\
        );

    \I__3928\ : LocalMux
    port map (
            O => \N__18367\,
            I => \transmit_module.TX_ADDR_3\
        );

    \I__3927\ : LocalMux
    port map (
            O => \N__18364\,
            I => \transmit_module.TX_ADDR_3\
        );

    \I__3926\ : LocalMux
    port map (
            O => \N__18361\,
            I => \transmit_module.TX_ADDR_3\
        );

    \I__3925\ : InMux
    port map (
            O => \N__18352\,
            I => \N__18349\
        );

    \I__3924\ : LocalMux
    port map (
            O => \N__18349\,
            I => \transmit_module.ADDR_Y_COMPONENT_3\
        );

    \I__3923\ : InMux
    port map (
            O => \N__18346\,
            I => \N__18343\
        );

    \I__3922\ : LocalMux
    port map (
            O => \N__18343\,
            I => \N__18340\
        );

    \I__3921\ : Odrv4
    port map (
            O => \N__18340\,
            I => \transmit_module.n193\
        );

    \I__3920\ : CascadeMux
    port map (
            O => \N__18337\,
            I => \N__18334\
        );

    \I__3919\ : InMux
    port map (
            O => \N__18334\,
            I => \N__18331\
        );

    \I__3918\ : LocalMux
    port map (
            O => \N__18331\,
            I => \transmit_module.ADDR_Y_COMPONENT_11\
        );

    \I__3917\ : InMux
    port map (
            O => \N__18328\,
            I => \N__18325\
        );

    \I__3916\ : LocalMux
    port map (
            O => \N__18325\,
            I => \transmit_module.ADDR_Y_COMPONENT_1\
        );

    \I__3915\ : InMux
    port map (
            O => \N__18322\,
            I => \N__18316\
        );

    \I__3914\ : InMux
    port map (
            O => \N__18321\,
            I => \N__18313\
        );

    \I__3913\ : InMux
    port map (
            O => \N__18320\,
            I => \N__18310\
        );

    \I__3912\ : InMux
    port map (
            O => \N__18319\,
            I => \N__18307\
        );

    \I__3911\ : LocalMux
    port map (
            O => \N__18316\,
            I => \N__18302\
        );

    \I__3910\ : LocalMux
    port map (
            O => \N__18313\,
            I => \N__18302\
        );

    \I__3909\ : LocalMux
    port map (
            O => \N__18310\,
            I => \N__18299\
        );

    \I__3908\ : LocalMux
    port map (
            O => \N__18307\,
            I => \transmit_module.TX_ADDR_1\
        );

    \I__3907\ : Odrv4
    port map (
            O => \N__18302\,
            I => \transmit_module.TX_ADDR_1\
        );

    \I__3906\ : Odrv4
    port map (
            O => \N__18299\,
            I => \transmit_module.TX_ADDR_1\
        );

    \I__3905\ : InMux
    port map (
            O => \N__18292\,
            I => \N__18288\
        );

    \I__3904\ : InMux
    port map (
            O => \N__18291\,
            I => \N__18285\
        );

    \I__3903\ : LocalMux
    port map (
            O => \N__18288\,
            I => \N__18282\
        );

    \I__3902\ : LocalMux
    port map (
            O => \N__18285\,
            I => \N__18279\
        );

    \I__3901\ : Odrv4
    port map (
            O => \N__18282\,
            I => \transmit_module.n187\
        );

    \I__3900\ : Odrv12
    port map (
            O => \N__18279\,
            I => \transmit_module.n187\
        );

    \I__3899\ : InMux
    port map (
            O => \N__18274\,
            I => \N__18271\
        );

    \I__3898\ : LocalMux
    port map (
            O => \N__18271\,
            I => \N__18268\
        );

    \I__3897\ : Odrv12
    port map (
            O => \N__18268\,
            I => \transmit_module.n218\
        );

    \I__3896\ : CascadeMux
    port map (
            O => \N__18265\,
            I => \N__18262\
        );

    \I__3895\ : CascadeBuf
    port map (
            O => \N__18262\,
            I => \N__18258\
        );

    \I__3894\ : CascadeMux
    port map (
            O => \N__18261\,
            I => \N__18255\
        );

    \I__3893\ : CascadeMux
    port map (
            O => \N__18258\,
            I => \N__18252\
        );

    \I__3892\ : CascadeBuf
    port map (
            O => \N__18255\,
            I => \N__18249\
        );

    \I__3891\ : CascadeBuf
    port map (
            O => \N__18252\,
            I => \N__18246\
        );

    \I__3890\ : CascadeMux
    port map (
            O => \N__18249\,
            I => \N__18243\
        );

    \I__3889\ : CascadeMux
    port map (
            O => \N__18246\,
            I => \N__18240\
        );

    \I__3888\ : CascadeBuf
    port map (
            O => \N__18243\,
            I => \N__18237\
        );

    \I__3887\ : CascadeBuf
    port map (
            O => \N__18240\,
            I => \N__18234\
        );

    \I__3886\ : CascadeMux
    port map (
            O => \N__18237\,
            I => \N__18231\
        );

    \I__3885\ : CascadeMux
    port map (
            O => \N__18234\,
            I => \N__18228\
        );

    \I__3884\ : CascadeBuf
    port map (
            O => \N__18231\,
            I => \N__18225\
        );

    \I__3883\ : CascadeBuf
    port map (
            O => \N__18228\,
            I => \N__18222\
        );

    \I__3882\ : CascadeMux
    port map (
            O => \N__18225\,
            I => \N__18219\
        );

    \I__3881\ : CascadeMux
    port map (
            O => \N__18222\,
            I => \N__18216\
        );

    \I__3880\ : CascadeBuf
    port map (
            O => \N__18219\,
            I => \N__18213\
        );

    \I__3879\ : CascadeBuf
    port map (
            O => \N__18216\,
            I => \N__18210\
        );

    \I__3878\ : CascadeMux
    port map (
            O => \N__18213\,
            I => \N__18207\
        );

    \I__3877\ : CascadeMux
    port map (
            O => \N__18210\,
            I => \N__18204\
        );

    \I__3876\ : CascadeBuf
    port map (
            O => \N__18207\,
            I => \N__18201\
        );

    \I__3875\ : CascadeBuf
    port map (
            O => \N__18204\,
            I => \N__18198\
        );

    \I__3874\ : CascadeMux
    port map (
            O => \N__18201\,
            I => \N__18195\
        );

    \I__3873\ : CascadeMux
    port map (
            O => \N__18198\,
            I => \N__18192\
        );

    \I__3872\ : CascadeBuf
    port map (
            O => \N__18195\,
            I => \N__18189\
        );

    \I__3871\ : CascadeBuf
    port map (
            O => \N__18192\,
            I => \N__18186\
        );

    \I__3870\ : CascadeMux
    port map (
            O => \N__18189\,
            I => \N__18183\
        );

    \I__3869\ : CascadeMux
    port map (
            O => \N__18186\,
            I => \N__18180\
        );

    \I__3868\ : CascadeBuf
    port map (
            O => \N__18183\,
            I => \N__18177\
        );

    \I__3867\ : CascadeBuf
    port map (
            O => \N__18180\,
            I => \N__18174\
        );

    \I__3866\ : CascadeMux
    port map (
            O => \N__18177\,
            I => \N__18171\
        );

    \I__3865\ : CascadeMux
    port map (
            O => \N__18174\,
            I => \N__18168\
        );

    \I__3864\ : CascadeBuf
    port map (
            O => \N__18171\,
            I => \N__18165\
        );

    \I__3863\ : CascadeBuf
    port map (
            O => \N__18168\,
            I => \N__18162\
        );

    \I__3862\ : CascadeMux
    port map (
            O => \N__18165\,
            I => \N__18159\
        );

    \I__3861\ : CascadeMux
    port map (
            O => \N__18162\,
            I => \N__18156\
        );

    \I__3860\ : CascadeBuf
    port map (
            O => \N__18159\,
            I => \N__18153\
        );

    \I__3859\ : CascadeBuf
    port map (
            O => \N__18156\,
            I => \N__18150\
        );

    \I__3858\ : CascadeMux
    port map (
            O => \N__18153\,
            I => \N__18147\
        );

    \I__3857\ : CascadeMux
    port map (
            O => \N__18150\,
            I => \N__18144\
        );

    \I__3856\ : CascadeBuf
    port map (
            O => \N__18147\,
            I => \N__18141\
        );

    \I__3855\ : CascadeBuf
    port map (
            O => \N__18144\,
            I => \N__18138\
        );

    \I__3854\ : CascadeMux
    port map (
            O => \N__18141\,
            I => \N__18135\
        );

    \I__3853\ : CascadeMux
    port map (
            O => \N__18138\,
            I => \N__18132\
        );

    \I__3852\ : CascadeBuf
    port map (
            O => \N__18135\,
            I => \N__18129\
        );

    \I__3851\ : CascadeBuf
    port map (
            O => \N__18132\,
            I => \N__18126\
        );

    \I__3850\ : CascadeMux
    port map (
            O => \N__18129\,
            I => \N__18123\
        );

    \I__3849\ : CascadeMux
    port map (
            O => \N__18126\,
            I => \N__18120\
        );

    \I__3848\ : CascadeBuf
    port map (
            O => \N__18123\,
            I => \N__18117\
        );

    \I__3847\ : CascadeBuf
    port map (
            O => \N__18120\,
            I => \N__18114\
        );

    \I__3846\ : CascadeMux
    port map (
            O => \N__18117\,
            I => \N__18111\
        );

    \I__3845\ : CascadeMux
    port map (
            O => \N__18114\,
            I => \N__18108\
        );

    \I__3844\ : CascadeBuf
    port map (
            O => \N__18111\,
            I => \N__18105\
        );

    \I__3843\ : CascadeBuf
    port map (
            O => \N__18108\,
            I => \N__18102\
        );

    \I__3842\ : CascadeMux
    port map (
            O => \N__18105\,
            I => \N__18099\
        );

    \I__3841\ : CascadeMux
    port map (
            O => \N__18102\,
            I => \N__18096\
        );

    \I__3840\ : CascadeBuf
    port map (
            O => \N__18099\,
            I => \N__18093\
        );

    \I__3839\ : CascadeBuf
    port map (
            O => \N__18096\,
            I => \N__18090\
        );

    \I__3838\ : CascadeMux
    port map (
            O => \N__18093\,
            I => \N__18087\
        );

    \I__3837\ : CascadeMux
    port map (
            O => \N__18090\,
            I => \N__18084\
        );

    \I__3836\ : CascadeBuf
    port map (
            O => \N__18087\,
            I => \N__18081\
        );

    \I__3835\ : InMux
    port map (
            O => \N__18084\,
            I => \N__18078\
        );

    \I__3834\ : CascadeMux
    port map (
            O => \N__18081\,
            I => \N__18075\
        );

    \I__3833\ : LocalMux
    port map (
            O => \N__18078\,
            I => \N__18072\
        );

    \I__3832\ : InMux
    port map (
            O => \N__18075\,
            I => \N__18069\
        );

    \I__3831\ : Span4Mux_v
    port map (
            O => \N__18072\,
            I => \N__18066\
        );

    \I__3830\ : LocalMux
    port map (
            O => \N__18069\,
            I => \N__18063\
        );

    \I__3829\ : Span4Mux_h
    port map (
            O => \N__18066\,
            I => \N__18060\
        );

    \I__3828\ : Span4Mux_v
    port map (
            O => \N__18063\,
            I => \N__18057\
        );

    \I__3827\ : Span4Mux_h
    port map (
            O => \N__18060\,
            I => \N__18052\
        );

    \I__3826\ : Span4Mux_h
    port map (
            O => \N__18057\,
            I => \N__18052\
        );

    \I__3825\ : Odrv4
    port map (
            O => \N__18052\,
            I => n27
        );

    \I__3824\ : InMux
    port map (
            O => \N__18049\,
            I => \N__18046\
        );

    \I__3823\ : LocalMux
    port map (
            O => \N__18046\,
            I => \N__18043\
        );

    \I__3822\ : Span4Mux_h
    port map (
            O => \N__18043\,
            I => \N__18040\
        );

    \I__3821\ : Sp12to4
    port map (
            O => \N__18040\,
            I => \N__18037\
        );

    \I__3820\ : Span12Mux_v
    port map (
            O => \N__18037\,
            I => \N__18034\
        );

    \I__3819\ : Odrv12
    port map (
            O => \N__18034\,
            I => \line_buffer.n678\
        );

    \I__3818\ : CascadeMux
    port map (
            O => \N__18031\,
            I => \N__18028\
        );

    \I__3817\ : InMux
    port map (
            O => \N__18028\,
            I => \N__18025\
        );

    \I__3816\ : LocalMux
    port map (
            O => \N__18025\,
            I => \N__18022\
        );

    \I__3815\ : Odrv12
    port map (
            O => \N__18022\,
            I => \line_buffer.n686\
        );

    \I__3814\ : InMux
    port map (
            O => \N__18019\,
            I => \N__18016\
        );

    \I__3813\ : LocalMux
    port map (
            O => \N__18016\,
            I => \N__18013\
        );

    \I__3812\ : Span4Mux_v
    port map (
            O => \N__18013\,
            I => \N__18010\
        );

    \I__3811\ : Span4Mux_h
    port map (
            O => \N__18010\,
            I => \N__18007\
        );

    \I__3810\ : Span4Mux_h
    port map (
            O => \N__18007\,
            I => \N__18004\
        );

    \I__3809\ : Odrv4
    port map (
            O => \N__18004\,
            I => \line_buffer.n614\
        );

    \I__3808\ : CascadeMux
    port map (
            O => \N__18001\,
            I => \line_buffer.n4188_cascade_\
        );

    \I__3807\ : InMux
    port map (
            O => \N__17998\,
            I => \N__17995\
        );

    \I__3806\ : LocalMux
    port map (
            O => \N__17995\,
            I => \N__17992\
        );

    \I__3805\ : Span4Mux_h
    port map (
            O => \N__17992\,
            I => \N__17989\
        );

    \I__3804\ : Sp12to4
    port map (
            O => \N__17989\,
            I => \N__17986\
        );

    \I__3803\ : Span12Mux_v
    port map (
            O => \N__17986\,
            I => \N__17983\
        );

    \I__3802\ : Odrv12
    port map (
            O => \N__17983\,
            I => \line_buffer.n622\
        );

    \I__3801\ : CascadeMux
    port map (
            O => \N__17980\,
            I => \line_buffer.n4191_cascade_\
        );

    \I__3800\ : InMux
    port map (
            O => \N__17977\,
            I => \N__17974\
        );

    \I__3799\ : LocalMux
    port map (
            O => \N__17974\,
            I => \line_buffer.n4179\
        );

    \I__3798\ : InMux
    port map (
            O => \N__17971\,
            I => \N__17968\
        );

    \I__3797\ : LocalMux
    port map (
            O => \N__17968\,
            I => \N__17965\
        );

    \I__3796\ : Span4Mux_h
    port map (
            O => \N__17965\,
            I => \N__17962\
        );

    \I__3795\ : Span4Mux_v
    port map (
            O => \N__17962\,
            I => \N__17959\
        );

    \I__3794\ : Odrv4
    port map (
            O => \N__17959\,
            I => \TX_DATA_5\
        );

    \I__3793\ : InMux
    port map (
            O => \N__17956\,
            I => \N__17952\
        );

    \I__3792\ : CascadeMux
    port map (
            O => \N__17955\,
            I => \N__17948\
        );

    \I__3791\ : LocalMux
    port map (
            O => \N__17952\,
            I => \N__17945\
        );

    \I__3790\ : InMux
    port map (
            O => \N__17951\,
            I => \N__17941\
        );

    \I__3789\ : InMux
    port map (
            O => \N__17948\,
            I => \N__17938\
        );

    \I__3788\ : Span4Mux_h
    port map (
            O => \N__17945\,
            I => \N__17935\
        );

    \I__3787\ : InMux
    port map (
            O => \N__17944\,
            I => \N__17932\
        );

    \I__3786\ : LocalMux
    port map (
            O => \N__17941\,
            I => \N__17925\
        );

    \I__3785\ : LocalMux
    port map (
            O => \N__17938\,
            I => \N__17925\
        );

    \I__3784\ : Span4Mux_v
    port map (
            O => \N__17935\,
            I => \N__17925\
        );

    \I__3783\ : LocalMux
    port map (
            O => \N__17932\,
            I => \transmit_module.TX_ADDR_10\
        );

    \I__3782\ : Odrv4
    port map (
            O => \N__17925\,
            I => \transmit_module.TX_ADDR_10\
        );

    \I__3781\ : InMux
    port map (
            O => \N__17920\,
            I => \N__17917\
        );

    \I__3780\ : LocalMux
    port map (
            O => \N__17917\,
            I => \N__17914\
        );

    \I__3779\ : Span4Mux_v
    port map (
            O => \N__17914\,
            I => \N__17911\
        );

    \I__3778\ : Span4Mux_v
    port map (
            O => \N__17911\,
            I => \N__17908\
        );

    \I__3777\ : Odrv4
    port map (
            O => \N__17908\,
            I => \transmit_module.n194\
        );

    \I__3776\ : InMux
    port map (
            O => \N__17905\,
            I => \transmit_module.n3665\
        );

    \I__3775\ : InMux
    port map (
            O => \N__17902\,
            I => \transmit_module.n3666\
        );

    \I__3774\ : InMux
    port map (
            O => \N__17899\,
            I => \transmit_module.n3667\
        );

    \I__3773\ : InMux
    port map (
            O => \N__17896\,
            I => \transmit_module.n3668\
        );

    \I__3772\ : CascadeMux
    port map (
            O => \N__17893\,
            I => \N__17890\
        );

    \I__3771\ : InMux
    port map (
            O => \N__17890\,
            I => \N__17887\
        );

    \I__3770\ : LocalMux
    port map (
            O => \N__17887\,
            I => \N__17881\
        );

    \I__3769\ : InMux
    port map (
            O => \N__17886\,
            I => \N__17878\
        );

    \I__3768\ : InMux
    port map (
            O => \N__17885\,
            I => \N__17873\
        );

    \I__3767\ : InMux
    port map (
            O => \N__17884\,
            I => \N__17873\
        );

    \I__3766\ : Odrv4
    port map (
            O => \N__17881\,
            I => \transmit_module.TX_ADDR_8\
        );

    \I__3765\ : LocalMux
    port map (
            O => \N__17878\,
            I => \transmit_module.TX_ADDR_8\
        );

    \I__3764\ : LocalMux
    port map (
            O => \N__17873\,
            I => \transmit_module.TX_ADDR_8\
        );

    \I__3763\ : InMux
    port map (
            O => \N__17866\,
            I => \N__17863\
        );

    \I__3762\ : LocalMux
    port map (
            O => \N__17863\,
            I => \N__17860\
        );

    \I__3761\ : Span4Mux_h
    port map (
            O => \N__17860\,
            I => \N__17857\
        );

    \I__3760\ : Odrv4
    port map (
            O => \N__17857\,
            I => \transmit_module.ADDR_Y_COMPONENT_8\
        );

    \I__3759\ : CascadeMux
    port map (
            O => \N__17854\,
            I => \N__17851\
        );

    \I__3758\ : InMux
    port map (
            O => \N__17851\,
            I => \N__17848\
        );

    \I__3757\ : LocalMux
    port map (
            O => \N__17848\,
            I => \N__17845\
        );

    \I__3756\ : Odrv4
    port map (
            O => \N__17845\,
            I => \transmit_module.n203\
        );

    \I__3755\ : CascadeMux
    port map (
            O => \N__17842\,
            I => \transmit_module.n218_cascade_\
        );

    \I__3754\ : InMux
    port map (
            O => \N__17839\,
            I => \N__17835\
        );

    \I__3753\ : InMux
    port map (
            O => \N__17838\,
            I => \N__17832\
        );

    \I__3752\ : LocalMux
    port map (
            O => \N__17835\,
            I => \N__17829\
        );

    \I__3751\ : LocalMux
    port map (
            O => \N__17832\,
            I => \transmit_module.n188\
        );

    \I__3750\ : Odrv12
    port map (
            O => \N__17829\,
            I => \transmit_module.n188\
        );

    \I__3749\ : InMux
    port map (
            O => \N__17824\,
            I => \N__17818\
        );

    \I__3748\ : InMux
    port map (
            O => \N__17823\,
            I => \N__17815\
        );

    \I__3747\ : InMux
    port map (
            O => \N__17822\,
            I => \N__17812\
        );

    \I__3746\ : InMux
    port map (
            O => \N__17821\,
            I => \N__17809\
        );

    \I__3745\ : LocalMux
    port map (
            O => \N__17818\,
            I => \N__17804\
        );

    \I__3744\ : LocalMux
    port map (
            O => \N__17815\,
            I => \N__17804\
        );

    \I__3743\ : LocalMux
    port map (
            O => \N__17812\,
            I => \transmit_module.TX_ADDR_2\
        );

    \I__3742\ : LocalMux
    port map (
            O => \N__17809\,
            I => \transmit_module.TX_ADDR_2\
        );

    \I__3741\ : Odrv4
    port map (
            O => \N__17804\,
            I => \transmit_module.TX_ADDR_2\
        );

    \I__3740\ : InMux
    port map (
            O => \N__17797\,
            I => \N__17794\
        );

    \I__3739\ : LocalMux
    port map (
            O => \N__17794\,
            I => \N__17791\
        );

    \I__3738\ : Span4Mux_h
    port map (
            O => \N__17791\,
            I => \N__17788\
        );

    \I__3737\ : Odrv4
    port map (
            O => \N__17788\,
            I => \transmit_module.n202\
        );

    \I__3736\ : InMux
    port map (
            O => \N__17785\,
            I => \transmit_module.n3657\
        );

    \I__3735\ : CascadeMux
    port map (
            O => \N__17782\,
            I => \N__17779\
        );

    \I__3734\ : InMux
    port map (
            O => \N__17779\,
            I => \N__17776\
        );

    \I__3733\ : LocalMux
    port map (
            O => \N__17776\,
            I => \N__17773\
        );

    \I__3732\ : Span4Mux_v
    port map (
            O => \N__17773\,
            I => \N__17770\
        );

    \I__3731\ : Odrv4
    port map (
            O => \N__17770\,
            I => \transmit_module.n201\
        );

    \I__3730\ : InMux
    port map (
            O => \N__17767\,
            I => \transmit_module.n3658\
        );

    \I__3729\ : InMux
    port map (
            O => \N__17764\,
            I => \transmit_module.n3659\
        );

    \I__3728\ : InMux
    port map (
            O => \N__17761\,
            I => \transmit_module.n3660\
        );

    \I__3727\ : InMux
    port map (
            O => \N__17758\,
            I => \N__17753\
        );

    \I__3726\ : InMux
    port map (
            O => \N__17757\,
            I => \N__17750\
        );

    \I__3725\ : CascadeMux
    port map (
            O => \N__17756\,
            I => \N__17747\
        );

    \I__3724\ : LocalMux
    port map (
            O => \N__17753\,
            I => \N__17742\
        );

    \I__3723\ : LocalMux
    port map (
            O => \N__17750\,
            I => \N__17742\
        );

    \I__3722\ : InMux
    port map (
            O => \N__17747\,
            I => \N__17738\
        );

    \I__3721\ : Span4Mux_v
    port map (
            O => \N__17742\,
            I => \N__17735\
        );

    \I__3720\ : InMux
    port map (
            O => \N__17741\,
            I => \N__17732\
        );

    \I__3719\ : LocalMux
    port map (
            O => \N__17738\,
            I => \transmit_module.TX_ADDR_6\
        );

    \I__3718\ : Odrv4
    port map (
            O => \N__17735\,
            I => \transmit_module.TX_ADDR_6\
        );

    \I__3717\ : LocalMux
    port map (
            O => \N__17732\,
            I => \transmit_module.TX_ADDR_6\
        );

    \I__3716\ : InMux
    port map (
            O => \N__17725\,
            I => \N__17722\
        );

    \I__3715\ : LocalMux
    port map (
            O => \N__17722\,
            I => \N__17719\
        );

    \I__3714\ : Odrv4
    port map (
            O => \N__17719\,
            I => \transmit_module.n198\
        );

    \I__3713\ : InMux
    port map (
            O => \N__17716\,
            I => \transmit_module.n3661\
        );

    \I__3712\ : InMux
    port map (
            O => \N__17713\,
            I => \N__17709\
        );

    \I__3711\ : CascadeMux
    port map (
            O => \N__17712\,
            I => \N__17705\
        );

    \I__3710\ : LocalMux
    port map (
            O => \N__17709\,
            I => \N__17701\
        );

    \I__3709\ : InMux
    port map (
            O => \N__17708\,
            I => \N__17698\
        );

    \I__3708\ : InMux
    port map (
            O => \N__17705\,
            I => \N__17695\
        );

    \I__3707\ : InMux
    port map (
            O => \N__17704\,
            I => \N__17692\
        );

    \I__3706\ : Odrv4
    port map (
            O => \N__17701\,
            I => \transmit_module.TX_ADDR_7\
        );

    \I__3705\ : LocalMux
    port map (
            O => \N__17698\,
            I => \transmit_module.TX_ADDR_7\
        );

    \I__3704\ : LocalMux
    port map (
            O => \N__17695\,
            I => \transmit_module.TX_ADDR_7\
        );

    \I__3703\ : LocalMux
    port map (
            O => \N__17692\,
            I => \transmit_module.TX_ADDR_7\
        );

    \I__3702\ : InMux
    port map (
            O => \N__17683\,
            I => \N__17680\
        );

    \I__3701\ : LocalMux
    port map (
            O => \N__17680\,
            I => \N__17677\
        );

    \I__3700\ : Span4Mux_h
    port map (
            O => \N__17677\,
            I => \N__17674\
        );

    \I__3699\ : Odrv4
    port map (
            O => \N__17674\,
            I => \transmit_module.n197\
        );

    \I__3698\ : InMux
    port map (
            O => \N__17671\,
            I => \transmit_module.n3662\
        );

    \I__3697\ : InMux
    port map (
            O => \N__17668\,
            I => \N__17665\
        );

    \I__3696\ : LocalMux
    port map (
            O => \N__17665\,
            I => \N__17662\
        );

    \I__3695\ : Span4Mux_h
    port map (
            O => \N__17662\,
            I => \N__17659\
        );

    \I__3694\ : Odrv4
    port map (
            O => \N__17659\,
            I => \transmit_module.n196\
        );

    \I__3693\ : InMux
    port map (
            O => \N__17656\,
            I => \bfn_15_18_0_\
        );

    \I__3692\ : InMux
    port map (
            O => \N__17653\,
            I => \N__17650\
        );

    \I__3691\ : LocalMux
    port map (
            O => \N__17650\,
            I => \N__17647\
        );

    \I__3690\ : Odrv4
    port map (
            O => \N__17647\,
            I => \transmit_module.n195\
        );

    \I__3689\ : InMux
    port map (
            O => \N__17644\,
            I => \transmit_module.n3664\
        );

    \I__3688\ : InMux
    port map (
            O => \N__17641\,
            I => \N__17638\
        );

    \I__3687\ : LocalMux
    port map (
            O => \N__17638\,
            I => \transmit_module.X_DELTA_PATTERN_7\
        );

    \I__3686\ : InMux
    port map (
            O => \N__17635\,
            I => \N__17632\
        );

    \I__3685\ : LocalMux
    port map (
            O => \N__17632\,
            I => \transmit_module.X_DELTA_PATTERN_6\
        );

    \I__3684\ : InMux
    port map (
            O => \N__17629\,
            I => \N__17626\
        );

    \I__3683\ : LocalMux
    port map (
            O => \N__17626\,
            I => \N__17623\
        );

    \I__3682\ : Odrv4
    port map (
            O => \N__17623\,
            I => \transmit_module.X_DELTA_PATTERN_14\
        );

    \I__3681\ : InMux
    port map (
            O => \N__17620\,
            I => \N__17617\
        );

    \I__3680\ : LocalMux
    port map (
            O => \N__17617\,
            I => \transmit_module.X_DELTA_PATTERN_2\
        );

    \I__3679\ : InMux
    port map (
            O => \N__17614\,
            I => \N__17611\
        );

    \I__3678\ : LocalMux
    port map (
            O => \N__17611\,
            I => \transmit_module.X_DELTA_PATTERN_1\
        );

    \I__3677\ : InMux
    port map (
            O => \N__17608\,
            I => \N__17605\
        );

    \I__3676\ : LocalMux
    port map (
            O => \N__17605\,
            I => \transmit_module.X_DELTA_PATTERN_3\
        );

    \I__3675\ : InMux
    port map (
            O => \N__17602\,
            I => \N__17599\
        );

    \I__3674\ : LocalMux
    port map (
            O => \N__17599\,
            I => \transmit_module.X_DELTA_PATTERN_15\
        );

    \I__3673\ : InMux
    port map (
            O => \N__17596\,
            I => \N__17593\
        );

    \I__3672\ : LocalMux
    port map (
            O => \N__17593\,
            I => \transmit_module.X_DELTA_PATTERN_5\
        );

    \I__3671\ : InMux
    port map (
            O => \N__17590\,
            I => \N__17587\
        );

    \I__3670\ : LocalMux
    port map (
            O => \N__17587\,
            I => \transmit_module.X_DELTA_PATTERN_4\
        );

    \I__3669\ : CEMux
    port map (
            O => \N__17584\,
            I => \N__17579\
        );

    \I__3668\ : CEMux
    port map (
            O => \N__17583\,
            I => \N__17575\
        );

    \I__3667\ : CEMux
    port map (
            O => \N__17582\,
            I => \N__17572\
        );

    \I__3666\ : LocalMux
    port map (
            O => \N__17579\,
            I => \N__17568\
        );

    \I__3665\ : CEMux
    port map (
            O => \N__17578\,
            I => \N__17565\
        );

    \I__3664\ : LocalMux
    port map (
            O => \N__17575\,
            I => \N__17562\
        );

    \I__3663\ : LocalMux
    port map (
            O => \N__17572\,
            I => \N__17559\
        );

    \I__3662\ : CEMux
    port map (
            O => \N__17571\,
            I => \N__17556\
        );

    \I__3661\ : Span4Mux_v
    port map (
            O => \N__17568\,
            I => \N__17551\
        );

    \I__3660\ : LocalMux
    port map (
            O => \N__17565\,
            I => \N__17551\
        );

    \I__3659\ : Span4Mux_v
    port map (
            O => \N__17562\,
            I => \N__17548\
        );

    \I__3658\ : Span4Mux_h
    port map (
            O => \N__17559\,
            I => \N__17541\
        );

    \I__3657\ : LocalMux
    port map (
            O => \N__17556\,
            I => \N__17541\
        );

    \I__3656\ : Span4Mux_h
    port map (
            O => \N__17551\,
            I => \N__17541\
        );

    \I__3655\ : Odrv4
    port map (
            O => \N__17548\,
            I => \transmit_module.n2315\
        );

    \I__3654\ : Odrv4
    port map (
            O => \N__17541\,
            I => \transmit_module.n2315\
        );

    \I__3653\ : CascadeMux
    port map (
            O => \N__17536\,
            I => \N__17532\
        );

    \I__3652\ : InMux
    port map (
            O => \N__17535\,
            I => \N__17529\
        );

    \I__3651\ : InMux
    port map (
            O => \N__17532\,
            I => \N__17526\
        );

    \I__3650\ : LocalMux
    port map (
            O => \N__17529\,
            I => \transmit_module.X_DELTA_PATTERN_0\
        );

    \I__3649\ : LocalMux
    port map (
            O => \N__17526\,
            I => \transmit_module.X_DELTA_PATTERN_0\
        );

    \I__3648\ : CascadeMux
    port map (
            O => \N__17521\,
            I => \N__17518\
        );

    \I__3647\ : InMux
    port map (
            O => \N__17518\,
            I => \N__17515\
        );

    \I__3646\ : LocalMux
    port map (
            O => \N__17515\,
            I => \N__17512\
        );

    \I__3645\ : Span4Mux_h
    port map (
            O => \N__17512\,
            I => \N__17509\
        );

    \I__3644\ : Odrv4
    port map (
            O => \N__17509\,
            I => \transmit_module.n204\
        );

    \I__3643\ : InMux
    port map (
            O => \N__17506\,
            I => \transmit_module.n3656\
        );

    \I__3642\ : InMux
    port map (
            O => \N__17503\,
            I => \N__17499\
        );

    \I__3641\ : InMux
    port map (
            O => \N__17502\,
            I => \N__17494\
        );

    \I__3640\ : LocalMux
    port map (
            O => \N__17499\,
            I => \N__17491\
        );

    \I__3639\ : InMux
    port map (
            O => \N__17498\,
            I => \N__17488\
        );

    \I__3638\ : InMux
    port map (
            O => \N__17497\,
            I => \N__17485\
        );

    \I__3637\ : LocalMux
    port map (
            O => \N__17494\,
            I => \receive_module.rx_counter.X_8\
        );

    \I__3636\ : Odrv12
    port map (
            O => \N__17491\,
            I => \receive_module.rx_counter.X_8\
        );

    \I__3635\ : LocalMux
    port map (
            O => \N__17488\,
            I => \receive_module.rx_counter.X_8\
        );

    \I__3634\ : LocalMux
    port map (
            O => \N__17485\,
            I => \receive_module.rx_counter.X_8\
        );

    \I__3633\ : InMux
    port map (
            O => \N__17476\,
            I => \N__17472\
        );

    \I__3632\ : InMux
    port map (
            O => \N__17475\,
            I => \N__17467\
        );

    \I__3631\ : LocalMux
    port map (
            O => \N__17472\,
            I => \N__17464\
        );

    \I__3630\ : InMux
    port map (
            O => \N__17471\,
            I => \N__17461\
        );

    \I__3629\ : InMux
    port map (
            O => \N__17470\,
            I => \N__17458\
        );

    \I__3628\ : LocalMux
    port map (
            O => \N__17467\,
            I => \receive_module.rx_counter.X_9\
        );

    \I__3627\ : Odrv4
    port map (
            O => \N__17464\,
            I => \receive_module.rx_counter.X_9\
        );

    \I__3626\ : LocalMux
    port map (
            O => \N__17461\,
            I => \receive_module.rx_counter.X_9\
        );

    \I__3625\ : LocalMux
    port map (
            O => \N__17458\,
            I => \receive_module.rx_counter.X_9\
        );

    \I__3624\ : InMux
    port map (
            O => \N__17449\,
            I => \N__17446\
        );

    \I__3623\ : LocalMux
    port map (
            O => \N__17446\,
            I => \receive_module.rx_counter.n4219\
        );

    \I__3622\ : CascadeMux
    port map (
            O => \N__17443\,
            I => \N__17438\
        );

    \I__3621\ : InMux
    port map (
            O => \N__17442\,
            I => \N__17434\
        );

    \I__3620\ : InMux
    port map (
            O => \N__17441\,
            I => \N__17431\
        );

    \I__3619\ : InMux
    port map (
            O => \N__17438\,
            I => \N__17426\
        );

    \I__3618\ : InMux
    port map (
            O => \N__17437\,
            I => \N__17426\
        );

    \I__3617\ : LocalMux
    port map (
            O => \N__17434\,
            I => \receive_module.rx_counter.X_7\
        );

    \I__3616\ : LocalMux
    port map (
            O => \N__17431\,
            I => \receive_module.rx_counter.X_7\
        );

    \I__3615\ : LocalMux
    port map (
            O => \N__17426\,
            I => \receive_module.rx_counter.X_7\
        );

    \I__3614\ : CascadeMux
    port map (
            O => \N__17419\,
            I => \receive_module.rx_counter.n4_adj_575_cascade_\
        );

    \I__3613\ : InMux
    port map (
            O => \N__17416\,
            I => \N__17413\
        );

    \I__3612\ : LocalMux
    port map (
            O => \N__17413\,
            I => \N__17409\
        );

    \I__3611\ : InMux
    port map (
            O => \N__17412\,
            I => \N__17404\
        );

    \I__3610\ : Span4Mux_h
    port map (
            O => \N__17409\,
            I => \N__17401\
        );

    \I__3609\ : InMux
    port map (
            O => \N__17408\,
            I => \N__17398\
        );

    \I__3608\ : InMux
    port map (
            O => \N__17407\,
            I => \N__17395\
        );

    \I__3607\ : LocalMux
    port map (
            O => \N__17404\,
            I => \receive_module.rx_counter.X_6\
        );

    \I__3606\ : Odrv4
    port map (
            O => \N__17401\,
            I => \receive_module.rx_counter.X_6\
        );

    \I__3605\ : LocalMux
    port map (
            O => \N__17398\,
            I => \receive_module.rx_counter.X_6\
        );

    \I__3604\ : LocalMux
    port map (
            O => \N__17395\,
            I => \receive_module.rx_counter.X_6\
        );

    \I__3603\ : InMux
    port map (
            O => \N__17386\,
            I => \N__17383\
        );

    \I__3602\ : LocalMux
    port map (
            O => \N__17383\,
            I => \N__17380\
        );

    \I__3601\ : Span4Mux_h
    port map (
            O => \N__17380\,
            I => \N__17377\
        );

    \I__3600\ : Odrv4
    port map (
            O => \N__17377\,
            I => \receive_module.rx_counter.O_VISIBLE_N_86\
        );

    \I__3599\ : InMux
    port map (
            O => \N__17374\,
            I => \N__17371\
        );

    \I__3598\ : LocalMux
    port map (
            O => \N__17371\,
            I => \N__17367\
        );

    \I__3597\ : InMux
    port map (
            O => \N__17370\,
            I => \N__17364\
        );

    \I__3596\ : Odrv4
    port map (
            O => \N__17367\,
            I => \receive_module.rx_counter.n11\
        );

    \I__3595\ : LocalMux
    port map (
            O => \N__17364\,
            I => \receive_module.rx_counter.n11\
        );

    \I__3594\ : IoInMux
    port map (
            O => \N__17359\,
            I => \N__17356\
        );

    \I__3593\ : LocalMux
    port map (
            O => \N__17356\,
            I => \N__17353\
        );

    \I__3592\ : Span4Mux_s1_v
    port map (
            O => \N__17353\,
            I => \N__17350\
        );

    \I__3591\ : Span4Mux_v
    port map (
            O => \N__17350\,
            I => \N__17347\
        );

    \I__3590\ : Span4Mux_v
    port map (
            O => \N__17347\,
            I => \N__17344\
        );

    \I__3589\ : Span4Mux_h
    port map (
            O => \N__17344\,
            I => \N__17340\
        );

    \I__3588\ : InMux
    port map (
            O => \N__17343\,
            I => \N__17337\
        );

    \I__3587\ : Odrv4
    port map (
            O => \N__17340\,
            I => \LED_c\
        );

    \I__3586\ : LocalMux
    port map (
            O => \N__17337\,
            I => \LED_c\
        );

    \I__3585\ : CEMux
    port map (
            O => \N__17332\,
            I => \N__17328\
        );

    \I__3584\ : CEMux
    port map (
            O => \N__17331\,
            I => \N__17325\
        );

    \I__3583\ : LocalMux
    port map (
            O => \N__17328\,
            I => \receive_module.rx_counter.n4222\
        );

    \I__3582\ : LocalMux
    port map (
            O => \N__17325\,
            I => \receive_module.rx_counter.n4222\
        );

    \I__3581\ : InMux
    port map (
            O => \N__17320\,
            I => \N__17317\
        );

    \I__3580\ : LocalMux
    port map (
            O => \N__17317\,
            I => \N__17314\
        );

    \I__3579\ : Span4Mux_v
    port map (
            O => \N__17314\,
            I => \N__17311\
        );

    \I__3578\ : Sp12to4
    port map (
            O => \N__17311\,
            I => \N__17308\
        );

    \I__3577\ : Span12Mux_h
    port map (
            O => \N__17308\,
            I => \N__17305\
        );

    \I__3576\ : Odrv12
    port map (
            O => \N__17305\,
            I => \line_buffer.n623\
        );

    \I__3575\ : InMux
    port map (
            O => \N__17302\,
            I => \N__17299\
        );

    \I__3574\ : LocalMux
    port map (
            O => \N__17299\,
            I => \N__17296\
        );

    \I__3573\ : Span4Mux_v
    port map (
            O => \N__17296\,
            I => \N__17293\
        );

    \I__3572\ : Span4Mux_v
    port map (
            O => \N__17293\,
            I => \N__17290\
        );

    \I__3571\ : Span4Mux_v
    port map (
            O => \N__17290\,
            I => \N__17287\
        );

    \I__3570\ : Sp12to4
    port map (
            O => \N__17287\,
            I => \N__17284\
        );

    \I__3569\ : Odrv12
    port map (
            O => \N__17284\,
            I => \line_buffer.n615\
        );

    \I__3568\ : InMux
    port map (
            O => \N__17281\,
            I => \N__17278\
        );

    \I__3567\ : LocalMux
    port map (
            O => \N__17278\,
            I => \N__17275\
        );

    \I__3566\ : Odrv4
    port map (
            O => \N__17275\,
            I => \line_buffer.n4071\
        );

    \I__3565\ : InMux
    port map (
            O => \N__17272\,
            I => \N__17269\
        );

    \I__3564\ : LocalMux
    port map (
            O => \N__17269\,
            I => \N__17266\
        );

    \I__3563\ : Span12Mux_h
    port map (
            O => \N__17266\,
            I => \N__17263\
        );

    \I__3562\ : Odrv12
    port map (
            O => \N__17263\,
            I => \line_buffer.n646\
        );

    \I__3561\ : CascadeMux
    port map (
            O => \N__17260\,
            I => \N__17257\
        );

    \I__3560\ : InMux
    port map (
            O => \N__17257\,
            I => \N__17254\
        );

    \I__3559\ : LocalMux
    port map (
            O => \N__17254\,
            I => \N__17251\
        );

    \I__3558\ : Span4Mux_v
    port map (
            O => \N__17251\,
            I => \N__17248\
        );

    \I__3557\ : Span4Mux_h
    port map (
            O => \N__17248\,
            I => \N__17245\
        );

    \I__3556\ : Span4Mux_h
    port map (
            O => \N__17245\,
            I => \N__17242\
        );

    \I__3555\ : Odrv4
    port map (
            O => \N__17242\,
            I => \line_buffer.n654\
        );

    \I__3554\ : InMux
    port map (
            O => \N__17239\,
            I => \N__17236\
        );

    \I__3553\ : LocalMux
    port map (
            O => \N__17236\,
            I => \N__17233\
        );

    \I__3552\ : Span4Mux_v
    port map (
            O => \N__17233\,
            I => \N__17230\
        );

    \I__3551\ : Span4Mux_h
    port map (
            O => \N__17230\,
            I => \N__17227\
        );

    \I__3550\ : Sp12to4
    port map (
            O => \N__17227\,
            I => \N__17224\
        );

    \I__3549\ : Span12Mux_v
    port map (
            O => \N__17224\,
            I => \N__17221\
        );

    \I__3548\ : Odrv12
    port map (
            O => \N__17221\,
            I => \line_buffer.n549\
        );

    \I__3547\ : CascadeMux
    port map (
            O => \N__17218\,
            I => \line_buffer.n4176_cascade_\
        );

    \I__3546\ : InMux
    port map (
            O => \N__17215\,
            I => \N__17212\
        );

    \I__3545\ : LocalMux
    port map (
            O => \N__17212\,
            I => \N__17209\
        );

    \I__3544\ : Span4Mux_v
    port map (
            O => \N__17209\,
            I => \N__17206\
        );

    \I__3543\ : Span4Mux_v
    port map (
            O => \N__17206\,
            I => \N__17203\
        );

    \I__3542\ : Sp12to4
    port map (
            O => \N__17203\,
            I => \N__17200\
        );

    \I__3541\ : Odrv12
    port map (
            O => \N__17200\,
            I => \line_buffer.n557\
        );

    \I__3540\ : InMux
    port map (
            O => \N__17197\,
            I => \N__17194\
        );

    \I__3539\ : LocalMux
    port map (
            O => \N__17194\,
            I => \transmit_module.X_DELTA_PATTERN_8\
        );

    \I__3538\ : InMux
    port map (
            O => \N__17191\,
            I => \receive_module.rx_counter.n3706\
        );

    \I__3537\ : InMux
    port map (
            O => \N__17188\,
            I => \N__17184\
        );

    \I__3536\ : InMux
    port map (
            O => \N__17187\,
            I => \N__17181\
        );

    \I__3535\ : LocalMux
    port map (
            O => \N__17184\,
            I => \receive_module.rx_counter.FRAME_COUNTER_2\
        );

    \I__3534\ : LocalMux
    port map (
            O => \N__17181\,
            I => \receive_module.rx_counter.FRAME_COUNTER_2\
        );

    \I__3533\ : InMux
    port map (
            O => \N__17176\,
            I => \receive_module.rx_counter.n3707\
        );

    \I__3532\ : InMux
    port map (
            O => \N__17173\,
            I => \N__17169\
        );

    \I__3531\ : InMux
    port map (
            O => \N__17172\,
            I => \N__17166\
        );

    \I__3530\ : LocalMux
    port map (
            O => \N__17169\,
            I => \receive_module.rx_counter.FRAME_COUNTER_3\
        );

    \I__3529\ : LocalMux
    port map (
            O => \N__17166\,
            I => \receive_module.rx_counter.FRAME_COUNTER_3\
        );

    \I__3528\ : InMux
    port map (
            O => \N__17161\,
            I => \receive_module.rx_counter.n3708\
        );

    \I__3527\ : InMux
    port map (
            O => \N__17158\,
            I => \N__17154\
        );

    \I__3526\ : InMux
    port map (
            O => \N__17157\,
            I => \N__17151\
        );

    \I__3525\ : LocalMux
    port map (
            O => \N__17154\,
            I => \receive_module.rx_counter.FRAME_COUNTER_4\
        );

    \I__3524\ : LocalMux
    port map (
            O => \N__17151\,
            I => \receive_module.rx_counter.FRAME_COUNTER_4\
        );

    \I__3523\ : InMux
    port map (
            O => \N__17146\,
            I => \receive_module.rx_counter.n3709\
        );

    \I__3522\ : InMux
    port map (
            O => \N__17143\,
            I => \receive_module.rx_counter.n3710\
        );

    \I__3521\ : InMux
    port map (
            O => \N__17140\,
            I => \N__17136\
        );

    \I__3520\ : InMux
    port map (
            O => \N__17139\,
            I => \N__17133\
        );

    \I__3519\ : LocalMux
    port map (
            O => \N__17136\,
            I => \receive_module.rx_counter.FRAME_COUNTER_5\
        );

    \I__3518\ : LocalMux
    port map (
            O => \N__17133\,
            I => \receive_module.rx_counter.FRAME_COUNTER_5\
        );

    \I__3517\ : SRMux
    port map (
            O => \N__17128\,
            I => \N__17125\
        );

    \I__3516\ : LocalMux
    port map (
            O => \N__17125\,
            I => \N__17122\
        );

    \I__3515\ : Odrv12
    port map (
            O => \N__17122\,
            I => \receive_module.rx_counter.n2605\
        );

    \I__3514\ : InMux
    port map (
            O => \N__17119\,
            I => \N__17113\
        );

    \I__3513\ : InMux
    port map (
            O => \N__17118\,
            I => \N__17113\
        );

    \I__3512\ : LocalMux
    port map (
            O => \N__17113\,
            I => \receive_module.rx_counter.old_VS\
        );

    \I__3511\ : InMux
    port map (
            O => \N__17110\,
            I => \N__17107\
        );

    \I__3510\ : LocalMux
    port map (
            O => \N__17107\,
            I => \N__17103\
        );

    \I__3509\ : InMux
    port map (
            O => \N__17106\,
            I => \N__17100\
        );

    \I__3508\ : Span4Mux_h
    port map (
            O => \N__17103\,
            I => \N__17094\
        );

    \I__3507\ : LocalMux
    port map (
            O => \N__17100\,
            I => \N__17091\
        );

    \I__3506\ : InMux
    port map (
            O => \N__17099\,
            I => \N__17084\
        );

    \I__3505\ : InMux
    port map (
            O => \N__17098\,
            I => \N__17084\
        );

    \I__3504\ : InMux
    port map (
            O => \N__17097\,
            I => \N__17084\
        );

    \I__3503\ : Sp12to4
    port map (
            O => \N__17094\,
            I => \N__17077\
        );

    \I__3502\ : Span12Mux_h
    port map (
            O => \N__17091\,
            I => \N__17077\
        );

    \I__3501\ : LocalMux
    port map (
            O => \N__17084\,
            I => \N__17077\
        );

    \I__3500\ : Odrv12
    port map (
            O => \N__17077\,
            I => \TVP_VSYNC_c\
        );

    \I__3499\ : CascadeMux
    port map (
            O => \N__17074\,
            I => \N__17068\
        );

    \I__3498\ : InMux
    port map (
            O => \N__17073\,
            I => \N__17065\
        );

    \I__3497\ : InMux
    port map (
            O => \N__17072\,
            I => \N__17062\
        );

    \I__3496\ : InMux
    port map (
            O => \N__17071\,
            I => \N__17057\
        );

    \I__3495\ : InMux
    port map (
            O => \N__17068\,
            I => \N__17057\
        );

    \I__3494\ : LocalMux
    port map (
            O => \N__17065\,
            I => \receive_module.rx_counter.X_5\
        );

    \I__3493\ : LocalMux
    port map (
            O => \N__17062\,
            I => \receive_module.rx_counter.X_5\
        );

    \I__3492\ : LocalMux
    port map (
            O => \N__17057\,
            I => \receive_module.rx_counter.X_5\
        );

    \I__3491\ : InMux
    port map (
            O => \N__17050\,
            I => \N__17044\
        );

    \I__3490\ : InMux
    port map (
            O => \N__17049\,
            I => \N__17041\
        );

    \I__3489\ : InMux
    port map (
            O => \N__17048\,
            I => \N__17036\
        );

    \I__3488\ : InMux
    port map (
            O => \N__17047\,
            I => \N__17036\
        );

    \I__3487\ : LocalMux
    port map (
            O => \N__17044\,
            I => \receive_module.rx_counter.X_4\
        );

    \I__3486\ : LocalMux
    port map (
            O => \N__17041\,
            I => \receive_module.rx_counter.X_4\
        );

    \I__3485\ : LocalMux
    port map (
            O => \N__17036\,
            I => \receive_module.rx_counter.X_4\
        );

    \I__3484\ : InMux
    port map (
            O => \N__17029\,
            I => \N__17023\
        );

    \I__3483\ : InMux
    port map (
            O => \N__17028\,
            I => \N__17020\
        );

    \I__3482\ : InMux
    port map (
            O => \N__17027\,
            I => \N__17015\
        );

    \I__3481\ : InMux
    port map (
            O => \N__17026\,
            I => \N__17015\
        );

    \I__3480\ : LocalMux
    port map (
            O => \N__17023\,
            I => \receive_module.rx_counter.X_3\
        );

    \I__3479\ : LocalMux
    port map (
            O => \N__17020\,
            I => \receive_module.rx_counter.X_3\
        );

    \I__3478\ : LocalMux
    port map (
            O => \N__17015\,
            I => \receive_module.rx_counter.X_3\
        );

    \I__3477\ : CascadeMux
    port map (
            O => \N__17008\,
            I => \N__17005\
        );

    \I__3476\ : InMux
    port map (
            O => \N__17005\,
            I => \N__17001\
        );

    \I__3475\ : CascadeMux
    port map (
            O => \N__17004\,
            I => \N__16998\
        );

    \I__3474\ : LocalMux
    port map (
            O => \N__17001\,
            I => \N__16995\
        );

    \I__3473\ : InMux
    port map (
            O => \N__16998\,
            I => \N__16992\
        );

    \I__3472\ : Odrv4
    port map (
            O => \N__16995\,
            I => \transmit_module.n180\
        );

    \I__3471\ : LocalMux
    port map (
            O => \N__16992\,
            I => \transmit_module.n180\
        );

    \I__3470\ : InMux
    port map (
            O => \N__16987\,
            I => \N__16983\
        );

    \I__3469\ : InMux
    port map (
            O => \N__16986\,
            I => \N__16980\
        );

    \I__3468\ : LocalMux
    port map (
            O => \N__16983\,
            I => \transmit_module.n211\
        );

    \I__3467\ : LocalMux
    port map (
            O => \N__16980\,
            I => \transmit_module.n211\
        );

    \I__3466\ : CascadeMux
    port map (
            O => \N__16975\,
            I => \N__16971\
        );

    \I__3465\ : CascadeMux
    port map (
            O => \N__16974\,
            I => \N__16968\
        );

    \I__3464\ : CascadeBuf
    port map (
            O => \N__16971\,
            I => \N__16965\
        );

    \I__3463\ : CascadeBuf
    port map (
            O => \N__16968\,
            I => \N__16962\
        );

    \I__3462\ : CascadeMux
    port map (
            O => \N__16965\,
            I => \N__16959\
        );

    \I__3461\ : CascadeMux
    port map (
            O => \N__16962\,
            I => \N__16956\
        );

    \I__3460\ : CascadeBuf
    port map (
            O => \N__16959\,
            I => \N__16953\
        );

    \I__3459\ : CascadeBuf
    port map (
            O => \N__16956\,
            I => \N__16950\
        );

    \I__3458\ : CascadeMux
    port map (
            O => \N__16953\,
            I => \N__16947\
        );

    \I__3457\ : CascadeMux
    port map (
            O => \N__16950\,
            I => \N__16944\
        );

    \I__3456\ : CascadeBuf
    port map (
            O => \N__16947\,
            I => \N__16941\
        );

    \I__3455\ : CascadeBuf
    port map (
            O => \N__16944\,
            I => \N__16938\
        );

    \I__3454\ : CascadeMux
    port map (
            O => \N__16941\,
            I => \N__16935\
        );

    \I__3453\ : CascadeMux
    port map (
            O => \N__16938\,
            I => \N__16932\
        );

    \I__3452\ : CascadeBuf
    port map (
            O => \N__16935\,
            I => \N__16929\
        );

    \I__3451\ : CascadeBuf
    port map (
            O => \N__16932\,
            I => \N__16926\
        );

    \I__3450\ : CascadeMux
    port map (
            O => \N__16929\,
            I => \N__16923\
        );

    \I__3449\ : CascadeMux
    port map (
            O => \N__16926\,
            I => \N__16920\
        );

    \I__3448\ : CascadeBuf
    port map (
            O => \N__16923\,
            I => \N__16917\
        );

    \I__3447\ : CascadeBuf
    port map (
            O => \N__16920\,
            I => \N__16914\
        );

    \I__3446\ : CascadeMux
    port map (
            O => \N__16917\,
            I => \N__16911\
        );

    \I__3445\ : CascadeMux
    port map (
            O => \N__16914\,
            I => \N__16908\
        );

    \I__3444\ : CascadeBuf
    port map (
            O => \N__16911\,
            I => \N__16905\
        );

    \I__3443\ : CascadeBuf
    port map (
            O => \N__16908\,
            I => \N__16902\
        );

    \I__3442\ : CascadeMux
    port map (
            O => \N__16905\,
            I => \N__16899\
        );

    \I__3441\ : CascadeMux
    port map (
            O => \N__16902\,
            I => \N__16896\
        );

    \I__3440\ : CascadeBuf
    port map (
            O => \N__16899\,
            I => \N__16893\
        );

    \I__3439\ : CascadeBuf
    port map (
            O => \N__16896\,
            I => \N__16890\
        );

    \I__3438\ : CascadeMux
    port map (
            O => \N__16893\,
            I => \N__16887\
        );

    \I__3437\ : CascadeMux
    port map (
            O => \N__16890\,
            I => \N__16884\
        );

    \I__3436\ : CascadeBuf
    port map (
            O => \N__16887\,
            I => \N__16881\
        );

    \I__3435\ : CascadeBuf
    port map (
            O => \N__16884\,
            I => \N__16878\
        );

    \I__3434\ : CascadeMux
    port map (
            O => \N__16881\,
            I => \N__16875\
        );

    \I__3433\ : CascadeMux
    port map (
            O => \N__16878\,
            I => \N__16872\
        );

    \I__3432\ : CascadeBuf
    port map (
            O => \N__16875\,
            I => \N__16869\
        );

    \I__3431\ : CascadeBuf
    port map (
            O => \N__16872\,
            I => \N__16866\
        );

    \I__3430\ : CascadeMux
    port map (
            O => \N__16869\,
            I => \N__16863\
        );

    \I__3429\ : CascadeMux
    port map (
            O => \N__16866\,
            I => \N__16860\
        );

    \I__3428\ : CascadeBuf
    port map (
            O => \N__16863\,
            I => \N__16857\
        );

    \I__3427\ : CascadeBuf
    port map (
            O => \N__16860\,
            I => \N__16854\
        );

    \I__3426\ : CascadeMux
    port map (
            O => \N__16857\,
            I => \N__16851\
        );

    \I__3425\ : CascadeMux
    port map (
            O => \N__16854\,
            I => \N__16848\
        );

    \I__3424\ : CascadeBuf
    port map (
            O => \N__16851\,
            I => \N__16845\
        );

    \I__3423\ : CascadeBuf
    port map (
            O => \N__16848\,
            I => \N__16842\
        );

    \I__3422\ : CascadeMux
    port map (
            O => \N__16845\,
            I => \N__16839\
        );

    \I__3421\ : CascadeMux
    port map (
            O => \N__16842\,
            I => \N__16836\
        );

    \I__3420\ : CascadeBuf
    port map (
            O => \N__16839\,
            I => \N__16833\
        );

    \I__3419\ : CascadeBuf
    port map (
            O => \N__16836\,
            I => \N__16830\
        );

    \I__3418\ : CascadeMux
    port map (
            O => \N__16833\,
            I => \N__16827\
        );

    \I__3417\ : CascadeMux
    port map (
            O => \N__16830\,
            I => \N__16824\
        );

    \I__3416\ : CascadeBuf
    port map (
            O => \N__16827\,
            I => \N__16821\
        );

    \I__3415\ : CascadeBuf
    port map (
            O => \N__16824\,
            I => \N__16818\
        );

    \I__3414\ : CascadeMux
    port map (
            O => \N__16821\,
            I => \N__16815\
        );

    \I__3413\ : CascadeMux
    port map (
            O => \N__16818\,
            I => \N__16812\
        );

    \I__3412\ : CascadeBuf
    port map (
            O => \N__16815\,
            I => \N__16809\
        );

    \I__3411\ : CascadeBuf
    port map (
            O => \N__16812\,
            I => \N__16806\
        );

    \I__3410\ : CascadeMux
    port map (
            O => \N__16809\,
            I => \N__16803\
        );

    \I__3409\ : CascadeMux
    port map (
            O => \N__16806\,
            I => \N__16800\
        );

    \I__3408\ : CascadeBuf
    port map (
            O => \N__16803\,
            I => \N__16797\
        );

    \I__3407\ : CascadeBuf
    port map (
            O => \N__16800\,
            I => \N__16794\
        );

    \I__3406\ : CascadeMux
    port map (
            O => \N__16797\,
            I => \N__16791\
        );

    \I__3405\ : CascadeMux
    port map (
            O => \N__16794\,
            I => \N__16788\
        );

    \I__3404\ : InMux
    port map (
            O => \N__16791\,
            I => \N__16785\
        );

    \I__3403\ : InMux
    port map (
            O => \N__16788\,
            I => \N__16782\
        );

    \I__3402\ : LocalMux
    port map (
            O => \N__16785\,
            I => \N__16779\
        );

    \I__3401\ : LocalMux
    port map (
            O => \N__16782\,
            I => \N__16776\
        );

    \I__3400\ : Span12Mux_s11_h
    port map (
            O => \N__16779\,
            I => \N__16773\
        );

    \I__3399\ : Span12Mux_s8_h
    port map (
            O => \N__16776\,
            I => \N__16770\
        );

    \I__3398\ : Span12Mux_v
    port map (
            O => \N__16773\,
            I => \N__16765\
        );

    \I__3397\ : Span12Mux_v
    port map (
            O => \N__16770\,
            I => \N__16765\
        );

    \I__3396\ : Odrv12
    port map (
            O => \N__16765\,
            I => n20
        );

    \I__3395\ : InMux
    port map (
            O => \N__16762\,
            I => \N__16757\
        );

    \I__3394\ : InMux
    port map (
            O => \N__16761\,
            I => \N__16752\
        );

    \I__3393\ : InMux
    port map (
            O => \N__16760\,
            I => \N__16749\
        );

    \I__3392\ : LocalMux
    port map (
            O => \N__16757\,
            I => \N__16746\
        );

    \I__3391\ : InMux
    port map (
            O => \N__16756\,
            I => \N__16743\
        );

    \I__3390\ : InMux
    port map (
            O => \N__16755\,
            I => \N__16740\
        );

    \I__3389\ : LocalMux
    port map (
            O => \N__16752\,
            I => \transmit_module.old_VGA_HS\
        );

    \I__3388\ : LocalMux
    port map (
            O => \N__16749\,
            I => \transmit_module.old_VGA_HS\
        );

    \I__3387\ : Odrv4
    port map (
            O => \N__16746\,
            I => \transmit_module.old_VGA_HS\
        );

    \I__3386\ : LocalMux
    port map (
            O => \N__16743\,
            I => \transmit_module.old_VGA_HS\
        );

    \I__3385\ : LocalMux
    port map (
            O => \N__16740\,
            I => \transmit_module.old_VGA_HS\
        );

    \I__3384\ : IoInMux
    port map (
            O => \N__16729\,
            I => \N__16726\
        );

    \I__3383\ : LocalMux
    port map (
            O => \N__16726\,
            I => \N__16723\
        );

    \I__3382\ : Span4Mux_s0_h
    port map (
            O => \N__16723\,
            I => \N__16720\
        );

    \I__3381\ : Span4Mux_h
    port map (
            O => \N__16720\,
            I => \N__16714\
        );

    \I__3380\ : InMux
    port map (
            O => \N__16719\,
            I => \N__16709\
        );

    \I__3379\ : InMux
    port map (
            O => \N__16718\,
            I => \N__16706\
        );

    \I__3378\ : InMux
    port map (
            O => \N__16717\,
            I => \N__16702\
        );

    \I__3377\ : Span4Mux_h
    port map (
            O => \N__16714\,
            I => \N__16699\
        );

    \I__3376\ : InMux
    port map (
            O => \N__16713\,
            I => \N__16694\
        );

    \I__3375\ : InMux
    port map (
            O => \N__16712\,
            I => \N__16694\
        );

    \I__3374\ : LocalMux
    port map (
            O => \N__16709\,
            I => \N__16689\
        );

    \I__3373\ : LocalMux
    port map (
            O => \N__16706\,
            I => \N__16689\
        );

    \I__3372\ : InMux
    port map (
            O => \N__16705\,
            I => \N__16686\
        );

    \I__3371\ : LocalMux
    port map (
            O => \N__16702\,
            I => \N__16683\
        );

    \I__3370\ : Span4Mux_h
    port map (
            O => \N__16699\,
            I => \N__16678\
        );

    \I__3369\ : LocalMux
    port map (
            O => \N__16694\,
            I => \N__16678\
        );

    \I__3368\ : Span12Mux_v
    port map (
            O => \N__16689\,
            I => \N__16675\
        );

    \I__3367\ : LocalMux
    port map (
            O => \N__16686\,
            I => \N__16668\
        );

    \I__3366\ : Span4Mux_v
    port map (
            O => \N__16683\,
            I => \N__16668\
        );

    \I__3365\ : Span4Mux_v
    port map (
            O => \N__16678\,
            I => \N__16668\
        );

    \I__3364\ : Odrv12
    port map (
            O => \N__16675\,
            I => \ADV_HSYNC_c\
        );

    \I__3363\ : Odrv4
    port map (
            O => \N__16668\,
            I => \ADV_HSYNC_c\
        );

    \I__3362\ : CascadeMux
    port map (
            O => \N__16663\,
            I => \N__16660\
        );

    \I__3361\ : InMux
    port map (
            O => \N__16660\,
            I => \N__16657\
        );

    \I__3360\ : LocalMux
    port map (
            O => \N__16657\,
            I => \transmit_module.n181\
        );

    \I__3359\ : InMux
    port map (
            O => \N__16654\,
            I => \N__16650\
        );

    \I__3358\ : InMux
    port map (
            O => \N__16653\,
            I => \N__16647\
        );

    \I__3357\ : LocalMux
    port map (
            O => \N__16650\,
            I => \transmit_module.n212\
        );

    \I__3356\ : LocalMux
    port map (
            O => \N__16647\,
            I => \transmit_module.n212\
        );

    \I__3355\ : CascadeMux
    port map (
            O => \N__16642\,
            I => \transmit_module.n181_cascade_\
        );

    \I__3354\ : CascadeMux
    port map (
            O => \N__16639\,
            I => \N__16635\
        );

    \I__3353\ : CascadeMux
    port map (
            O => \N__16638\,
            I => \N__16632\
        );

    \I__3352\ : CascadeBuf
    port map (
            O => \N__16635\,
            I => \N__16629\
        );

    \I__3351\ : CascadeBuf
    port map (
            O => \N__16632\,
            I => \N__16626\
        );

    \I__3350\ : CascadeMux
    port map (
            O => \N__16629\,
            I => \N__16623\
        );

    \I__3349\ : CascadeMux
    port map (
            O => \N__16626\,
            I => \N__16620\
        );

    \I__3348\ : CascadeBuf
    port map (
            O => \N__16623\,
            I => \N__16617\
        );

    \I__3347\ : CascadeBuf
    port map (
            O => \N__16620\,
            I => \N__16614\
        );

    \I__3346\ : CascadeMux
    port map (
            O => \N__16617\,
            I => \N__16611\
        );

    \I__3345\ : CascadeMux
    port map (
            O => \N__16614\,
            I => \N__16608\
        );

    \I__3344\ : CascadeBuf
    port map (
            O => \N__16611\,
            I => \N__16605\
        );

    \I__3343\ : CascadeBuf
    port map (
            O => \N__16608\,
            I => \N__16602\
        );

    \I__3342\ : CascadeMux
    port map (
            O => \N__16605\,
            I => \N__16599\
        );

    \I__3341\ : CascadeMux
    port map (
            O => \N__16602\,
            I => \N__16596\
        );

    \I__3340\ : CascadeBuf
    port map (
            O => \N__16599\,
            I => \N__16593\
        );

    \I__3339\ : CascadeBuf
    port map (
            O => \N__16596\,
            I => \N__16590\
        );

    \I__3338\ : CascadeMux
    port map (
            O => \N__16593\,
            I => \N__16587\
        );

    \I__3337\ : CascadeMux
    port map (
            O => \N__16590\,
            I => \N__16584\
        );

    \I__3336\ : CascadeBuf
    port map (
            O => \N__16587\,
            I => \N__16581\
        );

    \I__3335\ : CascadeBuf
    port map (
            O => \N__16584\,
            I => \N__16578\
        );

    \I__3334\ : CascadeMux
    port map (
            O => \N__16581\,
            I => \N__16575\
        );

    \I__3333\ : CascadeMux
    port map (
            O => \N__16578\,
            I => \N__16572\
        );

    \I__3332\ : CascadeBuf
    port map (
            O => \N__16575\,
            I => \N__16569\
        );

    \I__3331\ : CascadeBuf
    port map (
            O => \N__16572\,
            I => \N__16566\
        );

    \I__3330\ : CascadeMux
    port map (
            O => \N__16569\,
            I => \N__16563\
        );

    \I__3329\ : CascadeMux
    port map (
            O => \N__16566\,
            I => \N__16560\
        );

    \I__3328\ : CascadeBuf
    port map (
            O => \N__16563\,
            I => \N__16557\
        );

    \I__3327\ : CascadeBuf
    port map (
            O => \N__16560\,
            I => \N__16554\
        );

    \I__3326\ : CascadeMux
    port map (
            O => \N__16557\,
            I => \N__16551\
        );

    \I__3325\ : CascadeMux
    port map (
            O => \N__16554\,
            I => \N__16548\
        );

    \I__3324\ : CascadeBuf
    port map (
            O => \N__16551\,
            I => \N__16545\
        );

    \I__3323\ : CascadeBuf
    port map (
            O => \N__16548\,
            I => \N__16542\
        );

    \I__3322\ : CascadeMux
    port map (
            O => \N__16545\,
            I => \N__16539\
        );

    \I__3321\ : CascadeMux
    port map (
            O => \N__16542\,
            I => \N__16536\
        );

    \I__3320\ : CascadeBuf
    port map (
            O => \N__16539\,
            I => \N__16533\
        );

    \I__3319\ : CascadeBuf
    port map (
            O => \N__16536\,
            I => \N__16530\
        );

    \I__3318\ : CascadeMux
    port map (
            O => \N__16533\,
            I => \N__16527\
        );

    \I__3317\ : CascadeMux
    port map (
            O => \N__16530\,
            I => \N__16524\
        );

    \I__3316\ : CascadeBuf
    port map (
            O => \N__16527\,
            I => \N__16521\
        );

    \I__3315\ : CascadeBuf
    port map (
            O => \N__16524\,
            I => \N__16518\
        );

    \I__3314\ : CascadeMux
    port map (
            O => \N__16521\,
            I => \N__16515\
        );

    \I__3313\ : CascadeMux
    port map (
            O => \N__16518\,
            I => \N__16512\
        );

    \I__3312\ : CascadeBuf
    port map (
            O => \N__16515\,
            I => \N__16509\
        );

    \I__3311\ : CascadeBuf
    port map (
            O => \N__16512\,
            I => \N__16506\
        );

    \I__3310\ : CascadeMux
    port map (
            O => \N__16509\,
            I => \N__16503\
        );

    \I__3309\ : CascadeMux
    port map (
            O => \N__16506\,
            I => \N__16500\
        );

    \I__3308\ : CascadeBuf
    port map (
            O => \N__16503\,
            I => \N__16497\
        );

    \I__3307\ : CascadeBuf
    port map (
            O => \N__16500\,
            I => \N__16494\
        );

    \I__3306\ : CascadeMux
    port map (
            O => \N__16497\,
            I => \N__16491\
        );

    \I__3305\ : CascadeMux
    port map (
            O => \N__16494\,
            I => \N__16488\
        );

    \I__3304\ : CascadeBuf
    port map (
            O => \N__16491\,
            I => \N__16485\
        );

    \I__3303\ : CascadeBuf
    port map (
            O => \N__16488\,
            I => \N__16482\
        );

    \I__3302\ : CascadeMux
    port map (
            O => \N__16485\,
            I => \N__16479\
        );

    \I__3301\ : CascadeMux
    port map (
            O => \N__16482\,
            I => \N__16476\
        );

    \I__3300\ : CascadeBuf
    port map (
            O => \N__16479\,
            I => \N__16473\
        );

    \I__3299\ : CascadeBuf
    port map (
            O => \N__16476\,
            I => \N__16470\
        );

    \I__3298\ : CascadeMux
    port map (
            O => \N__16473\,
            I => \N__16467\
        );

    \I__3297\ : CascadeMux
    port map (
            O => \N__16470\,
            I => \N__16464\
        );

    \I__3296\ : CascadeBuf
    port map (
            O => \N__16467\,
            I => \N__16461\
        );

    \I__3295\ : CascadeBuf
    port map (
            O => \N__16464\,
            I => \N__16458\
        );

    \I__3294\ : CascadeMux
    port map (
            O => \N__16461\,
            I => \N__16455\
        );

    \I__3293\ : CascadeMux
    port map (
            O => \N__16458\,
            I => \N__16452\
        );

    \I__3292\ : InMux
    port map (
            O => \N__16455\,
            I => \N__16449\
        );

    \I__3291\ : InMux
    port map (
            O => \N__16452\,
            I => \N__16446\
        );

    \I__3290\ : LocalMux
    port map (
            O => \N__16449\,
            I => \N__16443\
        );

    \I__3289\ : LocalMux
    port map (
            O => \N__16446\,
            I => \N__16440\
        );

    \I__3288\ : Span12Mux_h
    port map (
            O => \N__16443\,
            I => \N__16435\
        );

    \I__3287\ : Span12Mux_h
    port map (
            O => \N__16440\,
            I => \N__16435\
        );

    \I__3286\ : Span12Mux_v
    port map (
            O => \N__16435\,
            I => \N__16432\
        );

    \I__3285\ : Odrv12
    port map (
            O => \N__16432\,
            I => n21
        );

    \I__3284\ : InMux
    port map (
            O => \N__16429\,
            I => \N__16426\
        );

    \I__3283\ : LocalMux
    port map (
            O => \N__16426\,
            I => \N__16423\
        );

    \I__3282\ : Odrv4
    port map (
            O => \N__16423\,
            I => \transmit_module.ADDR_Y_COMPONENT_7\
        );

    \I__3281\ : InMux
    port map (
            O => \N__16420\,
            I => \N__16417\
        );

    \I__3280\ : LocalMux
    port map (
            O => \N__16417\,
            I => \transmit_module.ADDR_Y_COMPONENT_6\
        );

    \I__3279\ : InMux
    port map (
            O => \N__16414\,
            I => \N__16410\
        );

    \I__3278\ : InMux
    port map (
            O => \N__16413\,
            I => \N__16407\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__16410\,
            I => \N__16404\
        );

    \I__3276\ : LocalMux
    port map (
            O => \N__16407\,
            I => \N__16401\
        );

    \I__3275\ : Span4Mux_v
    port map (
            O => \N__16404\,
            I => \N__16398\
        );

    \I__3274\ : Odrv12
    port map (
            O => \N__16401\,
            I => \transmit_module.n182\
        );

    \I__3273\ : Odrv4
    port map (
            O => \N__16398\,
            I => \transmit_module.n182\
        );

    \I__3272\ : InMux
    port map (
            O => \N__16393\,
            I => \N__16389\
        );

    \I__3271\ : InMux
    port map (
            O => \N__16392\,
            I => \N__16386\
        );

    \I__3270\ : LocalMux
    port map (
            O => \N__16389\,
            I => \receive_module.rx_counter.FRAME_COUNTER_0\
        );

    \I__3269\ : LocalMux
    port map (
            O => \N__16386\,
            I => \receive_module.rx_counter.FRAME_COUNTER_0\
        );

    \I__3268\ : InMux
    port map (
            O => \N__16381\,
            I => \bfn_15_8_0_\
        );

    \I__3267\ : InMux
    port map (
            O => \N__16378\,
            I => \N__16374\
        );

    \I__3266\ : InMux
    port map (
            O => \N__16377\,
            I => \N__16371\
        );

    \I__3265\ : LocalMux
    port map (
            O => \N__16374\,
            I => \receive_module.rx_counter.FRAME_COUNTER_1\
        );

    \I__3264\ : LocalMux
    port map (
            O => \N__16371\,
            I => \receive_module.rx_counter.FRAME_COUNTER_1\
        );

    \I__3263\ : InMux
    port map (
            O => \N__16366\,
            I => \N__16363\
        );

    \I__3262\ : LocalMux
    port map (
            O => \N__16363\,
            I => \transmit_module.ADDR_Y_COMPONENT_2\
        );

    \I__3261\ : InMux
    port map (
            O => \N__16360\,
            I => \N__16357\
        );

    \I__3260\ : LocalMux
    port map (
            O => \N__16357\,
            I => \N__16354\
        );

    \I__3259\ : Span4Mux_h
    port map (
            O => \N__16354\,
            I => \N__16351\
        );

    \I__3258\ : Odrv4
    port map (
            O => \N__16351\,
            I => \transmit_module.n219\
        );

    \I__3257\ : CascadeMux
    port map (
            O => \N__16348\,
            I => \transmit_module.n179_cascade_\
        );

    \I__3256\ : InMux
    port map (
            O => \N__16345\,
            I => \N__16342\
        );

    \I__3255\ : LocalMux
    port map (
            O => \N__16342\,
            I => \N__16338\
        );

    \I__3254\ : InMux
    port map (
            O => \N__16341\,
            I => \N__16335\
        );

    \I__3253\ : Span12Mux_s6_v
    port map (
            O => \N__16338\,
            I => \N__16332\
        );

    \I__3252\ : LocalMux
    port map (
            O => \N__16335\,
            I => \transmit_module.n213\
        );

    \I__3251\ : Odrv12
    port map (
            O => \N__16332\,
            I => \transmit_module.n213\
        );

    \I__3250\ : InMux
    port map (
            O => \N__16327\,
            I => \N__16324\
        );

    \I__3249\ : LocalMux
    port map (
            O => \N__16324\,
            I => \transmit_module.n179\
        );

    \I__3248\ : InMux
    port map (
            O => \N__16321\,
            I => \N__16317\
        );

    \I__3247\ : InMux
    port map (
            O => \N__16320\,
            I => \N__16314\
        );

    \I__3246\ : LocalMux
    port map (
            O => \N__16317\,
            I => \transmit_module.n210\
        );

    \I__3245\ : LocalMux
    port map (
            O => \N__16314\,
            I => \transmit_module.n210\
        );

    \I__3244\ : CascadeMux
    port map (
            O => \N__16309\,
            I => \N__16305\
        );

    \I__3243\ : CascadeMux
    port map (
            O => \N__16308\,
            I => \N__16302\
        );

    \I__3242\ : CascadeBuf
    port map (
            O => \N__16305\,
            I => \N__16299\
        );

    \I__3241\ : CascadeBuf
    port map (
            O => \N__16302\,
            I => \N__16296\
        );

    \I__3240\ : CascadeMux
    port map (
            O => \N__16299\,
            I => \N__16293\
        );

    \I__3239\ : CascadeMux
    port map (
            O => \N__16296\,
            I => \N__16290\
        );

    \I__3238\ : CascadeBuf
    port map (
            O => \N__16293\,
            I => \N__16287\
        );

    \I__3237\ : CascadeBuf
    port map (
            O => \N__16290\,
            I => \N__16284\
        );

    \I__3236\ : CascadeMux
    port map (
            O => \N__16287\,
            I => \N__16281\
        );

    \I__3235\ : CascadeMux
    port map (
            O => \N__16284\,
            I => \N__16278\
        );

    \I__3234\ : CascadeBuf
    port map (
            O => \N__16281\,
            I => \N__16275\
        );

    \I__3233\ : CascadeBuf
    port map (
            O => \N__16278\,
            I => \N__16272\
        );

    \I__3232\ : CascadeMux
    port map (
            O => \N__16275\,
            I => \N__16269\
        );

    \I__3231\ : CascadeMux
    port map (
            O => \N__16272\,
            I => \N__16266\
        );

    \I__3230\ : CascadeBuf
    port map (
            O => \N__16269\,
            I => \N__16263\
        );

    \I__3229\ : CascadeBuf
    port map (
            O => \N__16266\,
            I => \N__16260\
        );

    \I__3228\ : CascadeMux
    port map (
            O => \N__16263\,
            I => \N__16257\
        );

    \I__3227\ : CascadeMux
    port map (
            O => \N__16260\,
            I => \N__16254\
        );

    \I__3226\ : CascadeBuf
    port map (
            O => \N__16257\,
            I => \N__16251\
        );

    \I__3225\ : CascadeBuf
    port map (
            O => \N__16254\,
            I => \N__16248\
        );

    \I__3224\ : CascadeMux
    port map (
            O => \N__16251\,
            I => \N__16245\
        );

    \I__3223\ : CascadeMux
    port map (
            O => \N__16248\,
            I => \N__16242\
        );

    \I__3222\ : CascadeBuf
    port map (
            O => \N__16245\,
            I => \N__16239\
        );

    \I__3221\ : CascadeBuf
    port map (
            O => \N__16242\,
            I => \N__16236\
        );

    \I__3220\ : CascadeMux
    port map (
            O => \N__16239\,
            I => \N__16233\
        );

    \I__3219\ : CascadeMux
    port map (
            O => \N__16236\,
            I => \N__16230\
        );

    \I__3218\ : CascadeBuf
    port map (
            O => \N__16233\,
            I => \N__16227\
        );

    \I__3217\ : CascadeBuf
    port map (
            O => \N__16230\,
            I => \N__16224\
        );

    \I__3216\ : CascadeMux
    port map (
            O => \N__16227\,
            I => \N__16221\
        );

    \I__3215\ : CascadeMux
    port map (
            O => \N__16224\,
            I => \N__16218\
        );

    \I__3214\ : CascadeBuf
    port map (
            O => \N__16221\,
            I => \N__16215\
        );

    \I__3213\ : CascadeBuf
    port map (
            O => \N__16218\,
            I => \N__16212\
        );

    \I__3212\ : CascadeMux
    port map (
            O => \N__16215\,
            I => \N__16209\
        );

    \I__3211\ : CascadeMux
    port map (
            O => \N__16212\,
            I => \N__16206\
        );

    \I__3210\ : CascadeBuf
    port map (
            O => \N__16209\,
            I => \N__16203\
        );

    \I__3209\ : CascadeBuf
    port map (
            O => \N__16206\,
            I => \N__16200\
        );

    \I__3208\ : CascadeMux
    port map (
            O => \N__16203\,
            I => \N__16197\
        );

    \I__3207\ : CascadeMux
    port map (
            O => \N__16200\,
            I => \N__16194\
        );

    \I__3206\ : CascadeBuf
    port map (
            O => \N__16197\,
            I => \N__16191\
        );

    \I__3205\ : CascadeBuf
    port map (
            O => \N__16194\,
            I => \N__16188\
        );

    \I__3204\ : CascadeMux
    port map (
            O => \N__16191\,
            I => \N__16185\
        );

    \I__3203\ : CascadeMux
    port map (
            O => \N__16188\,
            I => \N__16182\
        );

    \I__3202\ : CascadeBuf
    port map (
            O => \N__16185\,
            I => \N__16179\
        );

    \I__3201\ : CascadeBuf
    port map (
            O => \N__16182\,
            I => \N__16176\
        );

    \I__3200\ : CascadeMux
    port map (
            O => \N__16179\,
            I => \N__16173\
        );

    \I__3199\ : CascadeMux
    port map (
            O => \N__16176\,
            I => \N__16170\
        );

    \I__3198\ : CascadeBuf
    port map (
            O => \N__16173\,
            I => \N__16167\
        );

    \I__3197\ : CascadeBuf
    port map (
            O => \N__16170\,
            I => \N__16164\
        );

    \I__3196\ : CascadeMux
    port map (
            O => \N__16167\,
            I => \N__16161\
        );

    \I__3195\ : CascadeMux
    port map (
            O => \N__16164\,
            I => \N__16158\
        );

    \I__3194\ : CascadeBuf
    port map (
            O => \N__16161\,
            I => \N__16155\
        );

    \I__3193\ : CascadeBuf
    port map (
            O => \N__16158\,
            I => \N__16152\
        );

    \I__3192\ : CascadeMux
    port map (
            O => \N__16155\,
            I => \N__16149\
        );

    \I__3191\ : CascadeMux
    port map (
            O => \N__16152\,
            I => \N__16146\
        );

    \I__3190\ : CascadeBuf
    port map (
            O => \N__16149\,
            I => \N__16143\
        );

    \I__3189\ : CascadeBuf
    port map (
            O => \N__16146\,
            I => \N__16140\
        );

    \I__3188\ : CascadeMux
    port map (
            O => \N__16143\,
            I => \N__16137\
        );

    \I__3187\ : CascadeMux
    port map (
            O => \N__16140\,
            I => \N__16134\
        );

    \I__3186\ : CascadeBuf
    port map (
            O => \N__16137\,
            I => \N__16131\
        );

    \I__3185\ : CascadeBuf
    port map (
            O => \N__16134\,
            I => \N__16128\
        );

    \I__3184\ : CascadeMux
    port map (
            O => \N__16131\,
            I => \N__16125\
        );

    \I__3183\ : CascadeMux
    port map (
            O => \N__16128\,
            I => \N__16122\
        );

    \I__3182\ : InMux
    port map (
            O => \N__16125\,
            I => \N__16119\
        );

    \I__3181\ : InMux
    port map (
            O => \N__16122\,
            I => \N__16116\
        );

    \I__3180\ : LocalMux
    port map (
            O => \N__16119\,
            I => \N__16113\
        );

    \I__3179\ : LocalMux
    port map (
            O => \N__16116\,
            I => \N__16110\
        );

    \I__3178\ : Span4Mux_h
    port map (
            O => \N__16113\,
            I => \N__16107\
        );

    \I__3177\ : Span4Mux_h
    port map (
            O => \N__16110\,
            I => \N__16104\
        );

    \I__3176\ : Sp12to4
    port map (
            O => \N__16107\,
            I => \N__16101\
        );

    \I__3175\ : Sp12to4
    port map (
            O => \N__16104\,
            I => \N__16098\
        );

    \I__3174\ : Span12Mux_v
    port map (
            O => \N__16101\,
            I => \N__16093\
        );

    \I__3173\ : Span12Mux_v
    port map (
            O => \N__16098\,
            I => \N__16093\
        );

    \I__3172\ : Odrv12
    port map (
            O => \N__16093\,
            I => n19
        );

    \I__3171\ : InMux
    port map (
            O => \N__16090\,
            I => \N__16087\
        );

    \I__3170\ : LocalMux
    port map (
            O => \N__16087\,
            I => \transmit_module.X_DELTA_PATTERN_13\
        );

    \I__3169\ : InMux
    port map (
            O => \N__16084\,
            I => \N__16081\
        );

    \I__3168\ : LocalMux
    port map (
            O => \N__16081\,
            I => \transmit_module.X_DELTA_PATTERN_9\
        );

    \I__3167\ : InMux
    port map (
            O => \N__16078\,
            I => \N__16075\
        );

    \I__3166\ : LocalMux
    port map (
            O => \N__16075\,
            I => \transmit_module.X_DELTA_PATTERN_12\
        );

    \I__3165\ : InMux
    port map (
            O => \N__16072\,
            I => \N__16069\
        );

    \I__3164\ : LocalMux
    port map (
            O => \N__16069\,
            I => \transmit_module.X_DELTA_PATTERN_11\
        );

    \I__3163\ : InMux
    port map (
            O => \N__16066\,
            I => \N__16063\
        );

    \I__3162\ : LocalMux
    port map (
            O => \N__16063\,
            I => \transmit_module.X_DELTA_PATTERN_10\
        );

    \I__3161\ : InMux
    port map (
            O => \N__16060\,
            I => \N__16057\
        );

    \I__3160\ : LocalMux
    port map (
            O => \N__16057\,
            I => \N__16054\
        );

    \I__3159\ : Odrv12
    port map (
            O => \N__16054\,
            I => \line_buffer.n4072\
        );

    \I__3158\ : InMux
    port map (
            O => \N__16051\,
            I => \N__16048\
        );

    \I__3157\ : LocalMux
    port map (
            O => \N__16048\,
            I => \N__16045\
        );

    \I__3156\ : Span4Mux_v
    port map (
            O => \N__16045\,
            I => \N__16042\
        );

    \I__3155\ : Odrv4
    port map (
            O => \N__16042\,
            I => \line_buffer.n4134\
        );

    \I__3154\ : CEMux
    port map (
            O => \N__16039\,
            I => \N__16033\
        );

    \I__3153\ : CEMux
    port map (
            O => \N__16038\,
            I => \N__16030\
        );

    \I__3152\ : CEMux
    port map (
            O => \N__16037\,
            I => \N__16026\
        );

    \I__3151\ : CEMux
    port map (
            O => \N__16036\,
            I => \N__16022\
        );

    \I__3150\ : LocalMux
    port map (
            O => \N__16033\,
            I => \N__16019\
        );

    \I__3149\ : LocalMux
    port map (
            O => \N__16030\,
            I => \N__16016\
        );

    \I__3148\ : CEMux
    port map (
            O => \N__16029\,
            I => \N__16013\
        );

    \I__3147\ : LocalMux
    port map (
            O => \N__16026\,
            I => \N__16010\
        );

    \I__3146\ : SRMux
    port map (
            O => \N__16025\,
            I => \N__16007\
        );

    \I__3145\ : LocalMux
    port map (
            O => \N__16022\,
            I => \N__16004\
        );

    \I__3144\ : Span4Mux_h
    port map (
            O => \N__16019\,
            I => \N__16001\
        );

    \I__3143\ : Span4Mux_v
    port map (
            O => \N__16016\,
            I => \N__15996\
        );

    \I__3142\ : LocalMux
    port map (
            O => \N__16013\,
            I => \N__15996\
        );

    \I__3141\ : Span4Mux_v
    port map (
            O => \N__16010\,
            I => \N__15993\
        );

    \I__3140\ : LocalMux
    port map (
            O => \N__16007\,
            I => \N__15990\
        );

    \I__3139\ : Span4Mux_v
    port map (
            O => \N__16004\,
            I => \N__15983\
        );

    \I__3138\ : Span4Mux_v
    port map (
            O => \N__16001\,
            I => \N__15983\
        );

    \I__3137\ : Span4Mux_h
    port map (
            O => \N__15996\,
            I => \N__15983\
        );

    \I__3136\ : Span4Mux_h
    port map (
            O => \N__15993\,
            I => \N__15978\
        );

    \I__3135\ : Span4Mux_v
    port map (
            O => \N__15990\,
            I => \N__15978\
        );

    \I__3134\ : Odrv4
    port map (
            O => \N__15983\,
            I => \transmit_module.n2361\
        );

    \I__3133\ : Odrv4
    port map (
            O => \N__15978\,
            I => \transmit_module.n2361\
        );

    \I__3132\ : InMux
    port map (
            O => \N__15973\,
            I => \receive_module.rx_counter.n3722\
        );

    \I__3131\ : InMux
    port map (
            O => \N__15970\,
            I => \receive_module.rx_counter.n3723\
        );

    \I__3130\ : InMux
    port map (
            O => \N__15967\,
            I => \receive_module.rx_counter.n3724\
        );

    \I__3129\ : InMux
    port map (
            O => \N__15964\,
            I => \receive_module.rx_counter.n3725\
        );

    \I__3128\ : InMux
    port map (
            O => \N__15961\,
            I => \receive_module.rx_counter.n3726\
        );

    \I__3127\ : InMux
    port map (
            O => \N__15958\,
            I => \bfn_14_10_0_\
        );

    \I__3126\ : InMux
    port map (
            O => \N__15955\,
            I => \receive_module.rx_counter.n3728\
        );

    \I__3125\ : SRMux
    port map (
            O => \N__15952\,
            I => \N__15949\
        );

    \I__3124\ : LocalMux
    port map (
            O => \N__15949\,
            I => \N__15945\
        );

    \I__3123\ : SRMux
    port map (
            O => \N__15948\,
            I => \N__15942\
        );

    \I__3122\ : Span4Mux_v
    port map (
            O => \N__15945\,
            I => \N__15939\
        );

    \I__3121\ : LocalMux
    port map (
            O => \N__15942\,
            I => \N__15934\
        );

    \I__3120\ : Span4Mux_v
    port map (
            O => \N__15939\,
            I => \N__15934\
        );

    \I__3119\ : Odrv4
    port map (
            O => \N__15934\,
            I => n4214
        );

    \I__3118\ : CascadeMux
    port map (
            O => \N__15931\,
            I => \N__15924\
        );

    \I__3117\ : InMux
    port map (
            O => \N__15930\,
            I => \N__15918\
        );

    \I__3116\ : InMux
    port map (
            O => \N__15929\,
            I => \N__15915\
        );

    \I__3115\ : InMux
    port map (
            O => \N__15928\,
            I => \N__15908\
        );

    \I__3114\ : InMux
    port map (
            O => \N__15927\,
            I => \N__15908\
        );

    \I__3113\ : InMux
    port map (
            O => \N__15924\,
            I => \N__15908\
        );

    \I__3112\ : InMux
    port map (
            O => \N__15923\,
            I => \N__15901\
        );

    \I__3111\ : InMux
    port map (
            O => \N__15922\,
            I => \N__15901\
        );

    \I__3110\ : InMux
    port map (
            O => \N__15921\,
            I => \N__15901\
        );

    \I__3109\ : LocalMux
    port map (
            O => \N__15918\,
            I => \RX_ADDR_11\
        );

    \I__3108\ : LocalMux
    port map (
            O => \N__15915\,
            I => \RX_ADDR_11\
        );

    \I__3107\ : LocalMux
    port map (
            O => \N__15908\,
            I => \RX_ADDR_11\
        );

    \I__3106\ : LocalMux
    port map (
            O => \N__15901\,
            I => \RX_ADDR_11\
        );

    \I__3105\ : InMux
    port map (
            O => \N__15892\,
            I => \N__15882\
        );

    \I__3104\ : InMux
    port map (
            O => \N__15891\,
            I => \N__15879\
        );

    \I__3103\ : InMux
    port map (
            O => \N__15890\,
            I => \N__15872\
        );

    \I__3102\ : InMux
    port map (
            O => \N__15889\,
            I => \N__15872\
        );

    \I__3101\ : InMux
    port map (
            O => \N__15888\,
            I => \N__15872\
        );

    \I__3100\ : InMux
    port map (
            O => \N__15887\,
            I => \N__15865\
        );

    \I__3099\ : InMux
    port map (
            O => \N__15886\,
            I => \N__15865\
        );

    \I__3098\ : InMux
    port map (
            O => \N__15885\,
            I => \N__15865\
        );

    \I__3097\ : LocalMux
    port map (
            O => \N__15882\,
            I => \RX_ADDR_12\
        );

    \I__3096\ : LocalMux
    port map (
            O => \N__15879\,
            I => \RX_ADDR_12\
        );

    \I__3095\ : LocalMux
    port map (
            O => \N__15872\,
            I => \RX_ADDR_12\
        );

    \I__3094\ : LocalMux
    port map (
            O => \N__15865\,
            I => \RX_ADDR_12\
        );

    \I__3093\ : IoInMux
    port map (
            O => \N__15856\,
            I => \N__15853\
        );

    \I__3092\ : LocalMux
    port map (
            O => \N__15853\,
            I => \N__15849\
        );

    \I__3091\ : CascadeMux
    port map (
            O => \N__15852\,
            I => \N__15845\
        );

    \I__3090\ : Span4Mux_s2_h
    port map (
            O => \N__15849\,
            I => \N__15839\
        );

    \I__3089\ : CascadeMux
    port map (
            O => \N__15848\,
            I => \N__15836\
        );

    \I__3088\ : InMux
    port map (
            O => \N__15845\,
            I => \N__15833\
        );

    \I__3087\ : CascadeMux
    port map (
            O => \N__15844\,
            I => \N__15830\
        );

    \I__3086\ : CascadeMux
    port map (
            O => \N__15843\,
            I => \N__15827\
        );

    \I__3085\ : CascadeMux
    port map (
            O => \N__15842\,
            I => \N__15824\
        );

    \I__3084\ : Span4Mux_h
    port map (
            O => \N__15839\,
            I => \N__15821\
        );

    \I__3083\ : InMux
    port map (
            O => \N__15836\,
            I => \N__15818\
        );

    \I__3082\ : LocalMux
    port map (
            O => \N__15833\,
            I => \N__15815\
        );

    \I__3081\ : InMux
    port map (
            O => \N__15830\,
            I => \N__15808\
        );

    \I__3080\ : InMux
    port map (
            O => \N__15827\,
            I => \N__15808\
        );

    \I__3079\ : InMux
    port map (
            O => \N__15824\,
            I => \N__15808\
        );

    \I__3078\ : Span4Mux_h
    port map (
            O => \N__15821\,
            I => \N__15803\
        );

    \I__3077\ : LocalMux
    port map (
            O => \N__15818\,
            I => \N__15796\
        );

    \I__3076\ : Span4Mux_v
    port map (
            O => \N__15815\,
            I => \N__15796\
        );

    \I__3075\ : LocalMux
    port map (
            O => \N__15808\,
            I => \N__15796\
        );

    \I__3074\ : CascadeMux
    port map (
            O => \N__15807\,
            I => \N__15792\
        );

    \I__3073\ : CascadeMux
    port map (
            O => \N__15806\,
            I => \N__15789\
        );

    \I__3072\ : Sp12to4
    port map (
            O => \N__15803\,
            I => \N__15786\
        );

    \I__3071\ : Span4Mux_h
    port map (
            O => \N__15796\,
            I => \N__15783\
        );

    \I__3070\ : InMux
    port map (
            O => \N__15795\,
            I => \N__15776\
        );

    \I__3069\ : InMux
    port map (
            O => \N__15792\,
            I => \N__15776\
        );

    \I__3068\ : InMux
    port map (
            O => \N__15789\,
            I => \N__15776\
        );

    \I__3067\ : Odrv12
    port map (
            O => \N__15786\,
            I => \DEBUG_c_5\
        );

    \I__3066\ : Odrv4
    port map (
            O => \N__15783\,
            I => \DEBUG_c_5\
        );

    \I__3065\ : LocalMux
    port map (
            O => \N__15776\,
            I => \DEBUG_c_5\
        );

    \I__3064\ : IoInMux
    port map (
            O => \N__15769\,
            I => \N__15766\
        );

    \I__3063\ : LocalMux
    port map (
            O => \N__15766\,
            I => \N__15763\
        );

    \I__3062\ : Span12Mux_s9_h
    port map (
            O => \N__15763\,
            I => \N__15752\
        );

    \I__3061\ : InMux
    port map (
            O => \N__15762\,
            I => \N__15749\
        );

    \I__3060\ : InMux
    port map (
            O => \N__15761\,
            I => \N__15746\
        );

    \I__3059\ : InMux
    port map (
            O => \N__15760\,
            I => \N__15739\
        );

    \I__3058\ : InMux
    port map (
            O => \N__15759\,
            I => \N__15739\
        );

    \I__3057\ : InMux
    port map (
            O => \N__15758\,
            I => \N__15739\
        );

    \I__3056\ : InMux
    port map (
            O => \N__15757\,
            I => \N__15732\
        );

    \I__3055\ : InMux
    port map (
            O => \N__15756\,
            I => \N__15732\
        );

    \I__3054\ : InMux
    port map (
            O => \N__15755\,
            I => \N__15732\
        );

    \I__3053\ : Odrv12
    port map (
            O => \N__15752\,
            I => \DEBUG_c_3\
        );

    \I__3052\ : LocalMux
    port map (
            O => \N__15749\,
            I => \DEBUG_c_3\
        );

    \I__3051\ : LocalMux
    port map (
            O => \N__15746\,
            I => \DEBUG_c_3\
        );

    \I__3050\ : LocalMux
    port map (
            O => \N__15739\,
            I => \DEBUG_c_3\
        );

    \I__3049\ : LocalMux
    port map (
            O => \N__15732\,
            I => \DEBUG_c_3\
        );

    \I__3048\ : SRMux
    port map (
            O => \N__15721\,
            I => \N__15716\
        );

    \I__3047\ : SRMux
    port map (
            O => \N__15720\,
            I => \N__15713\
        );

    \I__3046\ : SRMux
    port map (
            O => \N__15719\,
            I => \N__15709\
        );

    \I__3045\ : LocalMux
    port map (
            O => \N__15716\,
            I => \N__15704\
        );

    \I__3044\ : LocalMux
    port map (
            O => \N__15713\,
            I => \N__15704\
        );

    \I__3043\ : SRMux
    port map (
            O => \N__15712\,
            I => \N__15701\
        );

    \I__3042\ : LocalMux
    port map (
            O => \N__15709\,
            I => \N__15698\
        );

    \I__3041\ : Span4Mux_v
    port map (
            O => \N__15704\,
            I => \N__15693\
        );

    \I__3040\ : LocalMux
    port map (
            O => \N__15701\,
            I => \N__15693\
        );

    \I__3039\ : Span4Mux_v
    port map (
            O => \N__15698\,
            I => \N__15690\
        );

    \I__3038\ : Span4Mux_h
    port map (
            O => \N__15693\,
            I => \N__15687\
        );

    \I__3037\ : Sp12to4
    port map (
            O => \N__15690\,
            I => \N__15684\
        );

    \I__3036\ : Span4Mux_h
    port map (
            O => \N__15687\,
            I => \N__15681\
        );

    \I__3035\ : Span12Mux_h
    port map (
            O => \N__15684\,
            I => \N__15678\
        );

    \I__3034\ : Span4Mux_h
    port map (
            O => \N__15681\,
            I => \N__15675\
        );

    \I__3033\ : Odrv12
    port map (
            O => \N__15678\,
            I => n658
        );

    \I__3032\ : Odrv4
    port map (
            O => \N__15675\,
            I => n658
        );

    \I__3031\ : CascadeMux
    port map (
            O => \N__15670\,
            I => \N__15667\
        );

    \I__3030\ : InMux
    port map (
            O => \N__15667\,
            I => \N__15664\
        );

    \I__3029\ : LocalMux
    port map (
            O => \N__15664\,
            I => \N__15661\
        );

    \I__3028\ : Span4Mux_v
    port map (
            O => \N__15661\,
            I => \N__15658\
        );

    \I__3027\ : Span4Mux_v
    port map (
            O => \N__15658\,
            I => \N__15655\
        );

    \I__3026\ : Odrv4
    port map (
            O => \N__15655\,
            I => \line_buffer.n4101\
        );

    \I__3025\ : CascadeMux
    port map (
            O => \N__15652\,
            I => \N__15649\
        );

    \I__3024\ : CascadeBuf
    port map (
            O => \N__15649\,
            I => \N__15645\
        );

    \I__3023\ : CascadeMux
    port map (
            O => \N__15648\,
            I => \N__15642\
        );

    \I__3022\ : CascadeMux
    port map (
            O => \N__15645\,
            I => \N__15639\
        );

    \I__3021\ : CascadeBuf
    port map (
            O => \N__15642\,
            I => \N__15636\
        );

    \I__3020\ : CascadeBuf
    port map (
            O => \N__15639\,
            I => \N__15633\
        );

    \I__3019\ : CascadeMux
    port map (
            O => \N__15636\,
            I => \N__15630\
        );

    \I__3018\ : CascadeMux
    port map (
            O => \N__15633\,
            I => \N__15627\
        );

    \I__3017\ : CascadeBuf
    port map (
            O => \N__15630\,
            I => \N__15624\
        );

    \I__3016\ : CascadeBuf
    port map (
            O => \N__15627\,
            I => \N__15621\
        );

    \I__3015\ : CascadeMux
    port map (
            O => \N__15624\,
            I => \N__15618\
        );

    \I__3014\ : CascadeMux
    port map (
            O => \N__15621\,
            I => \N__15615\
        );

    \I__3013\ : CascadeBuf
    port map (
            O => \N__15618\,
            I => \N__15612\
        );

    \I__3012\ : CascadeBuf
    port map (
            O => \N__15615\,
            I => \N__15609\
        );

    \I__3011\ : CascadeMux
    port map (
            O => \N__15612\,
            I => \N__15606\
        );

    \I__3010\ : CascadeMux
    port map (
            O => \N__15609\,
            I => \N__15603\
        );

    \I__3009\ : CascadeBuf
    port map (
            O => \N__15606\,
            I => \N__15600\
        );

    \I__3008\ : CascadeBuf
    port map (
            O => \N__15603\,
            I => \N__15597\
        );

    \I__3007\ : CascadeMux
    port map (
            O => \N__15600\,
            I => \N__15594\
        );

    \I__3006\ : CascadeMux
    port map (
            O => \N__15597\,
            I => \N__15591\
        );

    \I__3005\ : CascadeBuf
    port map (
            O => \N__15594\,
            I => \N__15588\
        );

    \I__3004\ : CascadeBuf
    port map (
            O => \N__15591\,
            I => \N__15585\
        );

    \I__3003\ : CascadeMux
    port map (
            O => \N__15588\,
            I => \N__15582\
        );

    \I__3002\ : CascadeMux
    port map (
            O => \N__15585\,
            I => \N__15579\
        );

    \I__3001\ : CascadeBuf
    port map (
            O => \N__15582\,
            I => \N__15576\
        );

    \I__3000\ : CascadeBuf
    port map (
            O => \N__15579\,
            I => \N__15573\
        );

    \I__2999\ : CascadeMux
    port map (
            O => \N__15576\,
            I => \N__15570\
        );

    \I__2998\ : CascadeMux
    port map (
            O => \N__15573\,
            I => \N__15567\
        );

    \I__2997\ : CascadeBuf
    port map (
            O => \N__15570\,
            I => \N__15564\
        );

    \I__2996\ : CascadeBuf
    port map (
            O => \N__15567\,
            I => \N__15561\
        );

    \I__2995\ : CascadeMux
    port map (
            O => \N__15564\,
            I => \N__15558\
        );

    \I__2994\ : CascadeMux
    port map (
            O => \N__15561\,
            I => \N__15555\
        );

    \I__2993\ : CascadeBuf
    port map (
            O => \N__15558\,
            I => \N__15552\
        );

    \I__2992\ : CascadeBuf
    port map (
            O => \N__15555\,
            I => \N__15549\
        );

    \I__2991\ : CascadeMux
    port map (
            O => \N__15552\,
            I => \N__15546\
        );

    \I__2990\ : CascadeMux
    port map (
            O => \N__15549\,
            I => \N__15543\
        );

    \I__2989\ : CascadeBuf
    port map (
            O => \N__15546\,
            I => \N__15540\
        );

    \I__2988\ : CascadeBuf
    port map (
            O => \N__15543\,
            I => \N__15537\
        );

    \I__2987\ : CascadeMux
    port map (
            O => \N__15540\,
            I => \N__15534\
        );

    \I__2986\ : CascadeMux
    port map (
            O => \N__15537\,
            I => \N__15531\
        );

    \I__2985\ : CascadeBuf
    port map (
            O => \N__15534\,
            I => \N__15528\
        );

    \I__2984\ : CascadeBuf
    port map (
            O => \N__15531\,
            I => \N__15525\
        );

    \I__2983\ : CascadeMux
    port map (
            O => \N__15528\,
            I => \N__15522\
        );

    \I__2982\ : CascadeMux
    port map (
            O => \N__15525\,
            I => \N__15519\
        );

    \I__2981\ : CascadeBuf
    port map (
            O => \N__15522\,
            I => \N__15516\
        );

    \I__2980\ : CascadeBuf
    port map (
            O => \N__15519\,
            I => \N__15513\
        );

    \I__2979\ : CascadeMux
    port map (
            O => \N__15516\,
            I => \N__15510\
        );

    \I__2978\ : CascadeMux
    port map (
            O => \N__15513\,
            I => \N__15507\
        );

    \I__2977\ : CascadeBuf
    port map (
            O => \N__15510\,
            I => \N__15504\
        );

    \I__2976\ : CascadeBuf
    port map (
            O => \N__15507\,
            I => \N__15501\
        );

    \I__2975\ : CascadeMux
    port map (
            O => \N__15504\,
            I => \N__15498\
        );

    \I__2974\ : CascadeMux
    port map (
            O => \N__15501\,
            I => \N__15495\
        );

    \I__2973\ : CascadeBuf
    port map (
            O => \N__15498\,
            I => \N__15492\
        );

    \I__2972\ : CascadeBuf
    port map (
            O => \N__15495\,
            I => \N__15489\
        );

    \I__2971\ : CascadeMux
    port map (
            O => \N__15492\,
            I => \N__15486\
        );

    \I__2970\ : CascadeMux
    port map (
            O => \N__15489\,
            I => \N__15483\
        );

    \I__2969\ : CascadeBuf
    port map (
            O => \N__15486\,
            I => \N__15480\
        );

    \I__2968\ : CascadeBuf
    port map (
            O => \N__15483\,
            I => \N__15477\
        );

    \I__2967\ : CascadeMux
    port map (
            O => \N__15480\,
            I => \N__15474\
        );

    \I__2966\ : CascadeMux
    port map (
            O => \N__15477\,
            I => \N__15471\
        );

    \I__2965\ : CascadeBuf
    port map (
            O => \N__15474\,
            I => \N__15468\
        );

    \I__2964\ : InMux
    port map (
            O => \N__15471\,
            I => \N__15465\
        );

    \I__2963\ : CascadeMux
    port map (
            O => \N__15468\,
            I => \N__15462\
        );

    \I__2962\ : LocalMux
    port map (
            O => \N__15465\,
            I => \N__15459\
        );

    \I__2961\ : InMux
    port map (
            O => \N__15462\,
            I => \N__15456\
        );

    \I__2960\ : Span12Mux_s10_h
    port map (
            O => \N__15459\,
            I => \N__15453\
        );

    \I__2959\ : LocalMux
    port map (
            O => \N__15456\,
            I => \N__15450\
        );

    \I__2958\ : Odrv12
    port map (
            O => \N__15453\,
            I => n22
        );

    \I__2957\ : Odrv12
    port map (
            O => \N__15450\,
            I => n22
        );

    \I__2956\ : CascadeMux
    port map (
            O => \N__15445\,
            I => \receive_module.rx_counter.n5_cascade_\
        );

    \I__2955\ : InMux
    port map (
            O => \N__15442\,
            I => \N__15435\
        );

    \I__2954\ : InMux
    port map (
            O => \N__15441\,
            I => \N__15435\
        );

    \I__2953\ : InMux
    port map (
            O => \N__15440\,
            I => \N__15432\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__15435\,
            I => \N__15429\
        );

    \I__2951\ : LocalMux
    port map (
            O => \N__15432\,
            I => \N__15426\
        );

    \I__2950\ : Span4Mux_h
    port map (
            O => \N__15429\,
            I => \N__15423\
        );

    \I__2949\ : Span4Mux_h
    port map (
            O => \N__15426\,
            I => \N__15420\
        );

    \I__2948\ : Span4Mux_h
    port map (
            O => \N__15423\,
            I => \N__15417\
        );

    \I__2947\ : Span4Mux_h
    port map (
            O => \N__15420\,
            I => \N__15414\
        );

    \I__2946\ : Sp12to4
    port map (
            O => \N__15417\,
            I => \N__15411\
        );

    \I__2945\ : Span4Mux_v
    port map (
            O => \N__15414\,
            I => \N__15408\
        );

    \I__2944\ : Odrv12
    port map (
            O => \N__15411\,
            I => \TVP_HSYNC_c\
        );

    \I__2943\ : Odrv4
    port map (
            O => \N__15408\,
            I => \TVP_HSYNC_c\
        );

    \I__2942\ : InMux
    port map (
            O => \N__15403\,
            I => \N__15400\
        );

    \I__2941\ : LocalMux
    port map (
            O => \N__15400\,
            I => \receive_module.rx_counter.n4_adj_576\
        );

    \I__2940\ : CascadeMux
    port map (
            O => \N__15397\,
            I => \N__15393\
        );

    \I__2939\ : CascadeMux
    port map (
            O => \N__15396\,
            I => \N__15390\
        );

    \I__2938\ : CascadeBuf
    port map (
            O => \N__15393\,
            I => \N__15387\
        );

    \I__2937\ : CascadeBuf
    port map (
            O => \N__15390\,
            I => \N__15384\
        );

    \I__2936\ : CascadeMux
    port map (
            O => \N__15387\,
            I => \N__15381\
        );

    \I__2935\ : CascadeMux
    port map (
            O => \N__15384\,
            I => \N__15378\
        );

    \I__2934\ : CascadeBuf
    port map (
            O => \N__15381\,
            I => \N__15375\
        );

    \I__2933\ : CascadeBuf
    port map (
            O => \N__15378\,
            I => \N__15372\
        );

    \I__2932\ : CascadeMux
    port map (
            O => \N__15375\,
            I => \N__15369\
        );

    \I__2931\ : CascadeMux
    port map (
            O => \N__15372\,
            I => \N__15366\
        );

    \I__2930\ : CascadeBuf
    port map (
            O => \N__15369\,
            I => \N__15363\
        );

    \I__2929\ : CascadeBuf
    port map (
            O => \N__15366\,
            I => \N__15360\
        );

    \I__2928\ : CascadeMux
    port map (
            O => \N__15363\,
            I => \N__15357\
        );

    \I__2927\ : CascadeMux
    port map (
            O => \N__15360\,
            I => \N__15354\
        );

    \I__2926\ : CascadeBuf
    port map (
            O => \N__15357\,
            I => \N__15351\
        );

    \I__2925\ : CascadeBuf
    port map (
            O => \N__15354\,
            I => \N__15348\
        );

    \I__2924\ : CascadeMux
    port map (
            O => \N__15351\,
            I => \N__15345\
        );

    \I__2923\ : CascadeMux
    port map (
            O => \N__15348\,
            I => \N__15342\
        );

    \I__2922\ : CascadeBuf
    port map (
            O => \N__15345\,
            I => \N__15339\
        );

    \I__2921\ : CascadeBuf
    port map (
            O => \N__15342\,
            I => \N__15336\
        );

    \I__2920\ : CascadeMux
    port map (
            O => \N__15339\,
            I => \N__15333\
        );

    \I__2919\ : CascadeMux
    port map (
            O => \N__15336\,
            I => \N__15330\
        );

    \I__2918\ : CascadeBuf
    port map (
            O => \N__15333\,
            I => \N__15327\
        );

    \I__2917\ : CascadeBuf
    port map (
            O => \N__15330\,
            I => \N__15324\
        );

    \I__2916\ : CascadeMux
    port map (
            O => \N__15327\,
            I => \N__15321\
        );

    \I__2915\ : CascadeMux
    port map (
            O => \N__15324\,
            I => \N__15318\
        );

    \I__2914\ : CascadeBuf
    port map (
            O => \N__15321\,
            I => \N__15315\
        );

    \I__2913\ : CascadeBuf
    port map (
            O => \N__15318\,
            I => \N__15312\
        );

    \I__2912\ : CascadeMux
    port map (
            O => \N__15315\,
            I => \N__15309\
        );

    \I__2911\ : CascadeMux
    port map (
            O => \N__15312\,
            I => \N__15306\
        );

    \I__2910\ : CascadeBuf
    port map (
            O => \N__15309\,
            I => \N__15303\
        );

    \I__2909\ : CascadeBuf
    port map (
            O => \N__15306\,
            I => \N__15300\
        );

    \I__2908\ : CascadeMux
    port map (
            O => \N__15303\,
            I => \N__15297\
        );

    \I__2907\ : CascadeMux
    port map (
            O => \N__15300\,
            I => \N__15294\
        );

    \I__2906\ : CascadeBuf
    port map (
            O => \N__15297\,
            I => \N__15291\
        );

    \I__2905\ : CascadeBuf
    port map (
            O => \N__15294\,
            I => \N__15288\
        );

    \I__2904\ : CascadeMux
    port map (
            O => \N__15291\,
            I => \N__15285\
        );

    \I__2903\ : CascadeMux
    port map (
            O => \N__15288\,
            I => \N__15282\
        );

    \I__2902\ : CascadeBuf
    port map (
            O => \N__15285\,
            I => \N__15279\
        );

    \I__2901\ : CascadeBuf
    port map (
            O => \N__15282\,
            I => \N__15276\
        );

    \I__2900\ : CascadeMux
    port map (
            O => \N__15279\,
            I => \N__15273\
        );

    \I__2899\ : CascadeMux
    port map (
            O => \N__15276\,
            I => \N__15270\
        );

    \I__2898\ : CascadeBuf
    port map (
            O => \N__15273\,
            I => \N__15267\
        );

    \I__2897\ : CascadeBuf
    port map (
            O => \N__15270\,
            I => \N__15264\
        );

    \I__2896\ : CascadeMux
    port map (
            O => \N__15267\,
            I => \N__15261\
        );

    \I__2895\ : CascadeMux
    port map (
            O => \N__15264\,
            I => \N__15258\
        );

    \I__2894\ : CascadeBuf
    port map (
            O => \N__15261\,
            I => \N__15255\
        );

    \I__2893\ : CascadeBuf
    port map (
            O => \N__15258\,
            I => \N__15252\
        );

    \I__2892\ : CascadeMux
    port map (
            O => \N__15255\,
            I => \N__15249\
        );

    \I__2891\ : CascadeMux
    port map (
            O => \N__15252\,
            I => \N__15246\
        );

    \I__2890\ : CascadeBuf
    port map (
            O => \N__15249\,
            I => \N__15243\
        );

    \I__2889\ : CascadeBuf
    port map (
            O => \N__15246\,
            I => \N__15240\
        );

    \I__2888\ : CascadeMux
    port map (
            O => \N__15243\,
            I => \N__15237\
        );

    \I__2887\ : CascadeMux
    port map (
            O => \N__15240\,
            I => \N__15234\
        );

    \I__2886\ : CascadeBuf
    port map (
            O => \N__15237\,
            I => \N__15231\
        );

    \I__2885\ : CascadeBuf
    port map (
            O => \N__15234\,
            I => \N__15228\
        );

    \I__2884\ : CascadeMux
    port map (
            O => \N__15231\,
            I => \N__15225\
        );

    \I__2883\ : CascadeMux
    port map (
            O => \N__15228\,
            I => \N__15222\
        );

    \I__2882\ : CascadeBuf
    port map (
            O => \N__15225\,
            I => \N__15219\
        );

    \I__2881\ : CascadeBuf
    port map (
            O => \N__15222\,
            I => \N__15216\
        );

    \I__2880\ : CascadeMux
    port map (
            O => \N__15219\,
            I => \N__15213\
        );

    \I__2879\ : CascadeMux
    port map (
            O => \N__15216\,
            I => \N__15210\
        );

    \I__2878\ : InMux
    port map (
            O => \N__15213\,
            I => \N__15207\
        );

    \I__2877\ : InMux
    port map (
            O => \N__15210\,
            I => \N__15204\
        );

    \I__2876\ : LocalMux
    port map (
            O => \N__15207\,
            I => \N__15201\
        );

    \I__2875\ : LocalMux
    port map (
            O => \N__15204\,
            I => \N__15198\
        );

    \I__2874\ : Span4Mux_s3_v
    port map (
            O => \N__15201\,
            I => \N__15195\
        );

    \I__2873\ : Span4Mux_s3_v
    port map (
            O => \N__15198\,
            I => \N__15192\
        );

    \I__2872\ : Sp12to4
    port map (
            O => \N__15195\,
            I => \N__15189\
        );

    \I__2871\ : Sp12to4
    port map (
            O => \N__15192\,
            I => \N__15186\
        );

    \I__2870\ : Span12Mux_h
    port map (
            O => \N__15189\,
            I => \N__15182\
        );

    \I__2869\ : Span12Mux_v
    port map (
            O => \N__15186\,
            I => \N__15179\
        );

    \I__2868\ : InMux
    port map (
            O => \N__15185\,
            I => \N__15176\
        );

    \I__2867\ : Span12Mux_v
    port map (
            O => \N__15182\,
            I => \N__15171\
        );

    \I__2866\ : Span12Mux_h
    port map (
            O => \N__15179\,
            I => \N__15171\
        );

    \I__2865\ : LocalMux
    port map (
            O => \N__15176\,
            I => \RX_ADDR_0\
        );

    \I__2864\ : Odrv12
    port map (
            O => \N__15171\,
            I => \RX_ADDR_0\
        );

    \I__2863\ : InMux
    port map (
            O => \N__15166\,
            I => \bfn_14_9_0_\
        );

    \I__2862\ : CascadeMux
    port map (
            O => \N__15163\,
            I => \N__15159\
        );

    \I__2861\ : CascadeMux
    port map (
            O => \N__15162\,
            I => \N__15156\
        );

    \I__2860\ : CascadeBuf
    port map (
            O => \N__15159\,
            I => \N__15153\
        );

    \I__2859\ : CascadeBuf
    port map (
            O => \N__15156\,
            I => \N__15150\
        );

    \I__2858\ : CascadeMux
    port map (
            O => \N__15153\,
            I => \N__15147\
        );

    \I__2857\ : CascadeMux
    port map (
            O => \N__15150\,
            I => \N__15144\
        );

    \I__2856\ : CascadeBuf
    port map (
            O => \N__15147\,
            I => \N__15141\
        );

    \I__2855\ : CascadeBuf
    port map (
            O => \N__15144\,
            I => \N__15138\
        );

    \I__2854\ : CascadeMux
    port map (
            O => \N__15141\,
            I => \N__15135\
        );

    \I__2853\ : CascadeMux
    port map (
            O => \N__15138\,
            I => \N__15132\
        );

    \I__2852\ : CascadeBuf
    port map (
            O => \N__15135\,
            I => \N__15129\
        );

    \I__2851\ : CascadeBuf
    port map (
            O => \N__15132\,
            I => \N__15126\
        );

    \I__2850\ : CascadeMux
    port map (
            O => \N__15129\,
            I => \N__15123\
        );

    \I__2849\ : CascadeMux
    port map (
            O => \N__15126\,
            I => \N__15120\
        );

    \I__2848\ : CascadeBuf
    port map (
            O => \N__15123\,
            I => \N__15117\
        );

    \I__2847\ : CascadeBuf
    port map (
            O => \N__15120\,
            I => \N__15114\
        );

    \I__2846\ : CascadeMux
    port map (
            O => \N__15117\,
            I => \N__15111\
        );

    \I__2845\ : CascadeMux
    port map (
            O => \N__15114\,
            I => \N__15108\
        );

    \I__2844\ : CascadeBuf
    port map (
            O => \N__15111\,
            I => \N__15105\
        );

    \I__2843\ : CascadeBuf
    port map (
            O => \N__15108\,
            I => \N__15102\
        );

    \I__2842\ : CascadeMux
    port map (
            O => \N__15105\,
            I => \N__15099\
        );

    \I__2841\ : CascadeMux
    port map (
            O => \N__15102\,
            I => \N__15096\
        );

    \I__2840\ : CascadeBuf
    port map (
            O => \N__15099\,
            I => \N__15093\
        );

    \I__2839\ : CascadeBuf
    port map (
            O => \N__15096\,
            I => \N__15090\
        );

    \I__2838\ : CascadeMux
    port map (
            O => \N__15093\,
            I => \N__15087\
        );

    \I__2837\ : CascadeMux
    port map (
            O => \N__15090\,
            I => \N__15084\
        );

    \I__2836\ : CascadeBuf
    port map (
            O => \N__15087\,
            I => \N__15081\
        );

    \I__2835\ : CascadeBuf
    port map (
            O => \N__15084\,
            I => \N__15078\
        );

    \I__2834\ : CascadeMux
    port map (
            O => \N__15081\,
            I => \N__15075\
        );

    \I__2833\ : CascadeMux
    port map (
            O => \N__15078\,
            I => \N__15072\
        );

    \I__2832\ : CascadeBuf
    port map (
            O => \N__15075\,
            I => \N__15069\
        );

    \I__2831\ : CascadeBuf
    port map (
            O => \N__15072\,
            I => \N__15066\
        );

    \I__2830\ : CascadeMux
    port map (
            O => \N__15069\,
            I => \N__15063\
        );

    \I__2829\ : CascadeMux
    port map (
            O => \N__15066\,
            I => \N__15060\
        );

    \I__2828\ : CascadeBuf
    port map (
            O => \N__15063\,
            I => \N__15057\
        );

    \I__2827\ : CascadeBuf
    port map (
            O => \N__15060\,
            I => \N__15054\
        );

    \I__2826\ : CascadeMux
    port map (
            O => \N__15057\,
            I => \N__15051\
        );

    \I__2825\ : CascadeMux
    port map (
            O => \N__15054\,
            I => \N__15048\
        );

    \I__2824\ : CascadeBuf
    port map (
            O => \N__15051\,
            I => \N__15045\
        );

    \I__2823\ : CascadeBuf
    port map (
            O => \N__15048\,
            I => \N__15042\
        );

    \I__2822\ : CascadeMux
    port map (
            O => \N__15045\,
            I => \N__15039\
        );

    \I__2821\ : CascadeMux
    port map (
            O => \N__15042\,
            I => \N__15036\
        );

    \I__2820\ : CascadeBuf
    port map (
            O => \N__15039\,
            I => \N__15033\
        );

    \I__2819\ : CascadeBuf
    port map (
            O => \N__15036\,
            I => \N__15030\
        );

    \I__2818\ : CascadeMux
    port map (
            O => \N__15033\,
            I => \N__15027\
        );

    \I__2817\ : CascadeMux
    port map (
            O => \N__15030\,
            I => \N__15024\
        );

    \I__2816\ : CascadeBuf
    port map (
            O => \N__15027\,
            I => \N__15021\
        );

    \I__2815\ : CascadeBuf
    port map (
            O => \N__15024\,
            I => \N__15018\
        );

    \I__2814\ : CascadeMux
    port map (
            O => \N__15021\,
            I => \N__15015\
        );

    \I__2813\ : CascadeMux
    port map (
            O => \N__15018\,
            I => \N__15012\
        );

    \I__2812\ : CascadeBuf
    port map (
            O => \N__15015\,
            I => \N__15009\
        );

    \I__2811\ : CascadeBuf
    port map (
            O => \N__15012\,
            I => \N__15006\
        );

    \I__2810\ : CascadeMux
    port map (
            O => \N__15009\,
            I => \N__15003\
        );

    \I__2809\ : CascadeMux
    port map (
            O => \N__15006\,
            I => \N__15000\
        );

    \I__2808\ : CascadeBuf
    port map (
            O => \N__15003\,
            I => \N__14997\
        );

    \I__2807\ : CascadeBuf
    port map (
            O => \N__15000\,
            I => \N__14994\
        );

    \I__2806\ : CascadeMux
    port map (
            O => \N__14997\,
            I => \N__14991\
        );

    \I__2805\ : CascadeMux
    port map (
            O => \N__14994\,
            I => \N__14988\
        );

    \I__2804\ : CascadeBuf
    port map (
            O => \N__14991\,
            I => \N__14985\
        );

    \I__2803\ : CascadeBuf
    port map (
            O => \N__14988\,
            I => \N__14982\
        );

    \I__2802\ : CascadeMux
    port map (
            O => \N__14985\,
            I => \N__14979\
        );

    \I__2801\ : CascadeMux
    port map (
            O => \N__14982\,
            I => \N__14976\
        );

    \I__2800\ : InMux
    port map (
            O => \N__14979\,
            I => \N__14973\
        );

    \I__2799\ : InMux
    port map (
            O => \N__14976\,
            I => \N__14970\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__14973\,
            I => \N__14967\
        );

    \I__2797\ : LocalMux
    port map (
            O => \N__14970\,
            I => \N__14964\
        );

    \I__2796\ : Span4Mux_s2_v
    port map (
            O => \N__14967\,
            I => \N__14961\
        );

    \I__2795\ : Sp12to4
    port map (
            O => \N__14964\,
            I => \N__14958\
        );

    \I__2794\ : Sp12to4
    port map (
            O => \N__14961\,
            I => \N__14955\
        );

    \I__2793\ : Span12Mux_s11_v
    port map (
            O => \N__14958\,
            I => \N__14951\
        );

    \I__2792\ : Span12Mux_h
    port map (
            O => \N__14955\,
            I => \N__14948\
        );

    \I__2791\ : InMux
    port map (
            O => \N__14954\,
            I => \N__14945\
        );

    \I__2790\ : Span12Mux_v
    port map (
            O => \N__14951\,
            I => \N__14942\
        );

    \I__2789\ : Span12Mux_v
    port map (
            O => \N__14948\,
            I => \N__14939\
        );

    \I__2788\ : LocalMux
    port map (
            O => \N__14945\,
            I => \RX_ADDR_1\
        );

    \I__2787\ : Odrv12
    port map (
            O => \N__14942\,
            I => \RX_ADDR_1\
        );

    \I__2786\ : Odrv12
    port map (
            O => \N__14939\,
            I => \RX_ADDR_1\
        );

    \I__2785\ : InMux
    port map (
            O => \N__14932\,
            I => \receive_module.rx_counter.n3720\
        );

    \I__2784\ : CascadeMux
    port map (
            O => \N__14929\,
            I => \N__14926\
        );

    \I__2783\ : CascadeBuf
    port map (
            O => \N__14926\,
            I => \N__14922\
        );

    \I__2782\ : CascadeMux
    port map (
            O => \N__14925\,
            I => \N__14919\
        );

    \I__2781\ : CascadeMux
    port map (
            O => \N__14922\,
            I => \N__14916\
        );

    \I__2780\ : CascadeBuf
    port map (
            O => \N__14919\,
            I => \N__14913\
        );

    \I__2779\ : CascadeBuf
    port map (
            O => \N__14916\,
            I => \N__14910\
        );

    \I__2778\ : CascadeMux
    port map (
            O => \N__14913\,
            I => \N__14907\
        );

    \I__2777\ : CascadeMux
    port map (
            O => \N__14910\,
            I => \N__14904\
        );

    \I__2776\ : CascadeBuf
    port map (
            O => \N__14907\,
            I => \N__14901\
        );

    \I__2775\ : CascadeBuf
    port map (
            O => \N__14904\,
            I => \N__14898\
        );

    \I__2774\ : CascadeMux
    port map (
            O => \N__14901\,
            I => \N__14895\
        );

    \I__2773\ : CascadeMux
    port map (
            O => \N__14898\,
            I => \N__14892\
        );

    \I__2772\ : CascadeBuf
    port map (
            O => \N__14895\,
            I => \N__14889\
        );

    \I__2771\ : CascadeBuf
    port map (
            O => \N__14892\,
            I => \N__14886\
        );

    \I__2770\ : CascadeMux
    port map (
            O => \N__14889\,
            I => \N__14883\
        );

    \I__2769\ : CascadeMux
    port map (
            O => \N__14886\,
            I => \N__14880\
        );

    \I__2768\ : CascadeBuf
    port map (
            O => \N__14883\,
            I => \N__14877\
        );

    \I__2767\ : CascadeBuf
    port map (
            O => \N__14880\,
            I => \N__14874\
        );

    \I__2766\ : CascadeMux
    port map (
            O => \N__14877\,
            I => \N__14871\
        );

    \I__2765\ : CascadeMux
    port map (
            O => \N__14874\,
            I => \N__14868\
        );

    \I__2764\ : CascadeBuf
    port map (
            O => \N__14871\,
            I => \N__14865\
        );

    \I__2763\ : CascadeBuf
    port map (
            O => \N__14868\,
            I => \N__14862\
        );

    \I__2762\ : CascadeMux
    port map (
            O => \N__14865\,
            I => \N__14859\
        );

    \I__2761\ : CascadeMux
    port map (
            O => \N__14862\,
            I => \N__14856\
        );

    \I__2760\ : CascadeBuf
    port map (
            O => \N__14859\,
            I => \N__14853\
        );

    \I__2759\ : CascadeBuf
    port map (
            O => \N__14856\,
            I => \N__14850\
        );

    \I__2758\ : CascadeMux
    port map (
            O => \N__14853\,
            I => \N__14847\
        );

    \I__2757\ : CascadeMux
    port map (
            O => \N__14850\,
            I => \N__14844\
        );

    \I__2756\ : CascadeBuf
    port map (
            O => \N__14847\,
            I => \N__14841\
        );

    \I__2755\ : CascadeBuf
    port map (
            O => \N__14844\,
            I => \N__14838\
        );

    \I__2754\ : CascadeMux
    port map (
            O => \N__14841\,
            I => \N__14835\
        );

    \I__2753\ : CascadeMux
    port map (
            O => \N__14838\,
            I => \N__14832\
        );

    \I__2752\ : CascadeBuf
    port map (
            O => \N__14835\,
            I => \N__14829\
        );

    \I__2751\ : CascadeBuf
    port map (
            O => \N__14832\,
            I => \N__14826\
        );

    \I__2750\ : CascadeMux
    port map (
            O => \N__14829\,
            I => \N__14823\
        );

    \I__2749\ : CascadeMux
    port map (
            O => \N__14826\,
            I => \N__14820\
        );

    \I__2748\ : CascadeBuf
    port map (
            O => \N__14823\,
            I => \N__14817\
        );

    \I__2747\ : CascadeBuf
    port map (
            O => \N__14820\,
            I => \N__14814\
        );

    \I__2746\ : CascadeMux
    port map (
            O => \N__14817\,
            I => \N__14811\
        );

    \I__2745\ : CascadeMux
    port map (
            O => \N__14814\,
            I => \N__14808\
        );

    \I__2744\ : CascadeBuf
    port map (
            O => \N__14811\,
            I => \N__14805\
        );

    \I__2743\ : CascadeBuf
    port map (
            O => \N__14808\,
            I => \N__14802\
        );

    \I__2742\ : CascadeMux
    port map (
            O => \N__14805\,
            I => \N__14799\
        );

    \I__2741\ : CascadeMux
    port map (
            O => \N__14802\,
            I => \N__14796\
        );

    \I__2740\ : CascadeBuf
    port map (
            O => \N__14799\,
            I => \N__14793\
        );

    \I__2739\ : CascadeBuf
    port map (
            O => \N__14796\,
            I => \N__14790\
        );

    \I__2738\ : CascadeMux
    port map (
            O => \N__14793\,
            I => \N__14787\
        );

    \I__2737\ : CascadeMux
    port map (
            O => \N__14790\,
            I => \N__14784\
        );

    \I__2736\ : CascadeBuf
    port map (
            O => \N__14787\,
            I => \N__14781\
        );

    \I__2735\ : CascadeBuf
    port map (
            O => \N__14784\,
            I => \N__14778\
        );

    \I__2734\ : CascadeMux
    port map (
            O => \N__14781\,
            I => \N__14775\
        );

    \I__2733\ : CascadeMux
    port map (
            O => \N__14778\,
            I => \N__14772\
        );

    \I__2732\ : CascadeBuf
    port map (
            O => \N__14775\,
            I => \N__14769\
        );

    \I__2731\ : CascadeBuf
    port map (
            O => \N__14772\,
            I => \N__14766\
        );

    \I__2730\ : CascadeMux
    port map (
            O => \N__14769\,
            I => \N__14763\
        );

    \I__2729\ : CascadeMux
    port map (
            O => \N__14766\,
            I => \N__14760\
        );

    \I__2728\ : CascadeBuf
    port map (
            O => \N__14763\,
            I => \N__14757\
        );

    \I__2727\ : CascadeBuf
    port map (
            O => \N__14760\,
            I => \N__14754\
        );

    \I__2726\ : CascadeMux
    port map (
            O => \N__14757\,
            I => \N__14751\
        );

    \I__2725\ : CascadeMux
    port map (
            O => \N__14754\,
            I => \N__14748\
        );

    \I__2724\ : CascadeBuf
    port map (
            O => \N__14751\,
            I => \N__14745\
        );

    \I__2723\ : InMux
    port map (
            O => \N__14748\,
            I => \N__14742\
        );

    \I__2722\ : CascadeMux
    port map (
            O => \N__14745\,
            I => \N__14739\
        );

    \I__2721\ : LocalMux
    port map (
            O => \N__14742\,
            I => \N__14736\
        );

    \I__2720\ : InMux
    port map (
            O => \N__14739\,
            I => \N__14733\
        );

    \I__2719\ : Span4Mux_s3_v
    port map (
            O => \N__14736\,
            I => \N__14730\
        );

    \I__2718\ : LocalMux
    port map (
            O => \N__14733\,
            I => \N__14727\
        );

    \I__2717\ : Sp12to4
    port map (
            O => \N__14730\,
            I => \N__14724\
        );

    \I__2716\ : Span12Mux_s11_v
    port map (
            O => \N__14727\,
            I => \N__14720\
        );

    \I__2715\ : Span12Mux_v
    port map (
            O => \N__14724\,
            I => \N__14717\
        );

    \I__2714\ : InMux
    port map (
            O => \N__14723\,
            I => \N__14714\
        );

    \I__2713\ : Span12Mux_v
    port map (
            O => \N__14720\,
            I => \N__14711\
        );

    \I__2712\ : Span12Mux_h
    port map (
            O => \N__14717\,
            I => \N__14708\
        );

    \I__2711\ : LocalMux
    port map (
            O => \N__14714\,
            I => \RX_ADDR_2\
        );

    \I__2710\ : Odrv12
    port map (
            O => \N__14711\,
            I => \RX_ADDR_2\
        );

    \I__2709\ : Odrv12
    port map (
            O => \N__14708\,
            I => \RX_ADDR_2\
        );

    \I__2708\ : InMux
    port map (
            O => \N__14701\,
            I => \receive_module.rx_counter.n3721\
        );

    \I__2707\ : InMux
    port map (
            O => \N__14698\,
            I => \N__14695\
        );

    \I__2706\ : LocalMux
    port map (
            O => \N__14695\,
            I => \transmit_module.Y_DELTA_PATTERN_49\
        );

    \I__2705\ : InMux
    port map (
            O => \N__14692\,
            I => \N__14689\
        );

    \I__2704\ : LocalMux
    port map (
            O => \N__14689\,
            I => \transmit_module.Y_DELTA_PATTERN_54\
        );

    \I__2703\ : InMux
    port map (
            O => \N__14686\,
            I => \N__14683\
        );

    \I__2702\ : LocalMux
    port map (
            O => \N__14683\,
            I => \transmit_module.Y_DELTA_PATTERN_51\
        );

    \I__2701\ : InMux
    port map (
            O => \N__14680\,
            I => \N__14677\
        );

    \I__2700\ : LocalMux
    port map (
            O => \N__14677\,
            I => \transmit_module.Y_DELTA_PATTERN_50\
        );

    \I__2699\ : InMux
    port map (
            O => \N__14674\,
            I => \N__14671\
        );

    \I__2698\ : LocalMux
    port map (
            O => \N__14671\,
            I => \transmit_module.Y_DELTA_PATTERN_56\
        );

    \I__2697\ : InMux
    port map (
            O => \N__14668\,
            I => \N__14665\
        );

    \I__2696\ : LocalMux
    port map (
            O => \N__14665\,
            I => \transmit_module.Y_DELTA_PATTERN_55\
        );

    \I__2695\ : InMux
    port map (
            O => \N__14662\,
            I => \N__14659\
        );

    \I__2694\ : LocalMux
    port map (
            O => \N__14659\,
            I => \transmit_module.Y_DELTA_PATTERN_59\
        );

    \I__2693\ : InMux
    port map (
            O => \N__14656\,
            I => \N__14653\
        );

    \I__2692\ : LocalMux
    port map (
            O => \N__14653\,
            I => \transmit_module.Y_DELTA_PATTERN_58\
        );

    \I__2691\ : InMux
    port map (
            O => \N__14650\,
            I => \N__14647\
        );

    \I__2690\ : LocalMux
    port map (
            O => \N__14647\,
            I => \transmit_module.Y_DELTA_PATTERN_61\
        );

    \I__2689\ : InMux
    port map (
            O => \N__14644\,
            I => \N__14641\
        );

    \I__2688\ : LocalMux
    port map (
            O => \N__14641\,
            I => \transmit_module.Y_DELTA_PATTERN_60\
        );

    \I__2687\ : InMux
    port map (
            O => \N__14638\,
            I => \N__14635\
        );

    \I__2686\ : LocalMux
    port map (
            O => \N__14635\,
            I => \N__14632\
        );

    \I__2685\ : Span4Mux_h
    port map (
            O => \N__14632\,
            I => \N__14629\
        );

    \I__2684\ : Span4Mux_h
    port map (
            O => \N__14629\,
            I => \N__14626\
        );

    \I__2683\ : Span4Mux_h
    port map (
            O => \N__14626\,
            I => \N__14623\
        );

    \I__2682\ : Odrv4
    port map (
            O => \N__14623\,
            I => \line_buffer.n558\
        );

    \I__2681\ : InMux
    port map (
            O => \N__14620\,
            I => \N__14617\
        );

    \I__2680\ : LocalMux
    port map (
            O => \N__14617\,
            I => \N__14614\
        );

    \I__2679\ : Span4Mux_v
    port map (
            O => \N__14614\,
            I => \N__14611\
        );

    \I__2678\ : Span4Mux_h
    port map (
            O => \N__14611\,
            I => \N__14608\
        );

    \I__2677\ : Odrv4
    port map (
            O => \N__14608\,
            I => \line_buffer.n550\
        );

    \I__2676\ : SRMux
    port map (
            O => \N__14605\,
            I => \N__14601\
        );

    \I__2675\ : SRMux
    port map (
            O => \N__14604\,
            I => \N__14598\
        );

    \I__2674\ : LocalMux
    port map (
            O => \N__14601\,
            I => \N__14595\
        );

    \I__2673\ : LocalMux
    port map (
            O => \N__14598\,
            I => \N__14592\
        );

    \I__2672\ : Odrv4
    port map (
            O => \N__14595\,
            I => n2587
        );

    \I__2671\ : Odrv4
    port map (
            O => \N__14592\,
            I => n2587
        );

    \I__2670\ : InMux
    port map (
            O => \N__14587\,
            I => \N__14584\
        );

    \I__2669\ : LocalMux
    port map (
            O => \N__14584\,
            I => \transmit_module.Y_DELTA_PATTERN_43\
        );

    \I__2668\ : InMux
    port map (
            O => \N__14581\,
            I => \N__14578\
        );

    \I__2667\ : LocalMux
    port map (
            O => \N__14578\,
            I => \transmit_module.Y_DELTA_PATTERN_44\
        );

    \I__2666\ : InMux
    port map (
            O => \N__14575\,
            I => \N__14572\
        );

    \I__2665\ : LocalMux
    port map (
            O => \N__14572\,
            I => \transmit_module.Y_DELTA_PATTERN_46\
        );

    \I__2664\ : InMux
    port map (
            O => \N__14569\,
            I => \N__14566\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__14566\,
            I => \transmit_module.Y_DELTA_PATTERN_45\
        );

    \I__2662\ : InMux
    port map (
            O => \N__14563\,
            I => \N__14560\
        );

    \I__2661\ : LocalMux
    port map (
            O => \N__14560\,
            I => \transmit_module.Y_DELTA_PATTERN_47\
        );

    \I__2660\ : InMux
    port map (
            O => \N__14557\,
            I => \N__14554\
        );

    \I__2659\ : LocalMux
    port map (
            O => \N__14554\,
            I => \transmit_module.Y_DELTA_PATTERN_48\
        );

    \I__2658\ : InMux
    port map (
            O => \N__14551\,
            I => \N__14548\
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__14548\,
            I => \transmit_module.Y_DELTA_PATTERN_53\
        );

    \I__2656\ : InMux
    port map (
            O => \N__14545\,
            I => \N__14542\
        );

    \I__2655\ : LocalMux
    port map (
            O => \N__14542\,
            I => \transmit_module.Y_DELTA_PATTERN_52\
        );

    \I__2654\ : CascadeMux
    port map (
            O => \N__14539\,
            I => \line_buffer.n4185_cascade_\
        );

    \I__2653\ : InMux
    port map (
            O => \N__14536\,
            I => \N__14533\
        );

    \I__2652\ : LocalMux
    port map (
            O => \N__14533\,
            I => \N__14530\
        );

    \I__2651\ : Span4Mux_v
    port map (
            O => \N__14530\,
            I => \N__14527\
        );

    \I__2650\ : Odrv4
    port map (
            O => \N__14527\,
            I => \line_buffer.n4125\
        );

    \I__2649\ : IoInMux
    port map (
            O => \N__14524\,
            I => \N__14521\
        );

    \I__2648\ : LocalMux
    port map (
            O => \N__14521\,
            I => \N__14517\
        );

    \I__2647\ : IoInMux
    port map (
            O => \N__14520\,
            I => \N__14514\
        );

    \I__2646\ : IoSpan4Mux
    port map (
            O => \N__14517\,
            I => \N__14508\
        );

    \I__2645\ : LocalMux
    port map (
            O => \N__14514\,
            I => \N__14508\
        );

    \I__2644\ : IoInMux
    port map (
            O => \N__14513\,
            I => \N__14505\
        );

    \I__2643\ : IoSpan4Mux
    port map (
            O => \N__14508\,
            I => \N__14502\
        );

    \I__2642\ : LocalMux
    port map (
            O => \N__14505\,
            I => \N__14499\
        );

    \I__2641\ : Span4Mux_s0_h
    port map (
            O => \N__14502\,
            I => \N__14496\
        );

    \I__2640\ : Span4Mux_s3_v
    port map (
            O => \N__14499\,
            I => \N__14493\
        );

    \I__2639\ : Sp12to4
    port map (
            O => \N__14496\,
            I => \N__14490\
        );

    \I__2638\ : Sp12to4
    port map (
            O => \N__14493\,
            I => \N__14487\
        );

    \I__2637\ : Span12Mux_h
    port map (
            O => \N__14490\,
            I => \N__14482\
        );

    \I__2636\ : Span12Mux_h
    port map (
            O => \N__14487\,
            I => \N__14482\
        );

    \I__2635\ : Odrv12
    port map (
            O => \N__14482\,
            I => n1995
        );

    \I__2634\ : InMux
    port map (
            O => \N__14479\,
            I => \N__14476\
        );

    \I__2633\ : LocalMux
    port map (
            O => \N__14476\,
            I => \N__14473\
        );

    \I__2632\ : Span4Mux_h
    port map (
            O => \N__14473\,
            I => \N__14470\
        );

    \I__2631\ : Span4Mux_v
    port map (
            O => \N__14470\,
            I => \N__14467\
        );

    \I__2630\ : Odrv4
    port map (
            O => \N__14467\,
            I => \TX_DATA_2\
        );

    \I__2629\ : IoInMux
    port map (
            O => \N__14464\,
            I => \N__14459\
        );

    \I__2628\ : IoInMux
    port map (
            O => \N__14463\,
            I => \N__14456\
        );

    \I__2627\ : IoInMux
    port map (
            O => \N__14462\,
            I => \N__14453\
        );

    \I__2626\ : LocalMux
    port map (
            O => \N__14459\,
            I => \N__14450\
        );

    \I__2625\ : LocalMux
    port map (
            O => \N__14456\,
            I => \N__14447\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__14453\,
            I => \N__14444\
        );

    \I__2623\ : Span4Mux_s2_v
    port map (
            O => \N__14450\,
            I => \N__14441\
        );

    \I__2622\ : Span4Mux_s2_v
    port map (
            O => \N__14447\,
            I => \N__14438\
        );

    \I__2621\ : IoSpan4Mux
    port map (
            O => \N__14444\,
            I => \N__14435\
        );

    \I__2620\ : Sp12to4
    port map (
            O => \N__14441\,
            I => \N__14432\
        );

    \I__2619\ : Sp12to4
    port map (
            O => \N__14438\,
            I => \N__14429\
        );

    \I__2618\ : Sp12to4
    port map (
            O => \N__14435\,
            I => \N__14426\
        );

    \I__2617\ : Span12Mux_h
    port map (
            O => \N__14432\,
            I => \N__14419\
        );

    \I__2616\ : Span12Mux_h
    port map (
            O => \N__14429\,
            I => \N__14419\
        );

    \I__2615\ : Span12Mux_h
    port map (
            O => \N__14426\,
            I => \N__14419\
        );

    \I__2614\ : Odrv12
    port map (
            O => \N__14419\,
            I => n1994
        );

    \I__2613\ : IoInMux
    port map (
            O => \N__14416\,
            I => \N__14412\
        );

    \I__2612\ : IoInMux
    port map (
            O => \N__14415\,
            I => \N__14408\
        );

    \I__2611\ : LocalMux
    port map (
            O => \N__14412\,
            I => \N__14405\
        );

    \I__2610\ : IoInMux
    port map (
            O => \N__14411\,
            I => \N__14402\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__14408\,
            I => \N__14399\
        );

    \I__2608\ : IoSpan4Mux
    port map (
            O => \N__14405\,
            I => \N__14396\
        );

    \I__2607\ : LocalMux
    port map (
            O => \N__14402\,
            I => \N__14393\
        );

    \I__2606\ : IoSpan4Mux
    port map (
            O => \N__14399\,
            I => \N__14390\
        );

    \I__2605\ : Sp12to4
    port map (
            O => \N__14396\,
            I => \N__14387\
        );

    \I__2604\ : IoSpan4Mux
    port map (
            O => \N__14393\,
            I => \N__14384\
        );

    \I__2603\ : Span4Mux_s3_h
    port map (
            O => \N__14390\,
            I => \N__14381\
        );

    \I__2602\ : Span12Mux_v
    port map (
            O => \N__14387\,
            I => \N__14378\
        );

    \I__2601\ : Sp12to4
    port map (
            O => \N__14384\,
            I => \N__14375\
        );

    \I__2600\ : Span4Mux_h
    port map (
            O => \N__14381\,
            I => \N__14372\
        );

    \I__2599\ : Span12Mux_h
    port map (
            O => \N__14378\,
            I => \N__14367\
        );

    \I__2598\ : Span12Mux_v
    port map (
            O => \N__14375\,
            I => \N__14367\
        );

    \I__2597\ : Span4Mux_h
    port map (
            O => \N__14372\,
            I => \N__14364\
        );

    \I__2596\ : Odrv12
    port map (
            O => \N__14367\,
            I => n1993
        );

    \I__2595\ : Odrv4
    port map (
            O => \N__14364\,
            I => n1993
        );

    \I__2594\ : IoInMux
    port map (
            O => \N__14359\,
            I => \N__14356\
        );

    \I__2593\ : LocalMux
    port map (
            O => \N__14356\,
            I => \N__14353\
        );

    \I__2592\ : Span4Mux_s0_v
    port map (
            O => \N__14353\,
            I => \N__14348\
        );

    \I__2591\ : IoInMux
    port map (
            O => \N__14352\,
            I => \N__14345\
        );

    \I__2590\ : IoInMux
    port map (
            O => \N__14351\,
            I => \N__14342\
        );

    \I__2589\ : Span4Mux_v
    port map (
            O => \N__14348\,
            I => \N__14339\
        );

    \I__2588\ : LocalMux
    port map (
            O => \N__14345\,
            I => \N__14336\
        );

    \I__2587\ : LocalMux
    port map (
            O => \N__14342\,
            I => \N__14333\
        );

    \I__2586\ : Span4Mux_v
    port map (
            O => \N__14339\,
            I => \N__14330\
        );

    \I__2585\ : IoSpan4Mux
    port map (
            O => \N__14336\,
            I => \N__14327\
        );

    \I__2584\ : Span12Mux_s0_v
    port map (
            O => \N__14333\,
            I => \N__14324\
        );

    \I__2583\ : Sp12to4
    port map (
            O => \N__14330\,
            I => \N__14321\
        );

    \I__2582\ : Sp12to4
    port map (
            O => \N__14327\,
            I => \N__14318\
        );

    \I__2581\ : Span12Mux_v
    port map (
            O => \N__14324\,
            I => \N__14315\
        );

    \I__2580\ : Span12Mux_h
    port map (
            O => \N__14321\,
            I => \N__14310\
        );

    \I__2579\ : Span12Mux_h
    port map (
            O => \N__14318\,
            I => \N__14310\
        );

    \I__2578\ : Odrv12
    port map (
            O => \N__14315\,
            I => n1992
        );

    \I__2577\ : Odrv12
    port map (
            O => \N__14310\,
            I => n1992
        );

    \I__2576\ : IoInMux
    port map (
            O => \N__14305\,
            I => \N__14301\
        );

    \I__2575\ : IoInMux
    port map (
            O => \N__14304\,
            I => \N__14297\
        );

    \I__2574\ : LocalMux
    port map (
            O => \N__14301\,
            I => \N__14294\
        );

    \I__2573\ : IoInMux
    port map (
            O => \N__14300\,
            I => \N__14291\
        );

    \I__2572\ : LocalMux
    port map (
            O => \N__14297\,
            I => \N__14288\
        );

    \I__2571\ : Sp12to4
    port map (
            O => \N__14294\,
            I => \N__14285\
        );

    \I__2570\ : LocalMux
    port map (
            O => \N__14291\,
            I => \N__14282\
        );

    \I__2569\ : IoSpan4Mux
    port map (
            O => \N__14288\,
            I => \N__14279\
        );

    \I__2568\ : Span12Mux_v
    port map (
            O => \N__14285\,
            I => \N__14276\
        );

    \I__2567\ : Span12Mux_s0_h
    port map (
            O => \N__14282\,
            I => \N__14273\
        );

    \I__2566\ : Sp12to4
    port map (
            O => \N__14279\,
            I => \N__14270\
        );

    \I__2565\ : Span12Mux_h
    port map (
            O => \N__14276\,
            I => \N__14267\
        );

    \I__2564\ : Span12Mux_h
    port map (
            O => \N__14273\,
            I => \N__14264\
        );

    \I__2563\ : Span12Mux_v
    port map (
            O => \N__14270\,
            I => \N__14261\
        );

    \I__2562\ : Odrv12
    port map (
            O => \N__14267\,
            I => n1991
        );

    \I__2561\ : Odrv12
    port map (
            O => \N__14264\,
            I => n1991
        );

    \I__2560\ : Odrv12
    port map (
            O => \N__14261\,
            I => n1991
        );

    \I__2559\ : InMux
    port map (
            O => \N__14254\,
            I => \N__14251\
        );

    \I__2558\ : LocalMux
    port map (
            O => \N__14251\,
            I => \N__14248\
        );

    \I__2557\ : Odrv4
    port map (
            O => \N__14248\,
            I => \TX_DATA_6\
        );

    \I__2556\ : IoInMux
    port map (
            O => \N__14245\,
            I => \N__14240\
        );

    \I__2555\ : IoInMux
    port map (
            O => \N__14244\,
            I => \N__14237\
        );

    \I__2554\ : IoInMux
    port map (
            O => \N__14243\,
            I => \N__14234\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__14240\,
            I => \N__14231\
        );

    \I__2552\ : LocalMux
    port map (
            O => \N__14237\,
            I => \N__14228\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__14234\,
            I => \N__14225\
        );

    \I__2550\ : Span4Mux_s0_v
    port map (
            O => \N__14231\,
            I => \N__14222\
        );

    \I__2549\ : IoSpan4Mux
    port map (
            O => \N__14228\,
            I => \N__14219\
        );

    \I__2548\ : Span4Mux_s2_h
    port map (
            O => \N__14225\,
            I => \N__14216\
        );

    \I__2547\ : Sp12to4
    port map (
            O => \N__14222\,
            I => \N__14213\
        );

    \I__2546\ : Span4Mux_s0_v
    port map (
            O => \N__14219\,
            I => \N__14210\
        );

    \I__2545\ : Sp12to4
    port map (
            O => \N__14216\,
            I => \N__14207\
        );

    \I__2544\ : Span12Mux_s9_h
    port map (
            O => \N__14213\,
            I => \N__14204\
        );

    \I__2543\ : Sp12to4
    port map (
            O => \N__14210\,
            I => \N__14201\
        );

    \I__2542\ : Span12Mux_v
    port map (
            O => \N__14207\,
            I => \N__14198\
        );

    \I__2541\ : Span12Mux_v
    port map (
            O => \N__14204\,
            I => \N__14193\
        );

    \I__2540\ : Span12Mux_v
    port map (
            O => \N__14201\,
            I => \N__14193\
        );

    \I__2539\ : Odrv12
    port map (
            O => \N__14198\,
            I => n1990
        );

    \I__2538\ : Odrv12
    port map (
            O => \N__14193\,
            I => n1990
        );

    \I__2537\ : InMux
    port map (
            O => \N__14188\,
            I => \N__14185\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__14185\,
            I => \TX_DATA_7\
        );

    \I__2535\ : IoInMux
    port map (
            O => \N__14182\,
            I => \N__14178\
        );

    \I__2534\ : IoInMux
    port map (
            O => \N__14181\,
            I => \N__14175\
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__14178\,
            I => \N__14172\
        );

    \I__2532\ : LocalMux
    port map (
            O => \N__14175\,
            I => \N__14168\
        );

    \I__2531\ : IoSpan4Mux
    port map (
            O => \N__14172\,
            I => \N__14165\
        );

    \I__2530\ : IoInMux
    port map (
            O => \N__14171\,
            I => \N__14162\
        );

    \I__2529\ : IoSpan4Mux
    port map (
            O => \N__14168\,
            I => \N__14159\
        );

    \I__2528\ : Span4Mux_s2_h
    port map (
            O => \N__14165\,
            I => \N__14156\
        );

    \I__2527\ : LocalMux
    port map (
            O => \N__14162\,
            I => \N__14153\
        );

    \I__2526\ : Span4Mux_s0_h
    port map (
            O => \N__14159\,
            I => \N__14150\
        );

    \I__2525\ : Sp12to4
    port map (
            O => \N__14156\,
            I => \N__14147\
        );

    \I__2524\ : IoSpan4Mux
    port map (
            O => \N__14153\,
            I => \N__14144\
        );

    \I__2523\ : Sp12to4
    port map (
            O => \N__14150\,
            I => \N__14141\
        );

    \I__2522\ : Span12Mux_s10_h
    port map (
            O => \N__14147\,
            I => \N__14138\
        );

    \I__2521\ : Sp12to4
    port map (
            O => \N__14144\,
            I => \N__14135\
        );

    \I__2520\ : Span12Mux_h
    port map (
            O => \N__14141\,
            I => \N__14132\
        );

    \I__2519\ : Span12Mux_v
    port map (
            O => \N__14138\,
            I => \N__14127\
        );

    \I__2518\ : Span12Mux_v
    port map (
            O => \N__14135\,
            I => \N__14127\
        );

    \I__2517\ : Odrv12
    port map (
            O => \N__14132\,
            I => \ADV_B_c\
        );

    \I__2516\ : Odrv12
    port map (
            O => \N__14127\,
            I => \ADV_B_c\
        );

    \I__2515\ : InMux
    port map (
            O => \N__14122\,
            I => \N__14118\
        );

    \I__2514\ : InMux
    port map (
            O => \N__14121\,
            I => \N__14115\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__14118\,
            I => \transmit_module.n186\
        );

    \I__2512\ : LocalMux
    port map (
            O => \N__14115\,
            I => \transmit_module.n186\
        );

    \I__2511\ : CascadeMux
    port map (
            O => \N__14110\,
            I => \transmit_module.n4211_cascade_\
        );

    \I__2510\ : InMux
    port map (
            O => \N__14107\,
            I => \N__14103\
        );

    \I__2509\ : InMux
    port map (
            O => \N__14106\,
            I => \N__14100\
        );

    \I__2508\ : LocalMux
    port map (
            O => \N__14103\,
            I => \transmit_module.n217\
        );

    \I__2507\ : LocalMux
    port map (
            O => \N__14100\,
            I => \transmit_module.n217\
        );

    \I__2506\ : CascadeMux
    port map (
            O => \N__14095\,
            I => \N__14091\
        );

    \I__2505\ : CascadeMux
    port map (
            O => \N__14094\,
            I => \N__14088\
        );

    \I__2504\ : CascadeBuf
    port map (
            O => \N__14091\,
            I => \N__14085\
        );

    \I__2503\ : CascadeBuf
    port map (
            O => \N__14088\,
            I => \N__14082\
        );

    \I__2502\ : CascadeMux
    port map (
            O => \N__14085\,
            I => \N__14079\
        );

    \I__2501\ : CascadeMux
    port map (
            O => \N__14082\,
            I => \N__14076\
        );

    \I__2500\ : CascadeBuf
    port map (
            O => \N__14079\,
            I => \N__14073\
        );

    \I__2499\ : CascadeBuf
    port map (
            O => \N__14076\,
            I => \N__14070\
        );

    \I__2498\ : CascadeMux
    port map (
            O => \N__14073\,
            I => \N__14067\
        );

    \I__2497\ : CascadeMux
    port map (
            O => \N__14070\,
            I => \N__14064\
        );

    \I__2496\ : CascadeBuf
    port map (
            O => \N__14067\,
            I => \N__14061\
        );

    \I__2495\ : CascadeBuf
    port map (
            O => \N__14064\,
            I => \N__14058\
        );

    \I__2494\ : CascadeMux
    port map (
            O => \N__14061\,
            I => \N__14055\
        );

    \I__2493\ : CascadeMux
    port map (
            O => \N__14058\,
            I => \N__14052\
        );

    \I__2492\ : CascadeBuf
    port map (
            O => \N__14055\,
            I => \N__14049\
        );

    \I__2491\ : CascadeBuf
    port map (
            O => \N__14052\,
            I => \N__14046\
        );

    \I__2490\ : CascadeMux
    port map (
            O => \N__14049\,
            I => \N__14043\
        );

    \I__2489\ : CascadeMux
    port map (
            O => \N__14046\,
            I => \N__14040\
        );

    \I__2488\ : CascadeBuf
    port map (
            O => \N__14043\,
            I => \N__14037\
        );

    \I__2487\ : CascadeBuf
    port map (
            O => \N__14040\,
            I => \N__14034\
        );

    \I__2486\ : CascadeMux
    port map (
            O => \N__14037\,
            I => \N__14031\
        );

    \I__2485\ : CascadeMux
    port map (
            O => \N__14034\,
            I => \N__14028\
        );

    \I__2484\ : CascadeBuf
    port map (
            O => \N__14031\,
            I => \N__14025\
        );

    \I__2483\ : CascadeBuf
    port map (
            O => \N__14028\,
            I => \N__14022\
        );

    \I__2482\ : CascadeMux
    port map (
            O => \N__14025\,
            I => \N__14019\
        );

    \I__2481\ : CascadeMux
    port map (
            O => \N__14022\,
            I => \N__14016\
        );

    \I__2480\ : CascadeBuf
    port map (
            O => \N__14019\,
            I => \N__14013\
        );

    \I__2479\ : CascadeBuf
    port map (
            O => \N__14016\,
            I => \N__14010\
        );

    \I__2478\ : CascadeMux
    port map (
            O => \N__14013\,
            I => \N__14007\
        );

    \I__2477\ : CascadeMux
    port map (
            O => \N__14010\,
            I => \N__14004\
        );

    \I__2476\ : CascadeBuf
    port map (
            O => \N__14007\,
            I => \N__14001\
        );

    \I__2475\ : CascadeBuf
    port map (
            O => \N__14004\,
            I => \N__13998\
        );

    \I__2474\ : CascadeMux
    port map (
            O => \N__14001\,
            I => \N__13995\
        );

    \I__2473\ : CascadeMux
    port map (
            O => \N__13998\,
            I => \N__13992\
        );

    \I__2472\ : CascadeBuf
    port map (
            O => \N__13995\,
            I => \N__13989\
        );

    \I__2471\ : CascadeBuf
    port map (
            O => \N__13992\,
            I => \N__13986\
        );

    \I__2470\ : CascadeMux
    port map (
            O => \N__13989\,
            I => \N__13983\
        );

    \I__2469\ : CascadeMux
    port map (
            O => \N__13986\,
            I => \N__13980\
        );

    \I__2468\ : CascadeBuf
    port map (
            O => \N__13983\,
            I => \N__13977\
        );

    \I__2467\ : CascadeBuf
    port map (
            O => \N__13980\,
            I => \N__13974\
        );

    \I__2466\ : CascadeMux
    port map (
            O => \N__13977\,
            I => \N__13971\
        );

    \I__2465\ : CascadeMux
    port map (
            O => \N__13974\,
            I => \N__13968\
        );

    \I__2464\ : CascadeBuf
    port map (
            O => \N__13971\,
            I => \N__13965\
        );

    \I__2463\ : CascadeBuf
    port map (
            O => \N__13968\,
            I => \N__13962\
        );

    \I__2462\ : CascadeMux
    port map (
            O => \N__13965\,
            I => \N__13959\
        );

    \I__2461\ : CascadeMux
    port map (
            O => \N__13962\,
            I => \N__13956\
        );

    \I__2460\ : CascadeBuf
    port map (
            O => \N__13959\,
            I => \N__13953\
        );

    \I__2459\ : CascadeBuf
    port map (
            O => \N__13956\,
            I => \N__13950\
        );

    \I__2458\ : CascadeMux
    port map (
            O => \N__13953\,
            I => \N__13947\
        );

    \I__2457\ : CascadeMux
    port map (
            O => \N__13950\,
            I => \N__13944\
        );

    \I__2456\ : CascadeBuf
    port map (
            O => \N__13947\,
            I => \N__13941\
        );

    \I__2455\ : CascadeBuf
    port map (
            O => \N__13944\,
            I => \N__13938\
        );

    \I__2454\ : CascadeMux
    port map (
            O => \N__13941\,
            I => \N__13935\
        );

    \I__2453\ : CascadeMux
    port map (
            O => \N__13938\,
            I => \N__13932\
        );

    \I__2452\ : CascadeBuf
    port map (
            O => \N__13935\,
            I => \N__13929\
        );

    \I__2451\ : CascadeBuf
    port map (
            O => \N__13932\,
            I => \N__13926\
        );

    \I__2450\ : CascadeMux
    port map (
            O => \N__13929\,
            I => \N__13923\
        );

    \I__2449\ : CascadeMux
    port map (
            O => \N__13926\,
            I => \N__13920\
        );

    \I__2448\ : CascadeBuf
    port map (
            O => \N__13923\,
            I => \N__13917\
        );

    \I__2447\ : CascadeBuf
    port map (
            O => \N__13920\,
            I => \N__13914\
        );

    \I__2446\ : CascadeMux
    port map (
            O => \N__13917\,
            I => \N__13911\
        );

    \I__2445\ : CascadeMux
    port map (
            O => \N__13914\,
            I => \N__13908\
        );

    \I__2444\ : InMux
    port map (
            O => \N__13911\,
            I => \N__13905\
        );

    \I__2443\ : InMux
    port map (
            O => \N__13908\,
            I => \N__13902\
        );

    \I__2442\ : LocalMux
    port map (
            O => \N__13905\,
            I => \N__13899\
        );

    \I__2441\ : LocalMux
    port map (
            O => \N__13902\,
            I => \N__13896\
        );

    \I__2440\ : Span4Mux_h
    port map (
            O => \N__13899\,
            I => \N__13893\
        );

    \I__2439\ : Span12Mux_s10_v
    port map (
            O => \N__13896\,
            I => \N__13890\
        );

    \I__2438\ : Span4Mux_h
    port map (
            O => \N__13893\,
            I => \N__13887\
        );

    \I__2437\ : Span12Mux_h
    port map (
            O => \N__13890\,
            I => \N__13884\
        );

    \I__2436\ : Sp12to4
    port map (
            O => \N__13887\,
            I => \N__13881\
        );

    \I__2435\ : Odrv12
    port map (
            O => \N__13884\,
            I => n26
        );

    \I__2434\ : Odrv12
    port map (
            O => \N__13881\,
            I => n26
        );

    \I__2433\ : InMux
    port map (
            O => \N__13876\,
            I => \N__13873\
        );

    \I__2432\ : LocalMux
    port map (
            O => \N__13873\,
            I => \N__13870\
        );

    \I__2431\ : Span12Mux_v
    port map (
            O => \N__13870\,
            I => \N__13867\
        );

    \I__2430\ : Span12Mux_h
    port map (
            O => \N__13867\,
            I => \N__13864\
        );

    \I__2429\ : Odrv12
    port map (
            O => \N__13864\,
            I => \line_buffer.n559\
        );

    \I__2428\ : InMux
    port map (
            O => \N__13861\,
            I => \N__13858\
        );

    \I__2427\ : LocalMux
    port map (
            O => \N__13858\,
            I => \N__13855\
        );

    \I__2426\ : Odrv4
    port map (
            O => \N__13855\,
            I => \line_buffer.n4182\
        );

    \I__2425\ : CascadeMux
    port map (
            O => \N__13852\,
            I => \N__13849\
        );

    \I__2424\ : InMux
    port map (
            O => \N__13849\,
            I => \N__13846\
        );

    \I__2423\ : LocalMux
    port map (
            O => \N__13846\,
            I => \N__13843\
        );

    \I__2422\ : Span12Mux_h
    port map (
            O => \N__13843\,
            I => \N__13840\
        );

    \I__2421\ : Odrv12
    port map (
            O => \N__13840\,
            I => \line_buffer.n551\
        );

    \I__2420\ : InMux
    port map (
            O => \N__13837\,
            I => \N__13827\
        );

    \I__2419\ : InMux
    port map (
            O => \N__13836\,
            I => \N__13827\
        );

    \I__2418\ : InMux
    port map (
            O => \N__13835\,
            I => \N__13827\
        );

    \I__2417\ : InMux
    port map (
            O => \N__13834\,
            I => \N__13824\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__13827\,
            I => \N__13821\
        );

    \I__2415\ : LocalMux
    port map (
            O => \N__13824\,
            I => \transmit_module.video_signal_controller.VGA_X_9\
        );

    \I__2414\ : Odrv4
    port map (
            O => \N__13821\,
            I => \transmit_module.video_signal_controller.VGA_X_9\
        );

    \I__2413\ : InMux
    port map (
            O => \N__13816\,
            I => \transmit_module.video_signal_controller.n3696\
        );

    \I__2412\ : CascadeMux
    port map (
            O => \N__13813\,
            I => \N__13808\
        );

    \I__2411\ : InMux
    port map (
            O => \N__13812\,
            I => \N__13804\
        );

    \I__2410\ : InMux
    port map (
            O => \N__13811\,
            I => \N__13797\
        );

    \I__2409\ : InMux
    port map (
            O => \N__13808\,
            I => \N__13797\
        );

    \I__2408\ : InMux
    port map (
            O => \N__13807\,
            I => \N__13797\
        );

    \I__2407\ : LocalMux
    port map (
            O => \N__13804\,
            I => \transmit_module.video_signal_controller.VGA_X_10\
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__13797\,
            I => \transmit_module.video_signal_controller.VGA_X_10\
        );

    \I__2405\ : InMux
    port map (
            O => \N__13792\,
            I => \transmit_module.video_signal_controller.n3697\
        );

    \I__2404\ : InMux
    port map (
            O => \N__13789\,
            I => \transmit_module.video_signal_controller.n3698\
        );

    \I__2403\ : InMux
    port map (
            O => \N__13786\,
            I => \N__13780\
        );

    \I__2402\ : InMux
    port map (
            O => \N__13785\,
            I => \N__13773\
        );

    \I__2401\ : InMux
    port map (
            O => \N__13784\,
            I => \N__13773\
        );

    \I__2400\ : InMux
    port map (
            O => \N__13783\,
            I => \N__13773\
        );

    \I__2399\ : LocalMux
    port map (
            O => \N__13780\,
            I => \transmit_module.video_signal_controller.VGA_X_11\
        );

    \I__2398\ : LocalMux
    port map (
            O => \N__13773\,
            I => \transmit_module.video_signal_controller.VGA_X_11\
        );

    \I__2397\ : CEMux
    port map (
            O => \N__13768\,
            I => \N__13765\
        );

    \I__2396\ : LocalMux
    port map (
            O => \N__13765\,
            I => \N__13762\
        );

    \I__2395\ : Span4Mux_v
    port map (
            O => \N__13762\,
            I => \N__13758\
        );

    \I__2394\ : CEMux
    port map (
            O => \N__13761\,
            I => \N__13755\
        );

    \I__2393\ : Span4Mux_h
    port map (
            O => \N__13758\,
            I => \N__13748\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__13755\,
            I => \N__13748\
        );

    \I__2391\ : SRMux
    port map (
            O => \N__13754\,
            I => \N__13745\
        );

    \I__2390\ : SRMux
    port map (
            O => \N__13753\,
            I => \N__13742\
        );

    \I__2389\ : Span4Mux_v
    port map (
            O => \N__13748\,
            I => \N__13739\
        );

    \I__2388\ : LocalMux
    port map (
            O => \N__13745\,
            I => \N__13736\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__13742\,
            I => \N__13733\
        );

    \I__2386\ : Odrv4
    port map (
            O => \N__13739\,
            I => \transmit_module.video_signal_controller.n2274\
        );

    \I__2385\ : Odrv4
    port map (
            O => \N__13736\,
            I => \transmit_module.video_signal_controller.n2274\
        );

    \I__2384\ : Odrv4
    port map (
            O => \N__13733\,
            I => \transmit_module.video_signal_controller.n2274\
        );

    \I__2383\ : InMux
    port map (
            O => \N__13726\,
            I => \N__13723\
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__13723\,
            I => \N__13720\
        );

    \I__2381\ : Odrv4
    port map (
            O => \N__13720\,
            I => \line_buffer.n4102\
        );

    \I__2380\ : InMux
    port map (
            O => \N__13717\,
            I => \N__13714\
        );

    \I__2379\ : LocalMux
    port map (
            O => \N__13714\,
            I => \N__13711\
        );

    \I__2378\ : Span12Mux_v
    port map (
            O => \N__13711\,
            I => \N__13708\
        );

    \I__2377\ : Span12Mux_h
    port map (
            O => \N__13708\,
            I => \N__13705\
        );

    \I__2376\ : Odrv12
    port map (
            O => \N__13705\,
            I => \line_buffer.n648\
        );

    \I__2375\ : CascadeMux
    port map (
            O => \N__13702\,
            I => \N__13699\
        );

    \I__2374\ : InMux
    port map (
            O => \N__13699\,
            I => \N__13696\
        );

    \I__2373\ : LocalMux
    port map (
            O => \N__13696\,
            I => \N__13693\
        );

    \I__2372\ : Span4Mux_v
    port map (
            O => \N__13693\,
            I => \N__13690\
        );

    \I__2371\ : Span4Mux_h
    port map (
            O => \N__13690\,
            I => \N__13687\
        );

    \I__2370\ : Odrv4
    port map (
            O => \N__13687\,
            I => \line_buffer.n656\
        );

    \I__2369\ : InMux
    port map (
            O => \N__13684\,
            I => \N__13678\
        );

    \I__2368\ : InMux
    port map (
            O => \N__13683\,
            I => \N__13673\
        );

    \I__2367\ : InMux
    port map (
            O => \N__13682\,
            I => \N__13673\
        );

    \I__2366\ : InMux
    port map (
            O => \N__13681\,
            I => \N__13670\
        );

    \I__2365\ : LocalMux
    port map (
            O => \N__13678\,
            I => \transmit_module.video_signal_controller.VGA_X_1\
        );

    \I__2364\ : LocalMux
    port map (
            O => \N__13673\,
            I => \transmit_module.video_signal_controller.VGA_X_1\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__13670\,
            I => \transmit_module.video_signal_controller.VGA_X_1\
        );

    \I__2362\ : InMux
    port map (
            O => \N__13663\,
            I => \transmit_module.video_signal_controller.n3688\
        );

    \I__2361\ : CascadeMux
    port map (
            O => \N__13660\,
            I => \N__13656\
        );

    \I__2360\ : InMux
    port map (
            O => \N__13659\,
            I => \N__13651\
        );

    \I__2359\ : InMux
    port map (
            O => \N__13656\,
            I => \N__13646\
        );

    \I__2358\ : InMux
    port map (
            O => \N__13655\,
            I => \N__13646\
        );

    \I__2357\ : InMux
    port map (
            O => \N__13654\,
            I => \N__13643\
        );

    \I__2356\ : LocalMux
    port map (
            O => \N__13651\,
            I => \transmit_module.video_signal_controller.VGA_X_2\
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__13646\,
            I => \transmit_module.video_signal_controller.VGA_X_2\
        );

    \I__2354\ : LocalMux
    port map (
            O => \N__13643\,
            I => \transmit_module.video_signal_controller.VGA_X_2\
        );

    \I__2353\ : InMux
    port map (
            O => \N__13636\,
            I => \transmit_module.video_signal_controller.n3689\
        );

    \I__2352\ : InMux
    port map (
            O => \N__13633\,
            I => \N__13627\
        );

    \I__2351\ : InMux
    port map (
            O => \N__13632\,
            I => \N__13624\
        );

    \I__2350\ : InMux
    port map (
            O => \N__13631\,
            I => \N__13621\
        );

    \I__2349\ : InMux
    port map (
            O => \N__13630\,
            I => \N__13618\
        );

    \I__2348\ : LocalMux
    port map (
            O => \N__13627\,
            I => \transmit_module.video_signal_controller.VGA_X_3\
        );

    \I__2347\ : LocalMux
    port map (
            O => \N__13624\,
            I => \transmit_module.video_signal_controller.VGA_X_3\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__13621\,
            I => \transmit_module.video_signal_controller.VGA_X_3\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__13618\,
            I => \transmit_module.video_signal_controller.VGA_X_3\
        );

    \I__2344\ : InMux
    port map (
            O => \N__13609\,
            I => \transmit_module.video_signal_controller.n3690\
        );

    \I__2343\ : InMux
    port map (
            O => \N__13606\,
            I => \N__13600\
        );

    \I__2342\ : InMux
    port map (
            O => \N__13605\,
            I => \N__13593\
        );

    \I__2341\ : InMux
    port map (
            O => \N__13604\,
            I => \N__13593\
        );

    \I__2340\ : InMux
    port map (
            O => \N__13603\,
            I => \N__13593\
        );

    \I__2339\ : LocalMux
    port map (
            O => \N__13600\,
            I => \transmit_module.video_signal_controller.VGA_X_4\
        );

    \I__2338\ : LocalMux
    port map (
            O => \N__13593\,
            I => \transmit_module.video_signal_controller.VGA_X_4\
        );

    \I__2337\ : InMux
    port map (
            O => \N__13588\,
            I => \transmit_module.video_signal_controller.n3691\
        );

    \I__2336\ : InMux
    port map (
            O => \N__13585\,
            I => \N__13579\
        );

    \I__2335\ : InMux
    port map (
            O => \N__13584\,
            I => \N__13574\
        );

    \I__2334\ : InMux
    port map (
            O => \N__13583\,
            I => \N__13574\
        );

    \I__2333\ : InMux
    port map (
            O => \N__13582\,
            I => \N__13571\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__13579\,
            I => \transmit_module.video_signal_controller.VGA_X_5\
        );

    \I__2331\ : LocalMux
    port map (
            O => \N__13574\,
            I => \transmit_module.video_signal_controller.VGA_X_5\
        );

    \I__2330\ : LocalMux
    port map (
            O => \N__13571\,
            I => \transmit_module.video_signal_controller.VGA_X_5\
        );

    \I__2329\ : InMux
    port map (
            O => \N__13564\,
            I => \transmit_module.video_signal_controller.n3692\
        );

    \I__2328\ : InMux
    port map (
            O => \N__13561\,
            I => \N__13555\
        );

    \I__2327\ : InMux
    port map (
            O => \N__13560\,
            I => \N__13550\
        );

    \I__2326\ : InMux
    port map (
            O => \N__13559\,
            I => \N__13550\
        );

    \I__2325\ : InMux
    port map (
            O => \N__13558\,
            I => \N__13547\
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__13555\,
            I => \transmit_module.video_signal_controller.VGA_X_6\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__13550\,
            I => \transmit_module.video_signal_controller.VGA_X_6\
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__13547\,
            I => \transmit_module.video_signal_controller.VGA_X_6\
        );

    \I__2321\ : InMux
    port map (
            O => \N__13540\,
            I => \transmit_module.video_signal_controller.n3693\
        );

    \I__2320\ : InMux
    port map (
            O => \N__13537\,
            I => \N__13529\
        );

    \I__2319\ : InMux
    port map (
            O => \N__13536\,
            I => \N__13529\
        );

    \I__2318\ : InMux
    port map (
            O => \N__13535\,
            I => \N__13526\
        );

    \I__2317\ : InMux
    port map (
            O => \N__13534\,
            I => \N__13523\
        );

    \I__2316\ : LocalMux
    port map (
            O => \N__13529\,
            I => \transmit_module.video_signal_controller.VGA_X_7\
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__13526\,
            I => \transmit_module.video_signal_controller.VGA_X_7\
        );

    \I__2314\ : LocalMux
    port map (
            O => \N__13523\,
            I => \transmit_module.video_signal_controller.VGA_X_7\
        );

    \I__2313\ : InMux
    port map (
            O => \N__13516\,
            I => \transmit_module.video_signal_controller.n3694\
        );

    \I__2312\ : InMux
    port map (
            O => \N__13513\,
            I => \N__13510\
        );

    \I__2311\ : LocalMux
    port map (
            O => \N__13510\,
            I => \N__13504\
        );

    \I__2310\ : InMux
    port map (
            O => \N__13509\,
            I => \N__13501\
        );

    \I__2309\ : InMux
    port map (
            O => \N__13508\,
            I => \N__13496\
        );

    \I__2308\ : InMux
    port map (
            O => \N__13507\,
            I => \N__13496\
        );

    \I__2307\ : Odrv4
    port map (
            O => \N__13504\,
            I => \transmit_module.video_signal_controller.VGA_X_8\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__13501\,
            I => \transmit_module.video_signal_controller.VGA_X_8\
        );

    \I__2305\ : LocalMux
    port map (
            O => \N__13496\,
            I => \transmit_module.video_signal_controller.VGA_X_8\
        );

    \I__2304\ : InMux
    port map (
            O => \N__13489\,
            I => \bfn_13_16_0_\
        );

    \I__2303\ : SRMux
    port map (
            O => \N__13486\,
            I => \N__13482\
        );

    \I__2302\ : SRMux
    port map (
            O => \N__13485\,
            I => \N__13479\
        );

    \I__2301\ : LocalMux
    port map (
            O => \N__13482\,
            I => \N__13476\
        );

    \I__2300\ : LocalMux
    port map (
            O => \N__13479\,
            I => \N__13471\
        );

    \I__2299\ : Span4Mux_v
    port map (
            O => \N__13476\,
            I => \N__13468\
        );

    \I__2298\ : SRMux
    port map (
            O => \N__13475\,
            I => \N__13465\
        );

    \I__2297\ : SRMux
    port map (
            O => \N__13474\,
            I => \N__13462\
        );

    \I__2296\ : Span12Mux_s2_v
    port map (
            O => \N__13471\,
            I => \N__13455\
        );

    \I__2295\ : Sp12to4
    port map (
            O => \N__13468\,
            I => \N__13455\
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__13465\,
            I => \N__13455\
        );

    \I__2293\ : LocalMux
    port map (
            O => \N__13462\,
            I => \N__13452\
        );

    \I__2292\ : Span12Mux_v
    port map (
            O => \N__13455\,
            I => \N__13449\
        );

    \I__2291\ : Span4Mux_v
    port map (
            O => \N__13452\,
            I => \N__13446\
        );

    \I__2290\ : Span12Mux_h
    port map (
            O => \N__13449\,
            I => \N__13443\
        );

    \I__2289\ : Span4Mux_h
    port map (
            O => \N__13446\,
            I => \N__13440\
        );

    \I__2288\ : Odrv12
    port map (
            O => \N__13443\,
            I => n690
        );

    \I__2287\ : Odrv4
    port map (
            O => \N__13440\,
            I => n690
        );

    \I__2286\ : CascadeMux
    port map (
            O => \N__13435\,
            I => \N__13432\
        );

    \I__2285\ : InMux
    port map (
            O => \N__13432\,
            I => \N__13429\
        );

    \I__2284\ : LocalMux
    port map (
            O => \N__13429\,
            I => \db5.COUNTER_3\
        );

    \I__2283\ : InMux
    port map (
            O => \N__13426\,
            I => \N__13419\
        );

    \I__2282\ : InMux
    port map (
            O => \N__13425\,
            I => \N__13419\
        );

    \I__2281\ : InMux
    port map (
            O => \N__13424\,
            I => \N__13416\
        );

    \I__2280\ : LocalMux
    port map (
            O => \N__13419\,
            I => \N__13413\
        );

    \I__2279\ : LocalMux
    port map (
            O => \N__13416\,
            I => \db5.NEXT_COUNTER_3\
        );

    \I__2278\ : Odrv4
    port map (
            O => \N__13413\,
            I => \db5.NEXT_COUNTER_3\
        );

    \I__2277\ : InMux
    port map (
            O => \N__13408\,
            I => \N__13404\
        );

    \I__2276\ : InMux
    port map (
            O => \N__13407\,
            I => \N__13401\
        );

    \I__2275\ : LocalMux
    port map (
            O => \N__13404\,
            I => \N__13396\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__13401\,
            I => \N__13396\
        );

    \I__2273\ : Odrv4
    port map (
            O => \N__13396\,
            I => \db5.COUNTER_2\
        );

    \I__2272\ : CascadeMux
    port map (
            O => \N__13393\,
            I => \N__13390\
        );

    \I__2271\ : InMux
    port map (
            O => \N__13390\,
            I => \N__13381\
        );

    \I__2270\ : InMux
    port map (
            O => \N__13389\,
            I => \N__13381\
        );

    \I__2269\ : InMux
    port map (
            O => \N__13388\,
            I => \N__13381\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__13381\,
            I => \N__13378\
        );

    \I__2267\ : Odrv4
    port map (
            O => \N__13378\,
            I => \db5.NEXT_COUNTER_2\
        );

    \I__2266\ : InMux
    port map (
            O => \N__13375\,
            I => \N__13366\
        );

    \I__2265\ : InMux
    port map (
            O => \N__13374\,
            I => \N__13366\
        );

    \I__2264\ : InMux
    port map (
            O => \N__13373\,
            I => \N__13366\
        );

    \I__2263\ : LocalMux
    port map (
            O => \N__13366\,
            I => \db5.COUNTER_1\
        );

    \I__2262\ : CascadeMux
    port map (
            O => \N__13363\,
            I => \N__13360\
        );

    \I__2261\ : InMux
    port map (
            O => \N__13360\,
            I => \N__13357\
        );

    \I__2260\ : LocalMux
    port map (
            O => \N__13357\,
            I => \N__13353\
        );

    \I__2259\ : InMux
    port map (
            O => \N__13356\,
            I => \N__13350\
        );

    \I__2258\ : Odrv4
    port map (
            O => \N__13353\,
            I => \db5.NEXT_COUNTER_1\
        );

    \I__2257\ : LocalMux
    port map (
            O => \N__13350\,
            I => \db5.NEXT_COUNTER_1\
        );

    \I__2256\ : InMux
    port map (
            O => \N__13345\,
            I => \N__13333\
        );

    \I__2255\ : InMux
    port map (
            O => \N__13344\,
            I => \N__13333\
        );

    \I__2254\ : InMux
    port map (
            O => \N__13343\,
            I => \N__13333\
        );

    \I__2253\ : InMux
    port map (
            O => \N__13342\,
            I => \N__13333\
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__13333\,
            I => \N__13330\
        );

    \I__2251\ : Odrv4
    port map (
            O => \N__13330\,
            I => \db5.COUNTER_0\
        );

    \I__2250\ : InMux
    port map (
            O => \N__13327\,
            I => \N__13321\
        );

    \I__2249\ : InMux
    port map (
            O => \N__13326\,
            I => \N__13321\
        );

    \I__2248\ : LocalMux
    port map (
            O => \N__13321\,
            I => \N__13318\
        );

    \I__2247\ : Odrv4
    port map (
            O => \N__13318\,
            I => \db5.NEXT_COUNTER_0\
        );

    \I__2246\ : SRMux
    port map (
            O => \N__13315\,
            I => \N__13312\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__13312\,
            I => \N__13309\
        );

    \I__2244\ : Span4Mux_v
    port map (
            O => \N__13309\,
            I => \N__13306\
        );

    \I__2243\ : Odrv4
    port map (
            O => \N__13306\,
            I => \db5.n4221\
        );

    \I__2242\ : CascadeMux
    port map (
            O => \N__13303\,
            I => \N__13300\
        );

    \I__2241\ : InMux
    port map (
            O => \N__13300\,
            I => \N__13297\
        );

    \I__2240\ : LocalMux
    port map (
            O => \N__13297\,
            I => \transmit_module.video_signal_controller.n3997\
        );

    \I__2239\ : InMux
    port map (
            O => \N__13294\,
            I => \N__13291\
        );

    \I__2238\ : LocalMux
    port map (
            O => \N__13291\,
            I => \transmit_module.video_signal_controller.n3196\
        );

    \I__2237\ : InMux
    port map (
            O => \N__13288\,
            I => \N__13285\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__13285\,
            I => \N__13282\
        );

    \I__2235\ : Span4Mux_v
    port map (
            O => \N__13282\,
            I => \N__13279\
        );

    \I__2234\ : Span4Mux_v
    port map (
            O => \N__13279\,
            I => \N__13276\
        );

    \I__2233\ : Span4Mux_h
    port map (
            O => \N__13276\,
            I => \N__13273\
        );

    \I__2232\ : Odrv4
    port map (
            O => \N__13273\,
            I => \line_buffer.n655\
        );

    \I__2231\ : InMux
    port map (
            O => \N__13270\,
            I => \N__13267\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__13267\,
            I => \N__13264\
        );

    \I__2229\ : Span12Mux_v
    port map (
            O => \N__13264\,
            I => \N__13261\
        );

    \I__2228\ : Span12Mux_h
    port map (
            O => \N__13261\,
            I => \N__13258\
        );

    \I__2227\ : Odrv12
    port map (
            O => \N__13258\,
            I => \line_buffer.n647\
        );

    \I__2226\ : InMux
    port map (
            O => \N__13255\,
            I => \N__13250\
        );

    \I__2225\ : InMux
    port map (
            O => \N__13254\,
            I => \N__13245\
        );

    \I__2224\ : InMux
    port map (
            O => \N__13253\,
            I => \N__13245\
        );

    \I__2223\ : LocalMux
    port map (
            O => \N__13250\,
            I => \transmit_module.video_signal_controller.VGA_X_0\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__13245\,
            I => \transmit_module.video_signal_controller.VGA_X_0\
        );

    \I__2221\ : InMux
    port map (
            O => \N__13240\,
            I => \bfn_13_15_0_\
        );

    \I__2220\ : InMux
    port map (
            O => \N__13237\,
            I => \N__13234\
        );

    \I__2219\ : LocalMux
    port map (
            O => \N__13234\,
            I => \receive_module.n7\
        );

    \I__2218\ : CascadeMux
    port map (
            O => \N__13231\,
            I => \N__13228\
        );

    \I__2217\ : InMux
    port map (
            O => \N__13228\,
            I => \N__13225\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__13225\,
            I => \N__13222\
        );

    \I__2215\ : Span4Mux_v
    port map (
            O => \N__13222\,
            I => \N__13217\
        );

    \I__2214\ : InMux
    port map (
            O => \N__13221\,
            I => \N__13212\
        );

    \I__2213\ : InMux
    port map (
            O => \N__13220\,
            I => \N__13212\
        );

    \I__2212\ : Odrv4
    port map (
            O => \N__13217\,
            I => \receive_module.O_Y_3\
        );

    \I__2211\ : LocalMux
    port map (
            O => \N__13212\,
            I => \receive_module.O_Y_3\
        );

    \I__2210\ : CascadeMux
    port map (
            O => \N__13207\,
            I => \N__13203\
        );

    \I__2209\ : CascadeMux
    port map (
            O => \N__13206\,
            I => \N__13200\
        );

    \I__2208\ : CascadeBuf
    port map (
            O => \N__13203\,
            I => \N__13197\
        );

    \I__2207\ : CascadeBuf
    port map (
            O => \N__13200\,
            I => \N__13194\
        );

    \I__2206\ : CascadeMux
    port map (
            O => \N__13197\,
            I => \N__13191\
        );

    \I__2205\ : CascadeMux
    port map (
            O => \N__13194\,
            I => \N__13188\
        );

    \I__2204\ : CascadeBuf
    port map (
            O => \N__13191\,
            I => \N__13185\
        );

    \I__2203\ : CascadeBuf
    port map (
            O => \N__13188\,
            I => \N__13182\
        );

    \I__2202\ : CascadeMux
    port map (
            O => \N__13185\,
            I => \N__13179\
        );

    \I__2201\ : CascadeMux
    port map (
            O => \N__13182\,
            I => \N__13176\
        );

    \I__2200\ : CascadeBuf
    port map (
            O => \N__13179\,
            I => \N__13173\
        );

    \I__2199\ : CascadeBuf
    port map (
            O => \N__13176\,
            I => \N__13170\
        );

    \I__2198\ : CascadeMux
    port map (
            O => \N__13173\,
            I => \N__13167\
        );

    \I__2197\ : CascadeMux
    port map (
            O => \N__13170\,
            I => \N__13164\
        );

    \I__2196\ : CascadeBuf
    port map (
            O => \N__13167\,
            I => \N__13161\
        );

    \I__2195\ : CascadeBuf
    port map (
            O => \N__13164\,
            I => \N__13158\
        );

    \I__2194\ : CascadeMux
    port map (
            O => \N__13161\,
            I => \N__13155\
        );

    \I__2193\ : CascadeMux
    port map (
            O => \N__13158\,
            I => \N__13152\
        );

    \I__2192\ : CascadeBuf
    port map (
            O => \N__13155\,
            I => \N__13149\
        );

    \I__2191\ : CascadeBuf
    port map (
            O => \N__13152\,
            I => \N__13146\
        );

    \I__2190\ : CascadeMux
    port map (
            O => \N__13149\,
            I => \N__13143\
        );

    \I__2189\ : CascadeMux
    port map (
            O => \N__13146\,
            I => \N__13140\
        );

    \I__2188\ : CascadeBuf
    port map (
            O => \N__13143\,
            I => \N__13137\
        );

    \I__2187\ : CascadeBuf
    port map (
            O => \N__13140\,
            I => \N__13134\
        );

    \I__2186\ : CascadeMux
    port map (
            O => \N__13137\,
            I => \N__13131\
        );

    \I__2185\ : CascadeMux
    port map (
            O => \N__13134\,
            I => \N__13128\
        );

    \I__2184\ : CascadeBuf
    port map (
            O => \N__13131\,
            I => \N__13125\
        );

    \I__2183\ : CascadeBuf
    port map (
            O => \N__13128\,
            I => \N__13122\
        );

    \I__2182\ : CascadeMux
    port map (
            O => \N__13125\,
            I => \N__13119\
        );

    \I__2181\ : CascadeMux
    port map (
            O => \N__13122\,
            I => \N__13116\
        );

    \I__2180\ : CascadeBuf
    port map (
            O => \N__13119\,
            I => \N__13113\
        );

    \I__2179\ : CascadeBuf
    port map (
            O => \N__13116\,
            I => \N__13110\
        );

    \I__2178\ : CascadeMux
    port map (
            O => \N__13113\,
            I => \N__13107\
        );

    \I__2177\ : CascadeMux
    port map (
            O => \N__13110\,
            I => \N__13104\
        );

    \I__2176\ : CascadeBuf
    port map (
            O => \N__13107\,
            I => \N__13101\
        );

    \I__2175\ : CascadeBuf
    port map (
            O => \N__13104\,
            I => \N__13098\
        );

    \I__2174\ : CascadeMux
    port map (
            O => \N__13101\,
            I => \N__13095\
        );

    \I__2173\ : CascadeMux
    port map (
            O => \N__13098\,
            I => \N__13092\
        );

    \I__2172\ : CascadeBuf
    port map (
            O => \N__13095\,
            I => \N__13089\
        );

    \I__2171\ : CascadeBuf
    port map (
            O => \N__13092\,
            I => \N__13086\
        );

    \I__2170\ : CascadeMux
    port map (
            O => \N__13089\,
            I => \N__13083\
        );

    \I__2169\ : CascadeMux
    port map (
            O => \N__13086\,
            I => \N__13080\
        );

    \I__2168\ : CascadeBuf
    port map (
            O => \N__13083\,
            I => \N__13077\
        );

    \I__2167\ : CascadeBuf
    port map (
            O => \N__13080\,
            I => \N__13074\
        );

    \I__2166\ : CascadeMux
    port map (
            O => \N__13077\,
            I => \N__13071\
        );

    \I__2165\ : CascadeMux
    port map (
            O => \N__13074\,
            I => \N__13068\
        );

    \I__2164\ : CascadeBuf
    port map (
            O => \N__13071\,
            I => \N__13065\
        );

    \I__2163\ : CascadeBuf
    port map (
            O => \N__13068\,
            I => \N__13062\
        );

    \I__2162\ : CascadeMux
    port map (
            O => \N__13065\,
            I => \N__13059\
        );

    \I__2161\ : CascadeMux
    port map (
            O => \N__13062\,
            I => \N__13056\
        );

    \I__2160\ : CascadeBuf
    port map (
            O => \N__13059\,
            I => \N__13053\
        );

    \I__2159\ : CascadeBuf
    port map (
            O => \N__13056\,
            I => \N__13050\
        );

    \I__2158\ : CascadeMux
    port map (
            O => \N__13053\,
            I => \N__13047\
        );

    \I__2157\ : CascadeMux
    port map (
            O => \N__13050\,
            I => \N__13044\
        );

    \I__2156\ : CascadeBuf
    port map (
            O => \N__13047\,
            I => \N__13041\
        );

    \I__2155\ : CascadeBuf
    port map (
            O => \N__13044\,
            I => \N__13038\
        );

    \I__2154\ : CascadeMux
    port map (
            O => \N__13041\,
            I => \N__13035\
        );

    \I__2153\ : CascadeMux
    port map (
            O => \N__13038\,
            I => \N__13032\
        );

    \I__2152\ : CascadeBuf
    port map (
            O => \N__13035\,
            I => \N__13029\
        );

    \I__2151\ : CascadeBuf
    port map (
            O => \N__13032\,
            I => \N__13026\
        );

    \I__2150\ : CascadeMux
    port map (
            O => \N__13029\,
            I => \N__13023\
        );

    \I__2149\ : CascadeMux
    port map (
            O => \N__13026\,
            I => \N__13020\
        );

    \I__2148\ : InMux
    port map (
            O => \N__13023\,
            I => \N__13017\
        );

    \I__2147\ : InMux
    port map (
            O => \N__13020\,
            I => \N__13014\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__13017\,
            I => \N__13011\
        );

    \I__2145\ : LocalMux
    port map (
            O => \N__13014\,
            I => \N__13008\
        );

    \I__2144\ : Span4Mux_h
    port map (
            O => \N__13011\,
            I => \N__13005\
        );

    \I__2143\ : Span12Mux_s6_v
    port map (
            O => \N__13008\,
            I => \N__13002\
        );

    \I__2142\ : Sp12to4
    port map (
            O => \N__13005\,
            I => \N__12999\
        );

    \I__2141\ : Span12Mux_v
    port map (
            O => \N__13002\,
            I => \N__12996\
        );

    \I__2140\ : Span12Mux_s9_v
    port map (
            O => \N__12999\,
            I => \N__12993\
        );

    \I__2139\ : Span12Mux_h
    port map (
            O => \N__12996\,
            I => \N__12990\
        );

    \I__2138\ : Span12Mux_v
    port map (
            O => \N__12993\,
            I => \N__12987\
        );

    \I__2137\ : Odrv12
    port map (
            O => \N__12990\,
            I => \RX_ADDR_9\
        );

    \I__2136\ : Odrv12
    port map (
            O => \N__12987\,
            I => \RX_ADDR_9\
        );

    \I__2135\ : InMux
    port map (
            O => \N__12982\,
            I => \receive_module.n3701\
        );

    \I__2134\ : InMux
    port map (
            O => \N__12979\,
            I => \N__12976\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__12976\,
            I => \receive_module.n6\
        );

    \I__2132\ : CascadeMux
    port map (
            O => \N__12973\,
            I => \N__12970\
        );

    \I__2131\ : InMux
    port map (
            O => \N__12970\,
            I => \N__12967\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__12967\,
            I => \N__12964\
        );

    \I__2129\ : Span4Mux_h
    port map (
            O => \N__12964\,
            I => \N__12960\
        );

    \I__2128\ : InMux
    port map (
            O => \N__12963\,
            I => \N__12957\
        );

    \I__2127\ : Odrv4
    port map (
            O => \N__12960\,
            I => \receive_module.O_Y_4\
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__12957\,
            I => \receive_module.O_Y_4\
        );

    \I__2125\ : CascadeMux
    port map (
            O => \N__12952\,
            I => \N__12949\
        );

    \I__2124\ : CascadeBuf
    port map (
            O => \N__12949\,
            I => \N__12945\
        );

    \I__2123\ : CascadeMux
    port map (
            O => \N__12948\,
            I => \N__12942\
        );

    \I__2122\ : CascadeMux
    port map (
            O => \N__12945\,
            I => \N__12939\
        );

    \I__2121\ : CascadeBuf
    port map (
            O => \N__12942\,
            I => \N__12936\
        );

    \I__2120\ : CascadeBuf
    port map (
            O => \N__12939\,
            I => \N__12933\
        );

    \I__2119\ : CascadeMux
    port map (
            O => \N__12936\,
            I => \N__12930\
        );

    \I__2118\ : CascadeMux
    port map (
            O => \N__12933\,
            I => \N__12927\
        );

    \I__2117\ : CascadeBuf
    port map (
            O => \N__12930\,
            I => \N__12924\
        );

    \I__2116\ : CascadeBuf
    port map (
            O => \N__12927\,
            I => \N__12921\
        );

    \I__2115\ : CascadeMux
    port map (
            O => \N__12924\,
            I => \N__12918\
        );

    \I__2114\ : CascadeMux
    port map (
            O => \N__12921\,
            I => \N__12915\
        );

    \I__2113\ : CascadeBuf
    port map (
            O => \N__12918\,
            I => \N__12912\
        );

    \I__2112\ : CascadeBuf
    port map (
            O => \N__12915\,
            I => \N__12909\
        );

    \I__2111\ : CascadeMux
    port map (
            O => \N__12912\,
            I => \N__12906\
        );

    \I__2110\ : CascadeMux
    port map (
            O => \N__12909\,
            I => \N__12903\
        );

    \I__2109\ : CascadeBuf
    port map (
            O => \N__12906\,
            I => \N__12900\
        );

    \I__2108\ : CascadeBuf
    port map (
            O => \N__12903\,
            I => \N__12897\
        );

    \I__2107\ : CascadeMux
    port map (
            O => \N__12900\,
            I => \N__12894\
        );

    \I__2106\ : CascadeMux
    port map (
            O => \N__12897\,
            I => \N__12891\
        );

    \I__2105\ : CascadeBuf
    port map (
            O => \N__12894\,
            I => \N__12888\
        );

    \I__2104\ : CascadeBuf
    port map (
            O => \N__12891\,
            I => \N__12885\
        );

    \I__2103\ : CascadeMux
    port map (
            O => \N__12888\,
            I => \N__12882\
        );

    \I__2102\ : CascadeMux
    port map (
            O => \N__12885\,
            I => \N__12879\
        );

    \I__2101\ : CascadeBuf
    port map (
            O => \N__12882\,
            I => \N__12876\
        );

    \I__2100\ : CascadeBuf
    port map (
            O => \N__12879\,
            I => \N__12873\
        );

    \I__2099\ : CascadeMux
    port map (
            O => \N__12876\,
            I => \N__12870\
        );

    \I__2098\ : CascadeMux
    port map (
            O => \N__12873\,
            I => \N__12867\
        );

    \I__2097\ : CascadeBuf
    port map (
            O => \N__12870\,
            I => \N__12864\
        );

    \I__2096\ : CascadeBuf
    port map (
            O => \N__12867\,
            I => \N__12861\
        );

    \I__2095\ : CascadeMux
    port map (
            O => \N__12864\,
            I => \N__12858\
        );

    \I__2094\ : CascadeMux
    port map (
            O => \N__12861\,
            I => \N__12855\
        );

    \I__2093\ : CascadeBuf
    port map (
            O => \N__12858\,
            I => \N__12852\
        );

    \I__2092\ : CascadeBuf
    port map (
            O => \N__12855\,
            I => \N__12849\
        );

    \I__2091\ : CascadeMux
    port map (
            O => \N__12852\,
            I => \N__12846\
        );

    \I__2090\ : CascadeMux
    port map (
            O => \N__12849\,
            I => \N__12843\
        );

    \I__2089\ : CascadeBuf
    port map (
            O => \N__12846\,
            I => \N__12840\
        );

    \I__2088\ : CascadeBuf
    port map (
            O => \N__12843\,
            I => \N__12837\
        );

    \I__2087\ : CascadeMux
    port map (
            O => \N__12840\,
            I => \N__12834\
        );

    \I__2086\ : CascadeMux
    port map (
            O => \N__12837\,
            I => \N__12831\
        );

    \I__2085\ : CascadeBuf
    port map (
            O => \N__12834\,
            I => \N__12828\
        );

    \I__2084\ : CascadeBuf
    port map (
            O => \N__12831\,
            I => \N__12825\
        );

    \I__2083\ : CascadeMux
    port map (
            O => \N__12828\,
            I => \N__12822\
        );

    \I__2082\ : CascadeMux
    port map (
            O => \N__12825\,
            I => \N__12819\
        );

    \I__2081\ : CascadeBuf
    port map (
            O => \N__12822\,
            I => \N__12816\
        );

    \I__2080\ : CascadeBuf
    port map (
            O => \N__12819\,
            I => \N__12813\
        );

    \I__2079\ : CascadeMux
    port map (
            O => \N__12816\,
            I => \N__12810\
        );

    \I__2078\ : CascadeMux
    port map (
            O => \N__12813\,
            I => \N__12807\
        );

    \I__2077\ : CascadeBuf
    port map (
            O => \N__12810\,
            I => \N__12804\
        );

    \I__2076\ : CascadeBuf
    port map (
            O => \N__12807\,
            I => \N__12801\
        );

    \I__2075\ : CascadeMux
    port map (
            O => \N__12804\,
            I => \N__12798\
        );

    \I__2074\ : CascadeMux
    port map (
            O => \N__12801\,
            I => \N__12795\
        );

    \I__2073\ : CascadeBuf
    port map (
            O => \N__12798\,
            I => \N__12792\
        );

    \I__2072\ : CascadeBuf
    port map (
            O => \N__12795\,
            I => \N__12789\
        );

    \I__2071\ : CascadeMux
    port map (
            O => \N__12792\,
            I => \N__12786\
        );

    \I__2070\ : CascadeMux
    port map (
            O => \N__12789\,
            I => \N__12783\
        );

    \I__2069\ : CascadeBuf
    port map (
            O => \N__12786\,
            I => \N__12780\
        );

    \I__2068\ : CascadeBuf
    port map (
            O => \N__12783\,
            I => \N__12777\
        );

    \I__2067\ : CascadeMux
    port map (
            O => \N__12780\,
            I => \N__12774\
        );

    \I__2066\ : CascadeMux
    port map (
            O => \N__12777\,
            I => \N__12771\
        );

    \I__2065\ : CascadeBuf
    port map (
            O => \N__12774\,
            I => \N__12768\
        );

    \I__2064\ : InMux
    port map (
            O => \N__12771\,
            I => \N__12765\
        );

    \I__2063\ : CascadeMux
    port map (
            O => \N__12768\,
            I => \N__12762\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__12765\,
            I => \N__12759\
        );

    \I__2061\ : InMux
    port map (
            O => \N__12762\,
            I => \N__12756\
        );

    \I__2060\ : Span4Mux_s1_v
    port map (
            O => \N__12759\,
            I => \N__12753\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__12756\,
            I => \N__12750\
        );

    \I__2058\ : Span4Mux_h
    port map (
            O => \N__12753\,
            I => \N__12747\
        );

    \I__2057\ : Span12Mux_s5_v
    port map (
            O => \N__12750\,
            I => \N__12744\
        );

    \I__2056\ : Span4Mux_v
    port map (
            O => \N__12747\,
            I => \N__12741\
        );

    \I__2055\ : Span12Mux_h
    port map (
            O => \N__12744\,
            I => \N__12736\
        );

    \I__2054\ : Sp12to4
    port map (
            O => \N__12741\,
            I => \N__12736\
        );

    \I__2053\ : Span12Mux_v
    port map (
            O => \N__12736\,
            I => \N__12733\
        );

    \I__2052\ : Odrv12
    port map (
            O => \N__12733\,
            I => \RX_ADDR_10\
        );

    \I__2051\ : InMux
    port map (
            O => \N__12730\,
            I => \receive_module.n3702\
        );

    \I__2050\ : InMux
    port map (
            O => \N__12727\,
            I => \N__12724\
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__12724\,
            I => \receive_module.n5\
        );

    \I__2048\ : CascadeMux
    port map (
            O => \N__12721\,
            I => \N__12718\
        );

    \I__2047\ : InMux
    port map (
            O => \N__12718\,
            I => \N__12715\
        );

    \I__2046\ : LocalMux
    port map (
            O => \N__12715\,
            I => \N__12712\
        );

    \I__2045\ : Span4Mux_h
    port map (
            O => \N__12712\,
            I => \N__12709\
        );

    \I__2044\ : Odrv4
    port map (
            O => \N__12709\,
            I => \receive_module.O_Y_5\
        );

    \I__2043\ : InMux
    port map (
            O => \N__12706\,
            I => \receive_module.n3703\
        );

    \I__2042\ : InMux
    port map (
            O => \N__12703\,
            I => \N__12700\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__12700\,
            I => \receive_module.n4\
        );

    \I__2040\ : CascadeMux
    port map (
            O => \N__12697\,
            I => \N__12694\
        );

    \I__2039\ : InMux
    port map (
            O => \N__12694\,
            I => \N__12691\
        );

    \I__2038\ : LocalMux
    port map (
            O => \N__12691\,
            I => \N__12688\
        );

    \I__2037\ : Span4Mux_h
    port map (
            O => \N__12688\,
            I => \N__12685\
        );

    \I__2036\ : Odrv4
    port map (
            O => \N__12685\,
            I => \receive_module.O_Y_6\
        );

    \I__2035\ : InMux
    port map (
            O => \N__12682\,
            I => \receive_module.n3704\
        );

    \I__2034\ : InMux
    port map (
            O => \N__12679\,
            I => \N__12676\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__12676\,
            I => \receive_module.n3\
        );

    \I__2032\ : InMux
    port map (
            O => \N__12673\,
            I => \N__12670\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__12670\,
            I => \N__12667\
        );

    \I__2030\ : Span4Mux_v
    port map (
            O => \N__12667\,
            I => \N__12664\
        );

    \I__2029\ : Odrv4
    port map (
            O => \N__12664\,
            I => \receive_module.O_Y_7\
        );

    \I__2028\ : InMux
    port map (
            O => \N__12661\,
            I => \receive_module.n3705\
        );

    \I__2027\ : SRMux
    port map (
            O => \N__12658\,
            I => \N__12653\
        );

    \I__2026\ : SRMux
    port map (
            O => \N__12657\,
            I => \N__12650\
        );

    \I__2025\ : SRMux
    port map (
            O => \N__12656\,
            I => \N__12647\
        );

    \I__2024\ : LocalMux
    port map (
            O => \N__12653\,
            I => \N__12643\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__12650\,
            I => \N__12638\
        );

    \I__2022\ : LocalMux
    port map (
            O => \N__12647\,
            I => \N__12638\
        );

    \I__2021\ : SRMux
    port map (
            O => \N__12646\,
            I => \N__12635\
        );

    \I__2020\ : Span4Mux_v
    port map (
            O => \N__12643\,
            I => \N__12632\
        );

    \I__2019\ : Span4Mux_s3_v
    port map (
            O => \N__12638\,
            I => \N__12627\
        );

    \I__2018\ : LocalMux
    port map (
            O => \N__12635\,
            I => \N__12627\
        );

    \I__2017\ : Span4Mux_h
    port map (
            O => \N__12632\,
            I => \N__12624\
        );

    \I__2016\ : Span4Mux_v
    port map (
            O => \N__12627\,
            I => \N__12621\
        );

    \I__2015\ : Span4Mux_v
    port map (
            O => \N__12624\,
            I => \N__12618\
        );

    \I__2014\ : Span4Mux_h
    port map (
            O => \N__12621\,
            I => \N__12615\
        );

    \I__2013\ : Odrv4
    port map (
            O => \N__12618\,
            I => \line_buffer.n627\
        );

    \I__2012\ : Odrv4
    port map (
            O => \N__12615\,
            I => \line_buffer.n627\
        );

    \I__2011\ : SRMux
    port map (
            O => \N__12610\,
            I => \N__12607\
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__12607\,
            I => \N__12602\
        );

    \I__2009\ : SRMux
    port map (
            O => \N__12606\,
            I => \N__12599\
        );

    \I__2008\ : SRMux
    port map (
            O => \N__12605\,
            I => \N__12595\
        );

    \I__2007\ : Span4Mux_h
    port map (
            O => \N__12602\,
            I => \N__12592\
        );

    \I__2006\ : LocalMux
    port map (
            O => \N__12599\,
            I => \N__12589\
        );

    \I__2005\ : SRMux
    port map (
            O => \N__12598\,
            I => \N__12586\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__12595\,
            I => \N__12583\
        );

    \I__2003\ : Span4Mux_v
    port map (
            O => \N__12592\,
            I => \N__12578\
        );

    \I__2002\ : Span4Mux_h
    port map (
            O => \N__12589\,
            I => \N__12578\
        );

    \I__2001\ : LocalMux
    port map (
            O => \N__12586\,
            I => \N__12575\
        );

    \I__2000\ : Span12Mux_s10_v
    port map (
            O => \N__12583\,
            I => \N__12570\
        );

    \I__1999\ : Sp12to4
    port map (
            O => \N__12578\,
            I => \N__12570\
        );

    \I__1998\ : Span12Mux_v
    port map (
            O => \N__12575\,
            I => \N__12567\
        );

    \I__1997\ : Span12Mux_h
    port map (
            O => \N__12570\,
            I => \N__12562\
        );

    \I__1996\ : Span12Mux_h
    port map (
            O => \N__12567\,
            I => \N__12562\
        );

    \I__1995\ : Odrv12
    port map (
            O => \N__12562\,
            I => \line_buffer.n562\
        );

    \I__1994\ : InMux
    port map (
            O => \N__12559\,
            I => \receive_module.rx_counter.n3652\
        );

    \I__1993\ : InMux
    port map (
            O => \N__12556\,
            I => \receive_module.rx_counter.n3653\
        );

    \I__1992\ : InMux
    port map (
            O => \N__12553\,
            I => \receive_module.rx_counter.n3654\
        );

    \I__1991\ : InMux
    port map (
            O => \N__12550\,
            I => \receive_module.rx_counter.n3655\
        );

    \I__1990\ : InMux
    port map (
            O => \N__12547\,
            I => \N__12532\
        );

    \I__1989\ : InMux
    port map (
            O => \N__12546\,
            I => \N__12532\
        );

    \I__1988\ : InMux
    port map (
            O => \N__12545\,
            I => \N__12532\
        );

    \I__1987\ : InMux
    port map (
            O => \N__12544\,
            I => \N__12532\
        );

    \I__1986\ : InMux
    port map (
            O => \N__12543\,
            I => \N__12532\
        );

    \I__1985\ : LocalMux
    port map (
            O => \N__12532\,
            I => \receive_module.O_X_9\
        );

    \I__1984\ : CascadeMux
    port map (
            O => \N__12529\,
            I => \N__12526\
        );

    \I__1983\ : InMux
    port map (
            O => \N__12526\,
            I => \N__12523\
        );

    \I__1982\ : LocalMux
    port map (
            O => \N__12523\,
            I => \receive_module.rx_counter.n4\
        );

    \I__1981\ : InMux
    port map (
            O => \N__12520\,
            I => \N__12517\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__12517\,
            I => \N__12513\
        );

    \I__1979\ : CascadeMux
    port map (
            O => \N__12516\,
            I => \N__12509\
        );

    \I__1978\ : Span4Mux_h
    port map (
            O => \N__12513\,
            I => \N__12503\
        );

    \I__1977\ : InMux
    port map (
            O => \N__12512\,
            I => \N__12500\
        );

    \I__1976\ : InMux
    port map (
            O => \N__12509\,
            I => \N__12491\
        );

    \I__1975\ : InMux
    port map (
            O => \N__12508\,
            I => \N__12491\
        );

    \I__1974\ : InMux
    port map (
            O => \N__12507\,
            I => \N__12491\
        );

    \I__1973\ : InMux
    port map (
            O => \N__12506\,
            I => \N__12491\
        );

    \I__1972\ : Odrv4
    port map (
            O => \N__12503\,
            I => \receive_module.O_Y_0\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__12500\,
            I => \receive_module.O_Y_0\
        );

    \I__1970\ : LocalMux
    port map (
            O => \N__12491\,
            I => \receive_module.O_Y_0\
        );

    \I__1969\ : CascadeMux
    port map (
            O => \N__12484\,
            I => \N__12481\
        );

    \I__1968\ : InMux
    port map (
            O => \N__12481\,
            I => \N__12478\
        );

    \I__1967\ : LocalMux
    port map (
            O => \N__12478\,
            I => \receive_module.O_X_6\
        );

    \I__1966\ : CascadeMux
    port map (
            O => \N__12475\,
            I => \N__12472\
        );

    \I__1965\ : CascadeBuf
    port map (
            O => \N__12472\,
            I => \N__12469\
        );

    \I__1964\ : CascadeMux
    port map (
            O => \N__12469\,
            I => \N__12465\
        );

    \I__1963\ : CascadeMux
    port map (
            O => \N__12468\,
            I => \N__12462\
        );

    \I__1962\ : CascadeBuf
    port map (
            O => \N__12465\,
            I => \N__12459\
        );

    \I__1961\ : CascadeBuf
    port map (
            O => \N__12462\,
            I => \N__12456\
        );

    \I__1960\ : CascadeMux
    port map (
            O => \N__12459\,
            I => \N__12453\
        );

    \I__1959\ : CascadeMux
    port map (
            O => \N__12456\,
            I => \N__12450\
        );

    \I__1958\ : CascadeBuf
    port map (
            O => \N__12453\,
            I => \N__12447\
        );

    \I__1957\ : CascadeBuf
    port map (
            O => \N__12450\,
            I => \N__12444\
        );

    \I__1956\ : CascadeMux
    port map (
            O => \N__12447\,
            I => \N__12441\
        );

    \I__1955\ : CascadeMux
    port map (
            O => \N__12444\,
            I => \N__12438\
        );

    \I__1954\ : CascadeBuf
    port map (
            O => \N__12441\,
            I => \N__12435\
        );

    \I__1953\ : CascadeBuf
    port map (
            O => \N__12438\,
            I => \N__12432\
        );

    \I__1952\ : CascadeMux
    port map (
            O => \N__12435\,
            I => \N__12429\
        );

    \I__1951\ : CascadeMux
    port map (
            O => \N__12432\,
            I => \N__12426\
        );

    \I__1950\ : CascadeBuf
    port map (
            O => \N__12429\,
            I => \N__12423\
        );

    \I__1949\ : CascadeBuf
    port map (
            O => \N__12426\,
            I => \N__12420\
        );

    \I__1948\ : CascadeMux
    port map (
            O => \N__12423\,
            I => \N__12417\
        );

    \I__1947\ : CascadeMux
    port map (
            O => \N__12420\,
            I => \N__12414\
        );

    \I__1946\ : CascadeBuf
    port map (
            O => \N__12417\,
            I => \N__12411\
        );

    \I__1945\ : CascadeBuf
    port map (
            O => \N__12414\,
            I => \N__12408\
        );

    \I__1944\ : CascadeMux
    port map (
            O => \N__12411\,
            I => \N__12405\
        );

    \I__1943\ : CascadeMux
    port map (
            O => \N__12408\,
            I => \N__12402\
        );

    \I__1942\ : CascadeBuf
    port map (
            O => \N__12405\,
            I => \N__12399\
        );

    \I__1941\ : CascadeBuf
    port map (
            O => \N__12402\,
            I => \N__12396\
        );

    \I__1940\ : CascadeMux
    port map (
            O => \N__12399\,
            I => \N__12393\
        );

    \I__1939\ : CascadeMux
    port map (
            O => \N__12396\,
            I => \N__12390\
        );

    \I__1938\ : CascadeBuf
    port map (
            O => \N__12393\,
            I => \N__12387\
        );

    \I__1937\ : CascadeBuf
    port map (
            O => \N__12390\,
            I => \N__12384\
        );

    \I__1936\ : CascadeMux
    port map (
            O => \N__12387\,
            I => \N__12381\
        );

    \I__1935\ : CascadeMux
    port map (
            O => \N__12384\,
            I => \N__12378\
        );

    \I__1934\ : CascadeBuf
    port map (
            O => \N__12381\,
            I => \N__12375\
        );

    \I__1933\ : CascadeBuf
    port map (
            O => \N__12378\,
            I => \N__12372\
        );

    \I__1932\ : CascadeMux
    port map (
            O => \N__12375\,
            I => \N__12369\
        );

    \I__1931\ : CascadeMux
    port map (
            O => \N__12372\,
            I => \N__12366\
        );

    \I__1930\ : CascadeBuf
    port map (
            O => \N__12369\,
            I => \N__12363\
        );

    \I__1929\ : CascadeBuf
    port map (
            O => \N__12366\,
            I => \N__12360\
        );

    \I__1928\ : CascadeMux
    port map (
            O => \N__12363\,
            I => \N__12357\
        );

    \I__1927\ : CascadeMux
    port map (
            O => \N__12360\,
            I => \N__12354\
        );

    \I__1926\ : CascadeBuf
    port map (
            O => \N__12357\,
            I => \N__12351\
        );

    \I__1925\ : CascadeBuf
    port map (
            O => \N__12354\,
            I => \N__12348\
        );

    \I__1924\ : CascadeMux
    port map (
            O => \N__12351\,
            I => \N__12345\
        );

    \I__1923\ : CascadeMux
    port map (
            O => \N__12348\,
            I => \N__12342\
        );

    \I__1922\ : CascadeBuf
    port map (
            O => \N__12345\,
            I => \N__12339\
        );

    \I__1921\ : CascadeBuf
    port map (
            O => \N__12342\,
            I => \N__12336\
        );

    \I__1920\ : CascadeMux
    port map (
            O => \N__12339\,
            I => \N__12333\
        );

    \I__1919\ : CascadeMux
    port map (
            O => \N__12336\,
            I => \N__12330\
        );

    \I__1918\ : CascadeBuf
    port map (
            O => \N__12333\,
            I => \N__12327\
        );

    \I__1917\ : CascadeBuf
    port map (
            O => \N__12330\,
            I => \N__12324\
        );

    \I__1916\ : CascadeMux
    port map (
            O => \N__12327\,
            I => \N__12321\
        );

    \I__1915\ : CascadeMux
    port map (
            O => \N__12324\,
            I => \N__12318\
        );

    \I__1914\ : CascadeBuf
    port map (
            O => \N__12321\,
            I => \N__12315\
        );

    \I__1913\ : CascadeBuf
    port map (
            O => \N__12318\,
            I => \N__12312\
        );

    \I__1912\ : CascadeMux
    port map (
            O => \N__12315\,
            I => \N__12309\
        );

    \I__1911\ : CascadeMux
    port map (
            O => \N__12312\,
            I => \N__12306\
        );

    \I__1910\ : CascadeBuf
    port map (
            O => \N__12309\,
            I => \N__12303\
        );

    \I__1909\ : CascadeBuf
    port map (
            O => \N__12306\,
            I => \N__12300\
        );

    \I__1908\ : CascadeMux
    port map (
            O => \N__12303\,
            I => \N__12297\
        );

    \I__1907\ : CascadeMux
    port map (
            O => \N__12300\,
            I => \N__12294\
        );

    \I__1906\ : InMux
    port map (
            O => \N__12297\,
            I => \N__12291\
        );

    \I__1905\ : CascadeBuf
    port map (
            O => \N__12294\,
            I => \N__12288\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__12291\,
            I => \N__12285\
        );

    \I__1903\ : CascadeMux
    port map (
            O => \N__12288\,
            I => \N__12282\
        );

    \I__1902\ : Span4Mux_s1_v
    port map (
            O => \N__12285\,
            I => \N__12279\
        );

    \I__1901\ : InMux
    port map (
            O => \N__12282\,
            I => \N__12276\
        );

    \I__1900\ : Span4Mux_h
    port map (
            O => \N__12279\,
            I => \N__12273\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__12276\,
            I => \N__12270\
        );

    \I__1898\ : Sp12to4
    port map (
            O => \N__12273\,
            I => \N__12267\
        );

    \I__1897\ : Sp12to4
    port map (
            O => \N__12270\,
            I => \N__12264\
        );

    \I__1896\ : Span12Mux_s9_v
    port map (
            O => \N__12267\,
            I => \N__12261\
        );

    \I__1895\ : Span12Mux_s9_v
    port map (
            O => \N__12264\,
            I => \N__12258\
        );

    \I__1894\ : Span12Mux_v
    port map (
            O => \N__12261\,
            I => \N__12253\
        );

    \I__1893\ : Span12Mux_v
    port map (
            O => \N__12258\,
            I => \N__12253\
        );

    \I__1892\ : Odrv12
    port map (
            O => \N__12253\,
            I => \RX_ADDR_6\
        );

    \I__1891\ : InMux
    port map (
            O => \N__12250\,
            I => \N__12247\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__12247\,
            I => \receive_module.O_X_7\
        );

    \I__1889\ : CascadeMux
    port map (
            O => \N__12244\,
            I => \N__12241\
        );

    \I__1888\ : InMux
    port map (
            O => \N__12241\,
            I => \N__12238\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__12238\,
            I => \N__12231\
        );

    \I__1886\ : InMux
    port map (
            O => \N__12237\,
            I => \N__12222\
        );

    \I__1885\ : InMux
    port map (
            O => \N__12236\,
            I => \N__12222\
        );

    \I__1884\ : InMux
    port map (
            O => \N__12235\,
            I => \N__12222\
        );

    \I__1883\ : InMux
    port map (
            O => \N__12234\,
            I => \N__12222\
        );

    \I__1882\ : Span4Mux_h
    port map (
            O => \N__12231\,
            I => \N__12219\
        );

    \I__1881\ : LocalMux
    port map (
            O => \N__12222\,
            I => \receive_module.O_Y_1\
        );

    \I__1880\ : Odrv4
    port map (
            O => \N__12219\,
            I => \receive_module.O_Y_1\
        );

    \I__1879\ : CascadeMux
    port map (
            O => \N__12214\,
            I => \N__12210\
        );

    \I__1878\ : CascadeMux
    port map (
            O => \N__12213\,
            I => \N__12207\
        );

    \I__1877\ : CascadeBuf
    port map (
            O => \N__12210\,
            I => \N__12204\
        );

    \I__1876\ : CascadeBuf
    port map (
            O => \N__12207\,
            I => \N__12201\
        );

    \I__1875\ : CascadeMux
    port map (
            O => \N__12204\,
            I => \N__12198\
        );

    \I__1874\ : CascadeMux
    port map (
            O => \N__12201\,
            I => \N__12195\
        );

    \I__1873\ : CascadeBuf
    port map (
            O => \N__12198\,
            I => \N__12192\
        );

    \I__1872\ : CascadeBuf
    port map (
            O => \N__12195\,
            I => \N__12189\
        );

    \I__1871\ : CascadeMux
    port map (
            O => \N__12192\,
            I => \N__12186\
        );

    \I__1870\ : CascadeMux
    port map (
            O => \N__12189\,
            I => \N__12183\
        );

    \I__1869\ : CascadeBuf
    port map (
            O => \N__12186\,
            I => \N__12180\
        );

    \I__1868\ : CascadeBuf
    port map (
            O => \N__12183\,
            I => \N__12177\
        );

    \I__1867\ : CascadeMux
    port map (
            O => \N__12180\,
            I => \N__12174\
        );

    \I__1866\ : CascadeMux
    port map (
            O => \N__12177\,
            I => \N__12171\
        );

    \I__1865\ : CascadeBuf
    port map (
            O => \N__12174\,
            I => \N__12168\
        );

    \I__1864\ : CascadeBuf
    port map (
            O => \N__12171\,
            I => \N__12165\
        );

    \I__1863\ : CascadeMux
    port map (
            O => \N__12168\,
            I => \N__12162\
        );

    \I__1862\ : CascadeMux
    port map (
            O => \N__12165\,
            I => \N__12159\
        );

    \I__1861\ : CascadeBuf
    port map (
            O => \N__12162\,
            I => \N__12156\
        );

    \I__1860\ : CascadeBuf
    port map (
            O => \N__12159\,
            I => \N__12153\
        );

    \I__1859\ : CascadeMux
    port map (
            O => \N__12156\,
            I => \N__12150\
        );

    \I__1858\ : CascadeMux
    port map (
            O => \N__12153\,
            I => \N__12147\
        );

    \I__1857\ : CascadeBuf
    port map (
            O => \N__12150\,
            I => \N__12144\
        );

    \I__1856\ : CascadeBuf
    port map (
            O => \N__12147\,
            I => \N__12141\
        );

    \I__1855\ : CascadeMux
    port map (
            O => \N__12144\,
            I => \N__12138\
        );

    \I__1854\ : CascadeMux
    port map (
            O => \N__12141\,
            I => \N__12135\
        );

    \I__1853\ : CascadeBuf
    port map (
            O => \N__12138\,
            I => \N__12132\
        );

    \I__1852\ : CascadeBuf
    port map (
            O => \N__12135\,
            I => \N__12129\
        );

    \I__1851\ : CascadeMux
    port map (
            O => \N__12132\,
            I => \N__12126\
        );

    \I__1850\ : CascadeMux
    port map (
            O => \N__12129\,
            I => \N__12123\
        );

    \I__1849\ : CascadeBuf
    port map (
            O => \N__12126\,
            I => \N__12120\
        );

    \I__1848\ : CascadeBuf
    port map (
            O => \N__12123\,
            I => \N__12117\
        );

    \I__1847\ : CascadeMux
    port map (
            O => \N__12120\,
            I => \N__12114\
        );

    \I__1846\ : CascadeMux
    port map (
            O => \N__12117\,
            I => \N__12111\
        );

    \I__1845\ : CascadeBuf
    port map (
            O => \N__12114\,
            I => \N__12108\
        );

    \I__1844\ : CascadeBuf
    port map (
            O => \N__12111\,
            I => \N__12105\
        );

    \I__1843\ : CascadeMux
    port map (
            O => \N__12108\,
            I => \N__12102\
        );

    \I__1842\ : CascadeMux
    port map (
            O => \N__12105\,
            I => \N__12099\
        );

    \I__1841\ : CascadeBuf
    port map (
            O => \N__12102\,
            I => \N__12096\
        );

    \I__1840\ : CascadeBuf
    port map (
            O => \N__12099\,
            I => \N__12093\
        );

    \I__1839\ : CascadeMux
    port map (
            O => \N__12096\,
            I => \N__12090\
        );

    \I__1838\ : CascadeMux
    port map (
            O => \N__12093\,
            I => \N__12087\
        );

    \I__1837\ : CascadeBuf
    port map (
            O => \N__12090\,
            I => \N__12084\
        );

    \I__1836\ : CascadeBuf
    port map (
            O => \N__12087\,
            I => \N__12081\
        );

    \I__1835\ : CascadeMux
    port map (
            O => \N__12084\,
            I => \N__12078\
        );

    \I__1834\ : CascadeMux
    port map (
            O => \N__12081\,
            I => \N__12075\
        );

    \I__1833\ : CascadeBuf
    port map (
            O => \N__12078\,
            I => \N__12072\
        );

    \I__1832\ : CascadeBuf
    port map (
            O => \N__12075\,
            I => \N__12069\
        );

    \I__1831\ : CascadeMux
    port map (
            O => \N__12072\,
            I => \N__12066\
        );

    \I__1830\ : CascadeMux
    port map (
            O => \N__12069\,
            I => \N__12063\
        );

    \I__1829\ : CascadeBuf
    port map (
            O => \N__12066\,
            I => \N__12060\
        );

    \I__1828\ : CascadeBuf
    port map (
            O => \N__12063\,
            I => \N__12057\
        );

    \I__1827\ : CascadeMux
    port map (
            O => \N__12060\,
            I => \N__12054\
        );

    \I__1826\ : CascadeMux
    port map (
            O => \N__12057\,
            I => \N__12051\
        );

    \I__1825\ : CascadeBuf
    port map (
            O => \N__12054\,
            I => \N__12048\
        );

    \I__1824\ : CascadeBuf
    port map (
            O => \N__12051\,
            I => \N__12045\
        );

    \I__1823\ : CascadeMux
    port map (
            O => \N__12048\,
            I => \N__12042\
        );

    \I__1822\ : CascadeMux
    port map (
            O => \N__12045\,
            I => \N__12039\
        );

    \I__1821\ : CascadeBuf
    port map (
            O => \N__12042\,
            I => \N__12036\
        );

    \I__1820\ : CascadeBuf
    port map (
            O => \N__12039\,
            I => \N__12033\
        );

    \I__1819\ : CascadeMux
    port map (
            O => \N__12036\,
            I => \N__12030\
        );

    \I__1818\ : CascadeMux
    port map (
            O => \N__12033\,
            I => \N__12027\
        );

    \I__1817\ : InMux
    port map (
            O => \N__12030\,
            I => \N__12024\
        );

    \I__1816\ : InMux
    port map (
            O => \N__12027\,
            I => \N__12021\
        );

    \I__1815\ : LocalMux
    port map (
            O => \N__12024\,
            I => \N__12018\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__12021\,
            I => \N__12015\
        );

    \I__1813\ : Span12Mux_v
    port map (
            O => \N__12018\,
            I => \N__12012\
        );

    \I__1812\ : Span12Mux_s9_v
    port map (
            O => \N__12015\,
            I => \N__12009\
        );

    \I__1811\ : Span12Mux_h
    port map (
            O => \N__12012\,
            I => \N__12006\
        );

    \I__1810\ : Span12Mux_v
    port map (
            O => \N__12009\,
            I => \N__12003\
        );

    \I__1809\ : Odrv12
    port map (
            O => \N__12006\,
            I => \RX_ADDR_7\
        );

    \I__1808\ : Odrv12
    port map (
            O => \N__12003\,
            I => \RX_ADDR_7\
        );

    \I__1807\ : InMux
    port map (
            O => \N__11998\,
            I => \receive_module.n3699\
        );

    \I__1806\ : InMux
    port map (
            O => \N__11995\,
            I => \N__11992\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__11992\,
            I => \N__11989\
        );

    \I__1804\ : Span4Mux_v
    port map (
            O => \N__11989\,
            I => \N__11983\
        );

    \I__1803\ : InMux
    port map (
            O => \N__11988\,
            I => \N__11978\
        );

    \I__1802\ : InMux
    port map (
            O => \N__11987\,
            I => \N__11978\
        );

    \I__1801\ : InMux
    port map (
            O => \N__11986\,
            I => \N__11975\
        );

    \I__1800\ : Odrv4
    port map (
            O => \N__11983\,
            I => \receive_module.O_Y_2\
        );

    \I__1799\ : LocalMux
    port map (
            O => \N__11978\,
            I => \receive_module.O_Y_2\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__11975\,
            I => \receive_module.O_Y_2\
        );

    \I__1797\ : CascadeMux
    port map (
            O => \N__11968\,
            I => \N__11965\
        );

    \I__1796\ : InMux
    port map (
            O => \N__11965\,
            I => \N__11962\
        );

    \I__1795\ : LocalMux
    port map (
            O => \N__11962\,
            I => \receive_module.O_X_8\
        );

    \I__1794\ : CascadeMux
    port map (
            O => \N__11959\,
            I => \N__11955\
        );

    \I__1793\ : CascadeMux
    port map (
            O => \N__11958\,
            I => \N__11952\
        );

    \I__1792\ : CascadeBuf
    port map (
            O => \N__11955\,
            I => \N__11949\
        );

    \I__1791\ : CascadeBuf
    port map (
            O => \N__11952\,
            I => \N__11946\
        );

    \I__1790\ : CascadeMux
    port map (
            O => \N__11949\,
            I => \N__11943\
        );

    \I__1789\ : CascadeMux
    port map (
            O => \N__11946\,
            I => \N__11940\
        );

    \I__1788\ : CascadeBuf
    port map (
            O => \N__11943\,
            I => \N__11937\
        );

    \I__1787\ : CascadeBuf
    port map (
            O => \N__11940\,
            I => \N__11934\
        );

    \I__1786\ : CascadeMux
    port map (
            O => \N__11937\,
            I => \N__11931\
        );

    \I__1785\ : CascadeMux
    port map (
            O => \N__11934\,
            I => \N__11928\
        );

    \I__1784\ : CascadeBuf
    port map (
            O => \N__11931\,
            I => \N__11925\
        );

    \I__1783\ : CascadeBuf
    port map (
            O => \N__11928\,
            I => \N__11922\
        );

    \I__1782\ : CascadeMux
    port map (
            O => \N__11925\,
            I => \N__11919\
        );

    \I__1781\ : CascadeMux
    port map (
            O => \N__11922\,
            I => \N__11916\
        );

    \I__1780\ : CascadeBuf
    port map (
            O => \N__11919\,
            I => \N__11913\
        );

    \I__1779\ : CascadeBuf
    port map (
            O => \N__11916\,
            I => \N__11910\
        );

    \I__1778\ : CascadeMux
    port map (
            O => \N__11913\,
            I => \N__11907\
        );

    \I__1777\ : CascadeMux
    port map (
            O => \N__11910\,
            I => \N__11904\
        );

    \I__1776\ : CascadeBuf
    port map (
            O => \N__11907\,
            I => \N__11901\
        );

    \I__1775\ : CascadeBuf
    port map (
            O => \N__11904\,
            I => \N__11898\
        );

    \I__1774\ : CascadeMux
    port map (
            O => \N__11901\,
            I => \N__11895\
        );

    \I__1773\ : CascadeMux
    port map (
            O => \N__11898\,
            I => \N__11892\
        );

    \I__1772\ : CascadeBuf
    port map (
            O => \N__11895\,
            I => \N__11889\
        );

    \I__1771\ : CascadeBuf
    port map (
            O => \N__11892\,
            I => \N__11886\
        );

    \I__1770\ : CascadeMux
    port map (
            O => \N__11889\,
            I => \N__11883\
        );

    \I__1769\ : CascadeMux
    port map (
            O => \N__11886\,
            I => \N__11880\
        );

    \I__1768\ : CascadeBuf
    port map (
            O => \N__11883\,
            I => \N__11877\
        );

    \I__1767\ : CascadeBuf
    port map (
            O => \N__11880\,
            I => \N__11874\
        );

    \I__1766\ : CascadeMux
    port map (
            O => \N__11877\,
            I => \N__11871\
        );

    \I__1765\ : CascadeMux
    port map (
            O => \N__11874\,
            I => \N__11868\
        );

    \I__1764\ : CascadeBuf
    port map (
            O => \N__11871\,
            I => \N__11865\
        );

    \I__1763\ : CascadeBuf
    port map (
            O => \N__11868\,
            I => \N__11862\
        );

    \I__1762\ : CascadeMux
    port map (
            O => \N__11865\,
            I => \N__11859\
        );

    \I__1761\ : CascadeMux
    port map (
            O => \N__11862\,
            I => \N__11856\
        );

    \I__1760\ : CascadeBuf
    port map (
            O => \N__11859\,
            I => \N__11853\
        );

    \I__1759\ : CascadeBuf
    port map (
            O => \N__11856\,
            I => \N__11850\
        );

    \I__1758\ : CascadeMux
    port map (
            O => \N__11853\,
            I => \N__11847\
        );

    \I__1757\ : CascadeMux
    port map (
            O => \N__11850\,
            I => \N__11844\
        );

    \I__1756\ : CascadeBuf
    port map (
            O => \N__11847\,
            I => \N__11841\
        );

    \I__1755\ : CascadeBuf
    port map (
            O => \N__11844\,
            I => \N__11838\
        );

    \I__1754\ : CascadeMux
    port map (
            O => \N__11841\,
            I => \N__11835\
        );

    \I__1753\ : CascadeMux
    port map (
            O => \N__11838\,
            I => \N__11832\
        );

    \I__1752\ : CascadeBuf
    port map (
            O => \N__11835\,
            I => \N__11829\
        );

    \I__1751\ : CascadeBuf
    port map (
            O => \N__11832\,
            I => \N__11826\
        );

    \I__1750\ : CascadeMux
    port map (
            O => \N__11829\,
            I => \N__11823\
        );

    \I__1749\ : CascadeMux
    port map (
            O => \N__11826\,
            I => \N__11820\
        );

    \I__1748\ : CascadeBuf
    port map (
            O => \N__11823\,
            I => \N__11817\
        );

    \I__1747\ : CascadeBuf
    port map (
            O => \N__11820\,
            I => \N__11814\
        );

    \I__1746\ : CascadeMux
    port map (
            O => \N__11817\,
            I => \N__11811\
        );

    \I__1745\ : CascadeMux
    port map (
            O => \N__11814\,
            I => \N__11808\
        );

    \I__1744\ : CascadeBuf
    port map (
            O => \N__11811\,
            I => \N__11805\
        );

    \I__1743\ : CascadeBuf
    port map (
            O => \N__11808\,
            I => \N__11802\
        );

    \I__1742\ : CascadeMux
    port map (
            O => \N__11805\,
            I => \N__11799\
        );

    \I__1741\ : CascadeMux
    port map (
            O => \N__11802\,
            I => \N__11796\
        );

    \I__1740\ : CascadeBuf
    port map (
            O => \N__11799\,
            I => \N__11793\
        );

    \I__1739\ : CascadeBuf
    port map (
            O => \N__11796\,
            I => \N__11790\
        );

    \I__1738\ : CascadeMux
    port map (
            O => \N__11793\,
            I => \N__11787\
        );

    \I__1737\ : CascadeMux
    port map (
            O => \N__11790\,
            I => \N__11784\
        );

    \I__1736\ : CascadeBuf
    port map (
            O => \N__11787\,
            I => \N__11781\
        );

    \I__1735\ : CascadeBuf
    port map (
            O => \N__11784\,
            I => \N__11778\
        );

    \I__1734\ : CascadeMux
    port map (
            O => \N__11781\,
            I => \N__11775\
        );

    \I__1733\ : CascadeMux
    port map (
            O => \N__11778\,
            I => \N__11772\
        );

    \I__1732\ : InMux
    port map (
            O => \N__11775\,
            I => \N__11769\
        );

    \I__1731\ : InMux
    port map (
            O => \N__11772\,
            I => \N__11766\
        );

    \I__1730\ : LocalMux
    port map (
            O => \N__11769\,
            I => \N__11763\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__11766\,
            I => \N__11760\
        );

    \I__1728\ : Span4Mux_s1_v
    port map (
            O => \N__11763\,
            I => \N__11757\
        );

    \I__1727\ : Span12Mux_s7_v
    port map (
            O => \N__11760\,
            I => \N__11754\
        );

    \I__1726\ : Span4Mux_h
    port map (
            O => \N__11757\,
            I => \N__11751\
        );

    \I__1725\ : Span12Mux_h
    port map (
            O => \N__11754\,
            I => \N__11748\
        );

    \I__1724\ : Sp12to4
    port map (
            O => \N__11751\,
            I => \N__11745\
        );

    \I__1723\ : Span12Mux_v
    port map (
            O => \N__11748\,
            I => \N__11742\
        );

    \I__1722\ : Span12Mux_s11_v
    port map (
            O => \N__11745\,
            I => \N__11739\
        );

    \I__1721\ : Odrv12
    port map (
            O => \N__11742\,
            I => \RX_ADDR_8\
        );

    \I__1720\ : Odrv12
    port map (
            O => \N__11739\,
            I => \RX_ADDR_8\
        );

    \I__1719\ : InMux
    port map (
            O => \N__11734\,
            I => \receive_module.n3700\
        );

    \I__1718\ : InMux
    port map (
            O => \N__11731\,
            I => \N__11728\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__11728\,
            I => \transmit_module.ADDR_Y_COMPONENT_10\
        );

    \I__1716\ : InMux
    port map (
            O => \N__11725\,
            I => \N__11722\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__11722\,
            I => \N__11719\
        );

    \I__1714\ : Span4Mux_v
    port map (
            O => \N__11719\,
            I => \N__11716\
        );

    \I__1713\ : Odrv4
    port map (
            O => \N__11716\,
            I => \transmit_module.n209\
        );

    \I__1712\ : InMux
    port map (
            O => \N__11713\,
            I => \N__11710\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__11710\,
            I => \N__11706\
        );

    \I__1710\ : InMux
    port map (
            O => \N__11709\,
            I => \N__11703\
        );

    \I__1709\ : Span4Mux_v
    port map (
            O => \N__11706\,
            I => \N__11700\
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__11703\,
            I => \transmit_module.n178\
        );

    \I__1707\ : Odrv4
    port map (
            O => \N__11700\,
            I => \transmit_module.n178\
        );

    \I__1706\ : CascadeMux
    port map (
            O => \N__11695\,
            I => \transmit_module.n209_cascade_\
        );

    \I__1705\ : CEMux
    port map (
            O => \N__11692\,
            I => \N__11688\
        );

    \I__1704\ : CEMux
    port map (
            O => \N__11691\,
            I => \N__11685\
        );

    \I__1703\ : LocalMux
    port map (
            O => \N__11688\,
            I => \N__11682\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__11685\,
            I => \N__11679\
        );

    \I__1701\ : Span4Mux_h
    port map (
            O => \N__11682\,
            I => \N__11676\
        );

    \I__1700\ : Span4Mux_h
    port map (
            O => \N__11679\,
            I => \N__11673\
        );

    \I__1699\ : Odrv4
    port map (
            O => \N__11676\,
            I => n2283
        );

    \I__1698\ : Odrv4
    port map (
            O => \N__11673\,
            I => n2283
        );

    \I__1697\ : InMux
    port map (
            O => \N__11668\,
            I => \N__11665\
        );

    \I__1696\ : LocalMux
    port map (
            O => \N__11665\,
            I => \old_HS\
        );

    \I__1695\ : CascadeMux
    port map (
            O => \N__11662\,
            I => \N__11659\
        );

    \I__1694\ : CascadeBuf
    port map (
            O => \N__11659\,
            I => \N__11656\
        );

    \I__1693\ : CascadeMux
    port map (
            O => \N__11656\,
            I => \N__11652\
        );

    \I__1692\ : CascadeMux
    port map (
            O => \N__11655\,
            I => \N__11649\
        );

    \I__1691\ : CascadeBuf
    port map (
            O => \N__11652\,
            I => \N__11646\
        );

    \I__1690\ : CascadeBuf
    port map (
            O => \N__11649\,
            I => \N__11643\
        );

    \I__1689\ : CascadeMux
    port map (
            O => \N__11646\,
            I => \N__11640\
        );

    \I__1688\ : CascadeMux
    port map (
            O => \N__11643\,
            I => \N__11637\
        );

    \I__1687\ : CascadeBuf
    port map (
            O => \N__11640\,
            I => \N__11634\
        );

    \I__1686\ : CascadeBuf
    port map (
            O => \N__11637\,
            I => \N__11631\
        );

    \I__1685\ : CascadeMux
    port map (
            O => \N__11634\,
            I => \N__11628\
        );

    \I__1684\ : CascadeMux
    port map (
            O => \N__11631\,
            I => \N__11625\
        );

    \I__1683\ : CascadeBuf
    port map (
            O => \N__11628\,
            I => \N__11622\
        );

    \I__1682\ : CascadeBuf
    port map (
            O => \N__11625\,
            I => \N__11619\
        );

    \I__1681\ : CascadeMux
    port map (
            O => \N__11622\,
            I => \N__11616\
        );

    \I__1680\ : CascadeMux
    port map (
            O => \N__11619\,
            I => \N__11613\
        );

    \I__1679\ : CascadeBuf
    port map (
            O => \N__11616\,
            I => \N__11610\
        );

    \I__1678\ : CascadeBuf
    port map (
            O => \N__11613\,
            I => \N__11607\
        );

    \I__1677\ : CascadeMux
    port map (
            O => \N__11610\,
            I => \N__11604\
        );

    \I__1676\ : CascadeMux
    port map (
            O => \N__11607\,
            I => \N__11601\
        );

    \I__1675\ : CascadeBuf
    port map (
            O => \N__11604\,
            I => \N__11598\
        );

    \I__1674\ : CascadeBuf
    port map (
            O => \N__11601\,
            I => \N__11595\
        );

    \I__1673\ : CascadeMux
    port map (
            O => \N__11598\,
            I => \N__11592\
        );

    \I__1672\ : CascadeMux
    port map (
            O => \N__11595\,
            I => \N__11589\
        );

    \I__1671\ : CascadeBuf
    port map (
            O => \N__11592\,
            I => \N__11586\
        );

    \I__1670\ : CascadeBuf
    port map (
            O => \N__11589\,
            I => \N__11583\
        );

    \I__1669\ : CascadeMux
    port map (
            O => \N__11586\,
            I => \N__11580\
        );

    \I__1668\ : CascadeMux
    port map (
            O => \N__11583\,
            I => \N__11577\
        );

    \I__1667\ : CascadeBuf
    port map (
            O => \N__11580\,
            I => \N__11574\
        );

    \I__1666\ : CascadeBuf
    port map (
            O => \N__11577\,
            I => \N__11571\
        );

    \I__1665\ : CascadeMux
    port map (
            O => \N__11574\,
            I => \N__11568\
        );

    \I__1664\ : CascadeMux
    port map (
            O => \N__11571\,
            I => \N__11565\
        );

    \I__1663\ : CascadeBuf
    port map (
            O => \N__11568\,
            I => \N__11562\
        );

    \I__1662\ : CascadeBuf
    port map (
            O => \N__11565\,
            I => \N__11559\
        );

    \I__1661\ : CascadeMux
    port map (
            O => \N__11562\,
            I => \N__11556\
        );

    \I__1660\ : CascadeMux
    port map (
            O => \N__11559\,
            I => \N__11553\
        );

    \I__1659\ : CascadeBuf
    port map (
            O => \N__11556\,
            I => \N__11550\
        );

    \I__1658\ : CascadeBuf
    port map (
            O => \N__11553\,
            I => \N__11547\
        );

    \I__1657\ : CascadeMux
    port map (
            O => \N__11550\,
            I => \N__11544\
        );

    \I__1656\ : CascadeMux
    port map (
            O => \N__11547\,
            I => \N__11541\
        );

    \I__1655\ : CascadeBuf
    port map (
            O => \N__11544\,
            I => \N__11538\
        );

    \I__1654\ : CascadeBuf
    port map (
            O => \N__11541\,
            I => \N__11535\
        );

    \I__1653\ : CascadeMux
    port map (
            O => \N__11538\,
            I => \N__11532\
        );

    \I__1652\ : CascadeMux
    port map (
            O => \N__11535\,
            I => \N__11529\
        );

    \I__1651\ : CascadeBuf
    port map (
            O => \N__11532\,
            I => \N__11526\
        );

    \I__1650\ : CascadeBuf
    port map (
            O => \N__11529\,
            I => \N__11523\
        );

    \I__1649\ : CascadeMux
    port map (
            O => \N__11526\,
            I => \N__11520\
        );

    \I__1648\ : CascadeMux
    port map (
            O => \N__11523\,
            I => \N__11517\
        );

    \I__1647\ : CascadeBuf
    port map (
            O => \N__11520\,
            I => \N__11514\
        );

    \I__1646\ : CascadeBuf
    port map (
            O => \N__11517\,
            I => \N__11511\
        );

    \I__1645\ : CascadeMux
    port map (
            O => \N__11514\,
            I => \N__11508\
        );

    \I__1644\ : CascadeMux
    port map (
            O => \N__11511\,
            I => \N__11505\
        );

    \I__1643\ : CascadeBuf
    port map (
            O => \N__11508\,
            I => \N__11502\
        );

    \I__1642\ : CascadeBuf
    port map (
            O => \N__11505\,
            I => \N__11499\
        );

    \I__1641\ : CascadeMux
    port map (
            O => \N__11502\,
            I => \N__11496\
        );

    \I__1640\ : CascadeMux
    port map (
            O => \N__11499\,
            I => \N__11493\
        );

    \I__1639\ : CascadeBuf
    port map (
            O => \N__11496\,
            I => \N__11490\
        );

    \I__1638\ : CascadeBuf
    port map (
            O => \N__11493\,
            I => \N__11487\
        );

    \I__1637\ : CascadeMux
    port map (
            O => \N__11490\,
            I => \N__11484\
        );

    \I__1636\ : CascadeMux
    port map (
            O => \N__11487\,
            I => \N__11481\
        );

    \I__1635\ : InMux
    port map (
            O => \N__11484\,
            I => \N__11478\
        );

    \I__1634\ : CascadeBuf
    port map (
            O => \N__11481\,
            I => \N__11475\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__11478\,
            I => \N__11472\
        );

    \I__1632\ : CascadeMux
    port map (
            O => \N__11475\,
            I => \N__11469\
        );

    \I__1631\ : Span4Mux_s2_v
    port map (
            O => \N__11472\,
            I => \N__11466\
        );

    \I__1630\ : InMux
    port map (
            O => \N__11469\,
            I => \N__11463\
        );

    \I__1629\ : Span4Mux_h
    port map (
            O => \N__11466\,
            I => \N__11460\
        );

    \I__1628\ : LocalMux
    port map (
            O => \N__11463\,
            I => \N__11457\
        );

    \I__1627\ : Sp12to4
    port map (
            O => \N__11460\,
            I => \N__11454\
        );

    \I__1626\ : Span4Mux_s2_v
    port map (
            O => \N__11457\,
            I => \N__11451\
        );

    \I__1625\ : Span12Mux_s10_v
    port map (
            O => \N__11454\,
            I => \N__11448\
        );

    \I__1624\ : Sp12to4
    port map (
            O => \N__11451\,
            I => \N__11445\
        );

    \I__1623\ : Span12Mux_h
    port map (
            O => \N__11448\,
            I => \N__11440\
        );

    \I__1622\ : Span12Mux_s10_v
    port map (
            O => \N__11445\,
            I => \N__11440\
        );

    \I__1621\ : Span12Mux_v
    port map (
            O => \N__11440\,
            I => \N__11437\
        );

    \I__1620\ : Odrv12
    port map (
            O => \N__11437\,
            I => \RX_ADDR_3\
        );

    \I__1619\ : InMux
    port map (
            O => \N__11434\,
            I => \bfn_13_10_0_\
        );

    \I__1618\ : CascadeMux
    port map (
            O => \N__11431\,
            I => \N__11428\
        );

    \I__1617\ : CascadeBuf
    port map (
            O => \N__11428\,
            I => \N__11424\
        );

    \I__1616\ : CascadeMux
    port map (
            O => \N__11427\,
            I => \N__11421\
        );

    \I__1615\ : CascadeMux
    port map (
            O => \N__11424\,
            I => \N__11418\
        );

    \I__1614\ : CascadeBuf
    port map (
            O => \N__11421\,
            I => \N__11415\
        );

    \I__1613\ : CascadeBuf
    port map (
            O => \N__11418\,
            I => \N__11412\
        );

    \I__1612\ : CascadeMux
    port map (
            O => \N__11415\,
            I => \N__11409\
        );

    \I__1611\ : CascadeMux
    port map (
            O => \N__11412\,
            I => \N__11406\
        );

    \I__1610\ : CascadeBuf
    port map (
            O => \N__11409\,
            I => \N__11403\
        );

    \I__1609\ : CascadeBuf
    port map (
            O => \N__11406\,
            I => \N__11400\
        );

    \I__1608\ : CascadeMux
    port map (
            O => \N__11403\,
            I => \N__11397\
        );

    \I__1607\ : CascadeMux
    port map (
            O => \N__11400\,
            I => \N__11394\
        );

    \I__1606\ : CascadeBuf
    port map (
            O => \N__11397\,
            I => \N__11391\
        );

    \I__1605\ : CascadeBuf
    port map (
            O => \N__11394\,
            I => \N__11388\
        );

    \I__1604\ : CascadeMux
    port map (
            O => \N__11391\,
            I => \N__11385\
        );

    \I__1603\ : CascadeMux
    port map (
            O => \N__11388\,
            I => \N__11382\
        );

    \I__1602\ : CascadeBuf
    port map (
            O => \N__11385\,
            I => \N__11379\
        );

    \I__1601\ : CascadeBuf
    port map (
            O => \N__11382\,
            I => \N__11376\
        );

    \I__1600\ : CascadeMux
    port map (
            O => \N__11379\,
            I => \N__11373\
        );

    \I__1599\ : CascadeMux
    port map (
            O => \N__11376\,
            I => \N__11370\
        );

    \I__1598\ : CascadeBuf
    port map (
            O => \N__11373\,
            I => \N__11367\
        );

    \I__1597\ : CascadeBuf
    port map (
            O => \N__11370\,
            I => \N__11364\
        );

    \I__1596\ : CascadeMux
    port map (
            O => \N__11367\,
            I => \N__11361\
        );

    \I__1595\ : CascadeMux
    port map (
            O => \N__11364\,
            I => \N__11358\
        );

    \I__1594\ : CascadeBuf
    port map (
            O => \N__11361\,
            I => \N__11355\
        );

    \I__1593\ : CascadeBuf
    port map (
            O => \N__11358\,
            I => \N__11352\
        );

    \I__1592\ : CascadeMux
    port map (
            O => \N__11355\,
            I => \N__11349\
        );

    \I__1591\ : CascadeMux
    port map (
            O => \N__11352\,
            I => \N__11346\
        );

    \I__1590\ : CascadeBuf
    port map (
            O => \N__11349\,
            I => \N__11343\
        );

    \I__1589\ : CascadeBuf
    port map (
            O => \N__11346\,
            I => \N__11340\
        );

    \I__1588\ : CascadeMux
    port map (
            O => \N__11343\,
            I => \N__11337\
        );

    \I__1587\ : CascadeMux
    port map (
            O => \N__11340\,
            I => \N__11334\
        );

    \I__1586\ : CascadeBuf
    port map (
            O => \N__11337\,
            I => \N__11331\
        );

    \I__1585\ : CascadeBuf
    port map (
            O => \N__11334\,
            I => \N__11328\
        );

    \I__1584\ : CascadeMux
    port map (
            O => \N__11331\,
            I => \N__11325\
        );

    \I__1583\ : CascadeMux
    port map (
            O => \N__11328\,
            I => \N__11322\
        );

    \I__1582\ : CascadeBuf
    port map (
            O => \N__11325\,
            I => \N__11319\
        );

    \I__1581\ : CascadeBuf
    port map (
            O => \N__11322\,
            I => \N__11316\
        );

    \I__1580\ : CascadeMux
    port map (
            O => \N__11319\,
            I => \N__11313\
        );

    \I__1579\ : CascadeMux
    port map (
            O => \N__11316\,
            I => \N__11310\
        );

    \I__1578\ : CascadeBuf
    port map (
            O => \N__11313\,
            I => \N__11307\
        );

    \I__1577\ : CascadeBuf
    port map (
            O => \N__11310\,
            I => \N__11304\
        );

    \I__1576\ : CascadeMux
    port map (
            O => \N__11307\,
            I => \N__11301\
        );

    \I__1575\ : CascadeMux
    port map (
            O => \N__11304\,
            I => \N__11298\
        );

    \I__1574\ : CascadeBuf
    port map (
            O => \N__11301\,
            I => \N__11295\
        );

    \I__1573\ : CascadeBuf
    port map (
            O => \N__11298\,
            I => \N__11292\
        );

    \I__1572\ : CascadeMux
    port map (
            O => \N__11295\,
            I => \N__11289\
        );

    \I__1571\ : CascadeMux
    port map (
            O => \N__11292\,
            I => \N__11286\
        );

    \I__1570\ : CascadeBuf
    port map (
            O => \N__11289\,
            I => \N__11283\
        );

    \I__1569\ : CascadeBuf
    port map (
            O => \N__11286\,
            I => \N__11280\
        );

    \I__1568\ : CascadeMux
    port map (
            O => \N__11283\,
            I => \N__11277\
        );

    \I__1567\ : CascadeMux
    port map (
            O => \N__11280\,
            I => \N__11274\
        );

    \I__1566\ : CascadeBuf
    port map (
            O => \N__11277\,
            I => \N__11271\
        );

    \I__1565\ : CascadeBuf
    port map (
            O => \N__11274\,
            I => \N__11268\
        );

    \I__1564\ : CascadeMux
    port map (
            O => \N__11271\,
            I => \N__11265\
        );

    \I__1563\ : CascadeMux
    port map (
            O => \N__11268\,
            I => \N__11262\
        );

    \I__1562\ : CascadeBuf
    port map (
            O => \N__11265\,
            I => \N__11259\
        );

    \I__1561\ : CascadeBuf
    port map (
            O => \N__11262\,
            I => \N__11256\
        );

    \I__1560\ : CascadeMux
    port map (
            O => \N__11259\,
            I => \N__11253\
        );

    \I__1559\ : CascadeMux
    port map (
            O => \N__11256\,
            I => \N__11250\
        );

    \I__1558\ : CascadeBuf
    port map (
            O => \N__11253\,
            I => \N__11247\
        );

    \I__1557\ : InMux
    port map (
            O => \N__11250\,
            I => \N__11244\
        );

    \I__1556\ : CascadeMux
    port map (
            O => \N__11247\,
            I => \N__11241\
        );

    \I__1555\ : LocalMux
    port map (
            O => \N__11244\,
            I => \N__11238\
        );

    \I__1554\ : InMux
    port map (
            O => \N__11241\,
            I => \N__11235\
        );

    \I__1553\ : Span12Mux_s1_v
    port map (
            O => \N__11238\,
            I => \N__11232\
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__11235\,
            I => \N__11229\
        );

    \I__1551\ : Span12Mux_h
    port map (
            O => \N__11232\,
            I => \N__11226\
        );

    \I__1550\ : Span12Mux_s10_v
    port map (
            O => \N__11229\,
            I => \N__11223\
        );

    \I__1549\ : Span12Mux_v
    port map (
            O => \N__11226\,
            I => \N__11220\
        );

    \I__1548\ : Span12Mux_v
    port map (
            O => \N__11223\,
            I => \N__11217\
        );

    \I__1547\ : Odrv12
    port map (
            O => \N__11220\,
            I => \RX_ADDR_4\
        );

    \I__1546\ : Odrv12
    port map (
            O => \N__11217\,
            I => \RX_ADDR_4\
        );

    \I__1545\ : InMux
    port map (
            O => \N__11212\,
            I => \receive_module.rx_counter.n3650\
        );

    \I__1544\ : CascadeMux
    port map (
            O => \N__11209\,
            I => \N__11205\
        );

    \I__1543\ : CascadeMux
    port map (
            O => \N__11208\,
            I => \N__11202\
        );

    \I__1542\ : CascadeBuf
    port map (
            O => \N__11205\,
            I => \N__11199\
        );

    \I__1541\ : CascadeBuf
    port map (
            O => \N__11202\,
            I => \N__11196\
        );

    \I__1540\ : CascadeMux
    port map (
            O => \N__11199\,
            I => \N__11193\
        );

    \I__1539\ : CascadeMux
    port map (
            O => \N__11196\,
            I => \N__11190\
        );

    \I__1538\ : CascadeBuf
    port map (
            O => \N__11193\,
            I => \N__11187\
        );

    \I__1537\ : CascadeBuf
    port map (
            O => \N__11190\,
            I => \N__11184\
        );

    \I__1536\ : CascadeMux
    port map (
            O => \N__11187\,
            I => \N__11181\
        );

    \I__1535\ : CascadeMux
    port map (
            O => \N__11184\,
            I => \N__11178\
        );

    \I__1534\ : CascadeBuf
    port map (
            O => \N__11181\,
            I => \N__11175\
        );

    \I__1533\ : CascadeBuf
    port map (
            O => \N__11178\,
            I => \N__11172\
        );

    \I__1532\ : CascadeMux
    port map (
            O => \N__11175\,
            I => \N__11169\
        );

    \I__1531\ : CascadeMux
    port map (
            O => \N__11172\,
            I => \N__11166\
        );

    \I__1530\ : CascadeBuf
    port map (
            O => \N__11169\,
            I => \N__11163\
        );

    \I__1529\ : CascadeBuf
    port map (
            O => \N__11166\,
            I => \N__11160\
        );

    \I__1528\ : CascadeMux
    port map (
            O => \N__11163\,
            I => \N__11157\
        );

    \I__1527\ : CascadeMux
    port map (
            O => \N__11160\,
            I => \N__11154\
        );

    \I__1526\ : CascadeBuf
    port map (
            O => \N__11157\,
            I => \N__11151\
        );

    \I__1525\ : CascadeBuf
    port map (
            O => \N__11154\,
            I => \N__11148\
        );

    \I__1524\ : CascadeMux
    port map (
            O => \N__11151\,
            I => \N__11145\
        );

    \I__1523\ : CascadeMux
    port map (
            O => \N__11148\,
            I => \N__11142\
        );

    \I__1522\ : CascadeBuf
    port map (
            O => \N__11145\,
            I => \N__11139\
        );

    \I__1521\ : CascadeBuf
    port map (
            O => \N__11142\,
            I => \N__11136\
        );

    \I__1520\ : CascadeMux
    port map (
            O => \N__11139\,
            I => \N__11133\
        );

    \I__1519\ : CascadeMux
    port map (
            O => \N__11136\,
            I => \N__11130\
        );

    \I__1518\ : CascadeBuf
    port map (
            O => \N__11133\,
            I => \N__11127\
        );

    \I__1517\ : CascadeBuf
    port map (
            O => \N__11130\,
            I => \N__11124\
        );

    \I__1516\ : CascadeMux
    port map (
            O => \N__11127\,
            I => \N__11121\
        );

    \I__1515\ : CascadeMux
    port map (
            O => \N__11124\,
            I => \N__11118\
        );

    \I__1514\ : CascadeBuf
    port map (
            O => \N__11121\,
            I => \N__11115\
        );

    \I__1513\ : CascadeBuf
    port map (
            O => \N__11118\,
            I => \N__11112\
        );

    \I__1512\ : CascadeMux
    port map (
            O => \N__11115\,
            I => \N__11109\
        );

    \I__1511\ : CascadeMux
    port map (
            O => \N__11112\,
            I => \N__11106\
        );

    \I__1510\ : CascadeBuf
    port map (
            O => \N__11109\,
            I => \N__11103\
        );

    \I__1509\ : CascadeBuf
    port map (
            O => \N__11106\,
            I => \N__11100\
        );

    \I__1508\ : CascadeMux
    port map (
            O => \N__11103\,
            I => \N__11097\
        );

    \I__1507\ : CascadeMux
    port map (
            O => \N__11100\,
            I => \N__11094\
        );

    \I__1506\ : CascadeBuf
    port map (
            O => \N__11097\,
            I => \N__11091\
        );

    \I__1505\ : CascadeBuf
    port map (
            O => \N__11094\,
            I => \N__11088\
        );

    \I__1504\ : CascadeMux
    port map (
            O => \N__11091\,
            I => \N__11085\
        );

    \I__1503\ : CascadeMux
    port map (
            O => \N__11088\,
            I => \N__11082\
        );

    \I__1502\ : CascadeBuf
    port map (
            O => \N__11085\,
            I => \N__11079\
        );

    \I__1501\ : CascadeBuf
    port map (
            O => \N__11082\,
            I => \N__11076\
        );

    \I__1500\ : CascadeMux
    port map (
            O => \N__11079\,
            I => \N__11073\
        );

    \I__1499\ : CascadeMux
    port map (
            O => \N__11076\,
            I => \N__11070\
        );

    \I__1498\ : CascadeBuf
    port map (
            O => \N__11073\,
            I => \N__11067\
        );

    \I__1497\ : CascadeBuf
    port map (
            O => \N__11070\,
            I => \N__11064\
        );

    \I__1496\ : CascadeMux
    port map (
            O => \N__11067\,
            I => \N__11061\
        );

    \I__1495\ : CascadeMux
    port map (
            O => \N__11064\,
            I => \N__11058\
        );

    \I__1494\ : CascadeBuf
    port map (
            O => \N__11061\,
            I => \N__11055\
        );

    \I__1493\ : CascadeBuf
    port map (
            O => \N__11058\,
            I => \N__11052\
        );

    \I__1492\ : CascadeMux
    port map (
            O => \N__11055\,
            I => \N__11049\
        );

    \I__1491\ : CascadeMux
    port map (
            O => \N__11052\,
            I => \N__11046\
        );

    \I__1490\ : CascadeBuf
    port map (
            O => \N__11049\,
            I => \N__11043\
        );

    \I__1489\ : CascadeBuf
    port map (
            O => \N__11046\,
            I => \N__11040\
        );

    \I__1488\ : CascadeMux
    port map (
            O => \N__11043\,
            I => \N__11037\
        );

    \I__1487\ : CascadeMux
    port map (
            O => \N__11040\,
            I => \N__11034\
        );

    \I__1486\ : CascadeBuf
    port map (
            O => \N__11037\,
            I => \N__11031\
        );

    \I__1485\ : CascadeBuf
    port map (
            O => \N__11034\,
            I => \N__11028\
        );

    \I__1484\ : CascadeMux
    port map (
            O => \N__11031\,
            I => \N__11025\
        );

    \I__1483\ : CascadeMux
    port map (
            O => \N__11028\,
            I => \N__11022\
        );

    \I__1482\ : InMux
    port map (
            O => \N__11025\,
            I => \N__11019\
        );

    \I__1481\ : InMux
    port map (
            O => \N__11022\,
            I => \N__11016\
        );

    \I__1480\ : LocalMux
    port map (
            O => \N__11019\,
            I => \N__11013\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__11016\,
            I => \N__11010\
        );

    \I__1478\ : Span12Mux_v
    port map (
            O => \N__11013\,
            I => \N__11007\
        );

    \I__1477\ : Span12Mux_h
    port map (
            O => \N__11010\,
            I => \N__11004\
        );

    \I__1476\ : Span12Mux_h
    port map (
            O => \N__11007\,
            I => \N__10999\
        );

    \I__1475\ : Span12Mux_v
    port map (
            O => \N__11004\,
            I => \N__10999\
        );

    \I__1474\ : Odrv12
    port map (
            O => \N__10999\,
            I => \RX_ADDR_5\
        );

    \I__1473\ : InMux
    port map (
            O => \N__10996\,
            I => \receive_module.rx_counter.n3651\
        );

    \I__1472\ : InMux
    port map (
            O => \N__10993\,
            I => \N__10990\
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__10990\,
            I => \N__10987\
        );

    \I__1470\ : Span4Mux_v
    port map (
            O => \N__10987\,
            I => \N__10984\
        );

    \I__1469\ : Odrv4
    port map (
            O => \N__10984\,
            I => \transmit_module.Y_DELTA_PATTERN_81\
        );

    \I__1468\ : InMux
    port map (
            O => \N__10981\,
            I => \N__10978\
        );

    \I__1467\ : LocalMux
    port map (
            O => \N__10978\,
            I => \transmit_module.Y_DELTA_PATTERN_69\
        );

    \I__1466\ : InMux
    port map (
            O => \N__10975\,
            I => \N__10972\
        );

    \I__1465\ : LocalMux
    port map (
            O => \N__10972\,
            I => \transmit_module.Y_DELTA_PATTERN_68\
        );

    \I__1464\ : InMux
    port map (
            O => \N__10969\,
            I => \N__10966\
        );

    \I__1463\ : LocalMux
    port map (
            O => \N__10966\,
            I => \N__10963\
        );

    \I__1462\ : Odrv4
    port map (
            O => \N__10963\,
            I => \transmit_module.Y_DELTA_PATTERN_78\
        );

    \I__1461\ : InMux
    port map (
            O => \N__10960\,
            I => \N__10957\
        );

    \I__1460\ : LocalMux
    port map (
            O => \N__10957\,
            I => \transmit_module.Y_DELTA_PATTERN_62\
        );

    \I__1459\ : InMux
    port map (
            O => \N__10954\,
            I => \N__10951\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__10951\,
            I => \transmit_module.Y_DELTA_PATTERN_66\
        );

    \I__1457\ : InMux
    port map (
            O => \N__10948\,
            I => \N__10945\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__10945\,
            I => \transmit_module.Y_DELTA_PATTERN_65\
        );

    \I__1455\ : InMux
    port map (
            O => \N__10942\,
            I => \N__10939\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__10939\,
            I => \transmit_module.Y_DELTA_PATTERN_80\
        );

    \I__1453\ : InMux
    port map (
            O => \N__10936\,
            I => \N__10933\
        );

    \I__1452\ : LocalMux
    port map (
            O => \N__10933\,
            I => \transmit_module.Y_DELTA_PATTERN_79\
        );

    \I__1451\ : InMux
    port map (
            O => \N__10930\,
            I => \N__10927\
        );

    \I__1450\ : LocalMux
    port map (
            O => \N__10927\,
            I => \transmit_module.Y_DELTA_PATTERN_57\
        );

    \I__1449\ : CascadeMux
    port map (
            O => \N__10924\,
            I => \N__10919\
        );

    \I__1448\ : InMux
    port map (
            O => \N__10923\,
            I => \N__10916\
        );

    \I__1447\ : InMux
    port map (
            O => \N__10922\,
            I => \N__10913\
        );

    \I__1446\ : InMux
    port map (
            O => \N__10919\,
            I => \N__10910\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__10916\,
            I => \transmit_module.video_signal_controller.VGA_Y_11\
        );

    \I__1444\ : LocalMux
    port map (
            O => \N__10913\,
            I => \transmit_module.video_signal_controller.VGA_Y_11\
        );

    \I__1443\ : LocalMux
    port map (
            O => \N__10910\,
            I => \transmit_module.video_signal_controller.VGA_Y_11\
        );

    \I__1442\ : InMux
    port map (
            O => \N__10903\,
            I => \N__10898\
        );

    \I__1441\ : InMux
    port map (
            O => \N__10902\,
            I => \N__10895\
        );

    \I__1440\ : InMux
    port map (
            O => \N__10901\,
            I => \N__10892\
        );

    \I__1439\ : LocalMux
    port map (
            O => \N__10898\,
            I => \transmit_module.video_signal_controller.VGA_Y_10\
        );

    \I__1438\ : LocalMux
    port map (
            O => \N__10895\,
            I => \transmit_module.video_signal_controller.VGA_Y_10\
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__10892\,
            I => \transmit_module.video_signal_controller.VGA_Y_10\
        );

    \I__1436\ : InMux
    port map (
            O => \N__10885\,
            I => \N__10882\
        );

    \I__1435\ : LocalMux
    port map (
            O => \N__10882\,
            I => \transmit_module.video_signal_controller.n4218\
        );

    \I__1434\ : CascadeMux
    port map (
            O => \N__10879\,
            I => \transmit_module.n219_cascade_\
        );

    \I__1433\ : CascadeMux
    port map (
            O => \N__10876\,
            I => \N__10873\
        );

    \I__1432\ : CascadeBuf
    port map (
            O => \N__10873\,
            I => \N__10870\
        );

    \I__1431\ : CascadeMux
    port map (
            O => \N__10870\,
            I => \N__10866\
        );

    \I__1430\ : CascadeMux
    port map (
            O => \N__10869\,
            I => \N__10863\
        );

    \I__1429\ : CascadeBuf
    port map (
            O => \N__10866\,
            I => \N__10860\
        );

    \I__1428\ : CascadeBuf
    port map (
            O => \N__10863\,
            I => \N__10857\
        );

    \I__1427\ : CascadeMux
    port map (
            O => \N__10860\,
            I => \N__10854\
        );

    \I__1426\ : CascadeMux
    port map (
            O => \N__10857\,
            I => \N__10851\
        );

    \I__1425\ : CascadeBuf
    port map (
            O => \N__10854\,
            I => \N__10848\
        );

    \I__1424\ : CascadeBuf
    port map (
            O => \N__10851\,
            I => \N__10845\
        );

    \I__1423\ : CascadeMux
    port map (
            O => \N__10848\,
            I => \N__10842\
        );

    \I__1422\ : CascadeMux
    port map (
            O => \N__10845\,
            I => \N__10839\
        );

    \I__1421\ : CascadeBuf
    port map (
            O => \N__10842\,
            I => \N__10836\
        );

    \I__1420\ : CascadeBuf
    port map (
            O => \N__10839\,
            I => \N__10833\
        );

    \I__1419\ : CascadeMux
    port map (
            O => \N__10836\,
            I => \N__10830\
        );

    \I__1418\ : CascadeMux
    port map (
            O => \N__10833\,
            I => \N__10827\
        );

    \I__1417\ : CascadeBuf
    port map (
            O => \N__10830\,
            I => \N__10824\
        );

    \I__1416\ : CascadeBuf
    port map (
            O => \N__10827\,
            I => \N__10821\
        );

    \I__1415\ : CascadeMux
    port map (
            O => \N__10824\,
            I => \N__10818\
        );

    \I__1414\ : CascadeMux
    port map (
            O => \N__10821\,
            I => \N__10815\
        );

    \I__1413\ : CascadeBuf
    port map (
            O => \N__10818\,
            I => \N__10812\
        );

    \I__1412\ : CascadeBuf
    port map (
            O => \N__10815\,
            I => \N__10809\
        );

    \I__1411\ : CascadeMux
    port map (
            O => \N__10812\,
            I => \N__10806\
        );

    \I__1410\ : CascadeMux
    port map (
            O => \N__10809\,
            I => \N__10803\
        );

    \I__1409\ : CascadeBuf
    port map (
            O => \N__10806\,
            I => \N__10800\
        );

    \I__1408\ : CascadeBuf
    port map (
            O => \N__10803\,
            I => \N__10797\
        );

    \I__1407\ : CascadeMux
    port map (
            O => \N__10800\,
            I => \N__10794\
        );

    \I__1406\ : CascadeMux
    port map (
            O => \N__10797\,
            I => \N__10791\
        );

    \I__1405\ : CascadeBuf
    port map (
            O => \N__10794\,
            I => \N__10788\
        );

    \I__1404\ : CascadeBuf
    port map (
            O => \N__10791\,
            I => \N__10785\
        );

    \I__1403\ : CascadeMux
    port map (
            O => \N__10788\,
            I => \N__10782\
        );

    \I__1402\ : CascadeMux
    port map (
            O => \N__10785\,
            I => \N__10779\
        );

    \I__1401\ : CascadeBuf
    port map (
            O => \N__10782\,
            I => \N__10776\
        );

    \I__1400\ : CascadeBuf
    port map (
            O => \N__10779\,
            I => \N__10773\
        );

    \I__1399\ : CascadeMux
    port map (
            O => \N__10776\,
            I => \N__10770\
        );

    \I__1398\ : CascadeMux
    port map (
            O => \N__10773\,
            I => \N__10767\
        );

    \I__1397\ : CascadeBuf
    port map (
            O => \N__10770\,
            I => \N__10764\
        );

    \I__1396\ : CascadeBuf
    port map (
            O => \N__10767\,
            I => \N__10761\
        );

    \I__1395\ : CascadeMux
    port map (
            O => \N__10764\,
            I => \N__10758\
        );

    \I__1394\ : CascadeMux
    port map (
            O => \N__10761\,
            I => \N__10755\
        );

    \I__1393\ : CascadeBuf
    port map (
            O => \N__10758\,
            I => \N__10752\
        );

    \I__1392\ : CascadeBuf
    port map (
            O => \N__10755\,
            I => \N__10749\
        );

    \I__1391\ : CascadeMux
    port map (
            O => \N__10752\,
            I => \N__10746\
        );

    \I__1390\ : CascadeMux
    port map (
            O => \N__10749\,
            I => \N__10743\
        );

    \I__1389\ : CascadeBuf
    port map (
            O => \N__10746\,
            I => \N__10740\
        );

    \I__1388\ : CascadeBuf
    port map (
            O => \N__10743\,
            I => \N__10737\
        );

    \I__1387\ : CascadeMux
    port map (
            O => \N__10740\,
            I => \N__10734\
        );

    \I__1386\ : CascadeMux
    port map (
            O => \N__10737\,
            I => \N__10731\
        );

    \I__1385\ : CascadeBuf
    port map (
            O => \N__10734\,
            I => \N__10728\
        );

    \I__1384\ : CascadeBuf
    port map (
            O => \N__10731\,
            I => \N__10725\
        );

    \I__1383\ : CascadeMux
    port map (
            O => \N__10728\,
            I => \N__10722\
        );

    \I__1382\ : CascadeMux
    port map (
            O => \N__10725\,
            I => \N__10719\
        );

    \I__1381\ : CascadeBuf
    port map (
            O => \N__10722\,
            I => \N__10716\
        );

    \I__1380\ : CascadeBuf
    port map (
            O => \N__10719\,
            I => \N__10713\
        );

    \I__1379\ : CascadeMux
    port map (
            O => \N__10716\,
            I => \N__10710\
        );

    \I__1378\ : CascadeMux
    port map (
            O => \N__10713\,
            I => \N__10707\
        );

    \I__1377\ : CascadeBuf
    port map (
            O => \N__10710\,
            I => \N__10704\
        );

    \I__1376\ : CascadeBuf
    port map (
            O => \N__10707\,
            I => \N__10701\
        );

    \I__1375\ : CascadeMux
    port map (
            O => \N__10704\,
            I => \N__10698\
        );

    \I__1374\ : CascadeMux
    port map (
            O => \N__10701\,
            I => \N__10695\
        );

    \I__1373\ : InMux
    port map (
            O => \N__10698\,
            I => \N__10692\
        );

    \I__1372\ : CascadeBuf
    port map (
            O => \N__10695\,
            I => \N__10689\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__10692\,
            I => \N__10686\
        );

    \I__1370\ : CascadeMux
    port map (
            O => \N__10689\,
            I => \N__10683\
        );

    \I__1369\ : Span4Mux_h
    port map (
            O => \N__10686\,
            I => \N__10680\
        );

    \I__1368\ : InMux
    port map (
            O => \N__10683\,
            I => \N__10677\
        );

    \I__1367\ : Sp12to4
    port map (
            O => \N__10680\,
            I => \N__10674\
        );

    \I__1366\ : LocalMux
    port map (
            O => \N__10677\,
            I => \N__10671\
        );

    \I__1365\ : Span12Mux_v
    port map (
            O => \N__10674\,
            I => \N__10668\
        );

    \I__1364\ : Span4Mux_h
    port map (
            O => \N__10671\,
            I => \N__10665\
        );

    \I__1363\ : Span12Mux_h
    port map (
            O => \N__10668\,
            I => \N__10660\
        );

    \I__1362\ : Sp12to4
    port map (
            O => \N__10665\,
            I => \N__10660\
        );

    \I__1361\ : Odrv12
    port map (
            O => \N__10660\,
            I => n28
        );

    \I__1360\ : IoInMux
    port map (
            O => \N__10657\,
            I => \N__10654\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__10654\,
            I => \N__10651\
        );

    \I__1358\ : IoSpan4Mux
    port map (
            O => \N__10651\,
            I => \N__10648\
        );

    \I__1357\ : Span4Mux_s2_h
    port map (
            O => \N__10648\,
            I => \N__10645\
        );

    \I__1356\ : Sp12to4
    port map (
            O => \N__10645\,
            I => \N__10642\
        );

    \I__1355\ : Odrv12
    port map (
            O => \N__10642\,
            I => n4210
        );

    \I__1354\ : CascadeMux
    port map (
            O => \N__10639\,
            I => \n4210_cascade_\
        );

    \I__1353\ : InMux
    port map (
            O => \N__10636\,
            I => \N__10633\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__10633\,
            I => \transmit_module.Y_DELTA_PATTERN_64\
        );

    \I__1351\ : InMux
    port map (
            O => \N__10630\,
            I => \N__10627\
        );

    \I__1350\ : LocalMux
    port map (
            O => \N__10627\,
            I => \transmit_module.Y_DELTA_PATTERN_67\
        );

    \I__1349\ : InMux
    port map (
            O => \N__10624\,
            I => \N__10620\
        );

    \I__1348\ : InMux
    port map (
            O => \N__10623\,
            I => \N__10617\
        );

    \I__1347\ : LocalMux
    port map (
            O => \N__10620\,
            I => \transmit_module.video_signal_controller.VGA_Y_7\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__10617\,
            I => \transmit_module.video_signal_controller.VGA_Y_7\
        );

    \I__1345\ : InMux
    port map (
            O => \N__10612\,
            I => \transmit_module.video_signal_controller.n3683\
        );

    \I__1344\ : InMux
    port map (
            O => \N__10609\,
            I => \N__10605\
        );

    \I__1343\ : InMux
    port map (
            O => \N__10608\,
            I => \N__10602\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__10605\,
            I => \transmit_module.video_signal_controller.VGA_Y_8\
        );

    \I__1341\ : LocalMux
    port map (
            O => \N__10602\,
            I => \transmit_module.video_signal_controller.VGA_Y_8\
        );

    \I__1340\ : InMux
    port map (
            O => \N__10597\,
            I => \bfn_12_17_0_\
        );

    \I__1339\ : InMux
    port map (
            O => \N__10594\,
            I => \transmit_module.video_signal_controller.n3685\
        );

    \I__1338\ : InMux
    port map (
            O => \N__10591\,
            I => \transmit_module.video_signal_controller.n3686\
        );

    \I__1337\ : InMux
    port map (
            O => \N__10588\,
            I => \transmit_module.video_signal_controller.n3687\
        );

    \I__1336\ : SRMux
    port map (
            O => \N__10585\,
            I => \N__10581\
        );

    \I__1335\ : SRMux
    port map (
            O => \N__10584\,
            I => \N__10578\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__10581\,
            I => \N__10575\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__10578\,
            I => \N__10572\
        );

    \I__1332\ : Span4Mux_h
    port map (
            O => \N__10575\,
            I => \N__10569\
        );

    \I__1331\ : Span4Mux_v
    port map (
            O => \N__10572\,
            I => \N__10566\
        );

    \I__1330\ : Odrv4
    port map (
            O => \N__10569\,
            I => \transmit_module.video_signal_controller.n2594\
        );

    \I__1329\ : Odrv4
    port map (
            O => \N__10566\,
            I => \transmit_module.video_signal_controller.n2594\
        );

    \I__1328\ : InMux
    port map (
            O => \N__10561\,
            I => \N__10556\
        );

    \I__1327\ : InMux
    port map (
            O => \N__10560\,
            I => \N__10552\
        );

    \I__1326\ : InMux
    port map (
            O => \N__10559\,
            I => \N__10549\
        );

    \I__1325\ : LocalMux
    port map (
            O => \N__10556\,
            I => \N__10546\
        );

    \I__1324\ : InMux
    port map (
            O => \N__10555\,
            I => \N__10543\
        );

    \I__1323\ : LocalMux
    port map (
            O => \N__10552\,
            I => \transmit_module.video_signal_controller.VGA_Y_3\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__10549\,
            I => \transmit_module.video_signal_controller.VGA_Y_3\
        );

    \I__1321\ : Odrv4
    port map (
            O => \N__10546\,
            I => \transmit_module.video_signal_controller.VGA_Y_3\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__10543\,
            I => \transmit_module.video_signal_controller.VGA_Y_3\
        );

    \I__1319\ : InMux
    port map (
            O => \N__10534\,
            I => \N__10531\
        );

    \I__1318\ : LocalMux
    port map (
            O => \N__10531\,
            I => \transmit_module.video_signal_controller.n4215\
        );

    \I__1317\ : CascadeMux
    port map (
            O => \N__10528\,
            I => \N__10524\
        );

    \I__1316\ : CascadeMux
    port map (
            O => \N__10527\,
            I => \N__10521\
        );

    \I__1315\ : InMux
    port map (
            O => \N__10524\,
            I => \N__10517\
        );

    \I__1314\ : InMux
    port map (
            O => \N__10521\,
            I => \N__10513\
        );

    \I__1313\ : InMux
    port map (
            O => \N__10520\,
            I => \N__10510\
        );

    \I__1312\ : LocalMux
    port map (
            O => \N__10517\,
            I => \N__10507\
        );

    \I__1311\ : InMux
    port map (
            O => \N__10516\,
            I => \N__10504\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__10513\,
            I => \transmit_module.video_signal_controller.VGA_Y_4\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__10510\,
            I => \transmit_module.video_signal_controller.VGA_Y_4\
        );

    \I__1308\ : Odrv4
    port map (
            O => \N__10507\,
            I => \transmit_module.video_signal_controller.VGA_Y_4\
        );

    \I__1307\ : LocalMux
    port map (
            O => \N__10504\,
            I => \transmit_module.video_signal_controller.VGA_Y_4\
        );

    \I__1306\ : InMux
    port map (
            O => \N__10495\,
            I => \N__10491\
        );

    \I__1305\ : InMux
    port map (
            O => \N__10494\,
            I => \N__10488\
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__10491\,
            I => \transmit_module.video_signal_controller.n3892\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__10488\,
            I => \transmit_module.video_signal_controller.n3892\
        );

    \I__1302\ : InMux
    port map (
            O => \N__10483\,
            I => \N__10478\
        );

    \I__1301\ : InMux
    port map (
            O => \N__10482\,
            I => \N__10475\
        );

    \I__1300\ : InMux
    port map (
            O => \N__10481\,
            I => \N__10472\
        );

    \I__1299\ : LocalMux
    port map (
            O => \N__10478\,
            I => \transmit_module.video_signal_controller.VGA_Y_9\
        );

    \I__1298\ : LocalMux
    port map (
            O => \N__10475\,
            I => \transmit_module.video_signal_controller.VGA_Y_9\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__10472\,
            I => \transmit_module.video_signal_controller.VGA_Y_9\
        );

    \I__1296\ : CascadeMux
    port map (
            O => \N__10465\,
            I => \transmit_module.video_signal_controller.VGA_VISIBLE_Y_N_553_cascade_\
        );

    \I__1295\ : InMux
    port map (
            O => \N__10462\,
            I => \N__10459\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__10459\,
            I => \transmit_module.video_signal_controller.n3936\
        );

    \I__1293\ : CascadeMux
    port map (
            O => \N__10456\,
            I => \transmit_module.n3926_cascade_\
        );

    \I__1292\ : CascadeMux
    port map (
            O => \N__10453\,
            I => \transmit_module.video_signal_controller.n18_cascade_\
        );

    \I__1291\ : InMux
    port map (
            O => \N__10450\,
            I => \N__10447\
        );

    \I__1290\ : LocalMux
    port map (
            O => \N__10447\,
            I => \transmit_module.video_signal_controller.n2219\
        );

    \I__1289\ : InMux
    port map (
            O => \N__10444\,
            I => \N__10440\
        );

    \I__1288\ : InMux
    port map (
            O => \N__10443\,
            I => \N__10437\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__10440\,
            I => \transmit_module.video_signal_controller.VGA_Y_0\
        );

    \I__1286\ : LocalMux
    port map (
            O => \N__10437\,
            I => \transmit_module.video_signal_controller.VGA_Y_0\
        );

    \I__1285\ : InMux
    port map (
            O => \N__10432\,
            I => \bfn_12_16_0_\
        );

    \I__1284\ : CascadeMux
    port map (
            O => \N__10429\,
            I => \N__10424\
        );

    \I__1283\ : InMux
    port map (
            O => \N__10428\,
            I => \N__10420\
        );

    \I__1282\ : InMux
    port map (
            O => \N__10427\,
            I => \N__10417\
        );

    \I__1281\ : InMux
    port map (
            O => \N__10424\,
            I => \N__10412\
        );

    \I__1280\ : InMux
    port map (
            O => \N__10423\,
            I => \N__10412\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__10420\,
            I => \transmit_module.video_signal_controller.VGA_Y_1\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__10417\,
            I => \transmit_module.video_signal_controller.VGA_Y_1\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__10412\,
            I => \transmit_module.video_signal_controller.VGA_Y_1\
        );

    \I__1276\ : InMux
    port map (
            O => \N__10405\,
            I => \transmit_module.video_signal_controller.n3677\
        );

    \I__1275\ : InMux
    port map (
            O => \N__10402\,
            I => \N__10396\
        );

    \I__1274\ : InMux
    port map (
            O => \N__10401\,
            I => \N__10393\
        );

    \I__1273\ : InMux
    port map (
            O => \N__10400\,
            I => \N__10388\
        );

    \I__1272\ : InMux
    port map (
            O => \N__10399\,
            I => \N__10388\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__10396\,
            I => \transmit_module.video_signal_controller.VGA_Y_2\
        );

    \I__1270\ : LocalMux
    port map (
            O => \N__10393\,
            I => \transmit_module.video_signal_controller.VGA_Y_2\
        );

    \I__1269\ : LocalMux
    port map (
            O => \N__10388\,
            I => \transmit_module.video_signal_controller.VGA_Y_2\
        );

    \I__1268\ : InMux
    port map (
            O => \N__10381\,
            I => \transmit_module.video_signal_controller.n3678\
        );

    \I__1267\ : InMux
    port map (
            O => \N__10378\,
            I => \transmit_module.video_signal_controller.n3679\
        );

    \I__1266\ : InMux
    port map (
            O => \N__10375\,
            I => \transmit_module.video_signal_controller.n3680\
        );

    \I__1265\ : InMux
    port map (
            O => \N__10372\,
            I => \N__10367\
        );

    \I__1264\ : InMux
    port map (
            O => \N__10371\,
            I => \N__10364\
        );

    \I__1263\ : InMux
    port map (
            O => \N__10370\,
            I => \N__10361\
        );

    \I__1262\ : LocalMux
    port map (
            O => \N__10367\,
            I => \transmit_module.video_signal_controller.VGA_Y_5\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__10364\,
            I => \transmit_module.video_signal_controller.VGA_Y_5\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__10361\,
            I => \transmit_module.video_signal_controller.VGA_Y_5\
        );

    \I__1259\ : InMux
    port map (
            O => \N__10354\,
            I => \transmit_module.video_signal_controller.n3681\
        );

    \I__1258\ : InMux
    port map (
            O => \N__10351\,
            I => \N__10346\
        );

    \I__1257\ : InMux
    port map (
            O => \N__10350\,
            I => \N__10341\
        );

    \I__1256\ : InMux
    port map (
            O => \N__10349\,
            I => \N__10341\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__10346\,
            I => \transmit_module.video_signal_controller.VGA_Y_6\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__10341\,
            I => \transmit_module.video_signal_controller.VGA_Y_6\
        );

    \I__1253\ : InMux
    port map (
            O => \N__10336\,
            I => \transmit_module.video_signal_controller.n3682\
        );

    \I__1252\ : InMux
    port map (
            O => \N__10333\,
            I => \N__10330\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__10330\,
            I => \transmit_module.video_signal_controller.n4052\
        );

    \I__1250\ : CascadeMux
    port map (
            O => \N__10327\,
            I => \transmit_module.video_signal_controller.n4216_cascade_\
        );

    \I__1249\ : InMux
    port map (
            O => \N__10324\,
            I => \N__10321\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__10321\,
            I => \transmit_module.video_signal_controller.n12\
        );

    \I__1247\ : CascadeMux
    port map (
            O => \N__10318\,
            I => \transmit_module.video_signal_controller.n2274_cascade_\
        );

    \I__1246\ : InMux
    port map (
            O => \N__10315\,
            I => \N__10312\
        );

    \I__1245\ : LocalMux
    port map (
            O => \N__10312\,
            I => \transmit_module.video_signal_controller.SYNC_BUFF2\
        );

    \I__1244\ : CascadeMux
    port map (
            O => \N__10309\,
            I => \N__10306\
        );

    \I__1243\ : InMux
    port map (
            O => \N__10306\,
            I => \N__10303\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__10303\,
            I => \transmit_module.video_signal_controller.n3226\
        );

    \I__1241\ : CascadeMux
    port map (
            O => \N__10300\,
            I => \N__10297\
        );

    \I__1240\ : InMux
    port map (
            O => \N__10297\,
            I => \N__10294\
        );

    \I__1239\ : LocalMux
    port map (
            O => \N__10294\,
            I => \transmit_module.video_signal_controller.n2260\
        );

    \I__1238\ : InMux
    port map (
            O => \N__10291\,
            I => \N__10285\
        );

    \I__1237\ : InMux
    port map (
            O => \N__10290\,
            I => \N__10285\
        );

    \I__1236\ : LocalMux
    port map (
            O => \N__10285\,
            I => \transmit_module.video_signal_controller.n3917\
        );

    \I__1235\ : CascadeMux
    port map (
            O => \N__10282\,
            I => \transmit_module.video_signal_controller.n2260_cascade_\
        );

    \I__1234\ : InMux
    port map (
            O => \N__10279\,
            I => \N__10276\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__10276\,
            I => \transmit_module.video_signal_controller.n4217\
        );

    \I__1232\ : SRMux
    port map (
            O => \N__10273\,
            I => \N__10270\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__10270\,
            I => \N__10266\
        );

    \I__1230\ : SRMux
    port map (
            O => \N__10269\,
            I => \N__10263\
        );

    \I__1229\ : Span4Mux_v
    port map (
            O => \N__10266\,
            I => \N__10257\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__10263\,
            I => \N__10257\
        );

    \I__1227\ : SRMux
    port map (
            O => \N__10262\,
            I => \N__10254\
        );

    \I__1226\ : Span4Mux_v
    port map (
            O => \N__10257\,
            I => \N__10248\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__10254\,
            I => \N__10248\
        );

    \I__1224\ : SRMux
    port map (
            O => \N__10253\,
            I => \N__10245\
        );

    \I__1223\ : Span4Mux_v
    port map (
            O => \N__10248\,
            I => \N__10240\
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__10245\,
            I => \N__10240\
        );

    \I__1221\ : Span4Mux_h
    port map (
            O => \N__10240\,
            I => \N__10237\
        );

    \I__1220\ : Odrv4
    port map (
            O => \N__10237\,
            I => n691
        );

    \I__1219\ : SRMux
    port map (
            O => \N__10234\,
            I => \N__10231\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__10231\,
            I => \N__10228\
        );

    \I__1217\ : Span4Mux_s2_v
    port map (
            O => \N__10228\,
            I => \N__10222\
        );

    \I__1216\ : SRMux
    port map (
            O => \N__10227\,
            I => \N__10219\
        );

    \I__1215\ : SRMux
    port map (
            O => \N__10226\,
            I => \N__10216\
        );

    \I__1214\ : SRMux
    port map (
            O => \N__10225\,
            I => \N__10213\
        );

    \I__1213\ : Span4Mux_v
    port map (
            O => \N__10222\,
            I => \N__10206\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__10219\,
            I => \N__10206\
        );

    \I__1211\ : LocalMux
    port map (
            O => \N__10216\,
            I => \N__10206\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__10213\,
            I => \N__10203\
        );

    \I__1209\ : Span4Mux_v
    port map (
            O => \N__10206\,
            I => \N__10198\
        );

    \I__1208\ : Span4Mux_v
    port map (
            O => \N__10203\,
            I => \N__10198\
        );

    \I__1207\ : Span4Mux_h
    port map (
            O => \N__10198\,
            I => \N__10195\
        );

    \I__1206\ : Sp12to4
    port map (
            O => \N__10195\,
            I => \N__10192\
        );

    \I__1205\ : Odrv12
    port map (
            O => \N__10192\,
            I => \line_buffer.n626\
        );

    \I__1204\ : SRMux
    port map (
            O => \N__10189\,
            I => \N__10185\
        );

    \I__1203\ : SRMux
    port map (
            O => \N__10188\,
            I => \N__10182\
        );

    \I__1202\ : LocalMux
    port map (
            O => \N__10185\,
            I => \N__10175\
        );

    \I__1201\ : LocalMux
    port map (
            O => \N__10182\,
            I => \N__10175\
        );

    \I__1200\ : SRMux
    port map (
            O => \N__10181\,
            I => \N__10172\
        );

    \I__1199\ : SRMux
    port map (
            O => \N__10180\,
            I => \N__10169\
        );

    \I__1198\ : Span4Mux_v
    port map (
            O => \N__10175\,
            I => \N__10164\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__10172\,
            I => \N__10164\
        );

    \I__1196\ : LocalMux
    port map (
            O => \N__10169\,
            I => \N__10161\
        );

    \I__1195\ : Span4Mux_v
    port map (
            O => \N__10164\,
            I => \N__10158\
        );

    \I__1194\ : Span4Mux_h
    port map (
            O => \N__10161\,
            I => \N__10155\
        );

    \I__1193\ : Span4Mux_v
    port map (
            O => \N__10158\,
            I => \N__10152\
        );

    \I__1192\ : Sp12to4
    port map (
            O => \N__10155\,
            I => \N__10149\
        );

    \I__1191\ : Span4Mux_v
    port map (
            O => \N__10152\,
            I => \N__10146\
        );

    \I__1190\ : Span12Mux_h
    port map (
            O => \N__10149\,
            I => \N__10143\
        );

    \I__1189\ : Span4Mux_v
    port map (
            O => \N__10146\,
            I => \N__10140\
        );

    \I__1188\ : Odrv12
    port map (
            O => \N__10143\,
            I => \line_buffer.n561\
        );

    \I__1187\ : Odrv4
    port map (
            O => \N__10140\,
            I => \line_buffer.n561\
        );

    \I__1186\ : CascadeMux
    port map (
            O => \N__10135\,
            I => \transmit_module.video_signal_controller.n3978_cascade_\
        );

    \I__1185\ : CascadeMux
    port map (
            O => \N__10132\,
            I => \receive_module.n4212_cascade_\
        );

    \I__1184\ : CascadeMux
    port map (
            O => \N__10129\,
            I => \receive_module.n4213_cascade_\
        );

    \I__1183\ : InMux
    port map (
            O => \N__10126\,
            I => \N__10123\
        );

    \I__1182\ : LocalMux
    port map (
            O => \N__10123\,
            I => \receive_module.rx_counter.n3204\
        );

    \I__1181\ : SRMux
    port map (
            O => \N__10120\,
            I => \N__10117\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__10117\,
            I => \N__10114\
        );

    \I__1179\ : Span4Mux_v
    port map (
            O => \N__10114\,
            I => \N__10109\
        );

    \I__1178\ : SRMux
    port map (
            O => \N__10113\,
            I => \N__10106\
        );

    \I__1177\ : SRMux
    port map (
            O => \N__10112\,
            I => \N__10102\
        );

    \I__1176\ : Span4Mux_v
    port map (
            O => \N__10109\,
            I => \N__10099\
        );

    \I__1175\ : LocalMux
    port map (
            O => \N__10106\,
            I => \N__10096\
        );

    \I__1174\ : SRMux
    port map (
            O => \N__10105\,
            I => \N__10093\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__10102\,
            I => \N__10090\
        );

    \I__1172\ : Span4Mux_v
    port map (
            O => \N__10099\,
            I => \N__10083\
        );

    \I__1171\ : Span4Mux_v
    port map (
            O => \N__10096\,
            I => \N__10083\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__10093\,
            I => \N__10083\
        );

    \I__1169\ : Span4Mux_h
    port map (
            O => \N__10090\,
            I => \N__10078\
        );

    \I__1168\ : Span4Mux_h
    port map (
            O => \N__10083\,
            I => \N__10078\
        );

    \I__1167\ : Odrv4
    port map (
            O => \N__10078\,
            I => n659
        );

    \I__1166\ : IoInMux
    port map (
            O => \N__10075\,
            I => \N__10072\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__10072\,
            I => \N__10069\
        );

    \I__1164\ : Span4Mux_s3_h
    port map (
            O => \N__10069\,
            I => \N__10066\
        );

    \I__1163\ : Span4Mux_v
    port map (
            O => \N__10066\,
            I => \N__10063\
        );

    \I__1162\ : Span4Mux_h
    port map (
            O => \N__10063\,
            I => \N__10060\
        );

    \I__1161\ : Span4Mux_h
    port map (
            O => \N__10060\,
            I => \N__10057\
        );

    \I__1160\ : Odrv4
    port map (
            O => \N__10057\,
            I => \DEBUG_c_0\
        );

    \I__1159\ : IoInMux
    port map (
            O => \N__10054\,
            I => \N__10051\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__10051\,
            I => \N__10048\
        );

    \I__1157\ : IoSpan4Mux
    port map (
            O => \N__10048\,
            I => \N__10044\
        );

    \I__1156\ : IoInMux
    port map (
            O => \N__10047\,
            I => \N__10041\
        );

    \I__1155\ : Span4Mux_s1_v
    port map (
            O => \N__10044\,
            I => \N__10037\
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__10041\,
            I => \N__10034\
        );

    \I__1153\ : IoInMux
    port map (
            O => \N__10040\,
            I => \N__10031\
        );

    \I__1152\ : Span4Mux_v
    port map (
            O => \N__10037\,
            I => \N__10026\
        );

    \I__1151\ : Span4Mux_s2_h
    port map (
            O => \N__10034\,
            I => \N__10026\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__10031\,
            I => \N__10023\
        );

    \I__1149\ : Span4Mux_h
    port map (
            O => \N__10026\,
            I => \N__10020\
        );

    \I__1148\ : Span4Mux_s1_v
    port map (
            O => \N__10023\,
            I => \N__10017\
        );

    \I__1147\ : Span4Mux_h
    port map (
            O => \N__10020\,
            I => \N__10012\
        );

    \I__1146\ : Span4Mux_v
    port map (
            O => \N__10017\,
            I => \N__10012\
        );

    \I__1145\ : Span4Mux_v
    port map (
            O => \N__10012\,
            I => \N__10009\
        );

    \I__1144\ : Odrv4
    port map (
            O => \N__10009\,
            I => n1996
        );

    \I__1143\ : InMux
    port map (
            O => \N__10006\,
            I => \N__10003\
        );

    \I__1142\ : LocalMux
    port map (
            O => \N__10003\,
            I => \transmit_module.Y_DELTA_PATTERN_70\
        );

    \I__1141\ : InMux
    port map (
            O => \N__10000\,
            I => \N__9997\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__9997\,
            I => \N__9994\
        );

    \I__1139\ : Odrv4
    port map (
            O => \N__9994\,
            I => \transmit_module.Y_DELTA_PATTERN_72\
        );

    \I__1138\ : InMux
    port map (
            O => \N__9991\,
            I => \N__9988\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__9988\,
            I => \transmit_module.Y_DELTA_PATTERN_71\
        );

    \I__1136\ : InMux
    port map (
            O => \N__9985\,
            I => \N__9982\
        );

    \I__1135\ : LocalMux
    port map (
            O => \N__9982\,
            I => \transmit_module.Y_DELTA_PATTERN_63\
        );

    \I__1134\ : CascadeMux
    port map (
            O => \N__9979\,
            I => \N__9976\
        );

    \I__1133\ : CascadeBuf
    port map (
            O => \N__9976\,
            I => \N__9972\
        );

    \I__1132\ : CascadeMux
    port map (
            O => \N__9975\,
            I => \N__9969\
        );

    \I__1131\ : CascadeMux
    port map (
            O => \N__9972\,
            I => \N__9966\
        );

    \I__1130\ : CascadeBuf
    port map (
            O => \N__9969\,
            I => \N__9963\
        );

    \I__1129\ : CascadeBuf
    port map (
            O => \N__9966\,
            I => \N__9960\
        );

    \I__1128\ : CascadeMux
    port map (
            O => \N__9963\,
            I => \N__9957\
        );

    \I__1127\ : CascadeMux
    port map (
            O => \N__9960\,
            I => \N__9954\
        );

    \I__1126\ : CascadeBuf
    port map (
            O => \N__9957\,
            I => \N__9951\
        );

    \I__1125\ : CascadeBuf
    port map (
            O => \N__9954\,
            I => \N__9948\
        );

    \I__1124\ : CascadeMux
    port map (
            O => \N__9951\,
            I => \N__9945\
        );

    \I__1123\ : CascadeMux
    port map (
            O => \N__9948\,
            I => \N__9942\
        );

    \I__1122\ : CascadeBuf
    port map (
            O => \N__9945\,
            I => \N__9939\
        );

    \I__1121\ : CascadeBuf
    port map (
            O => \N__9942\,
            I => \N__9936\
        );

    \I__1120\ : CascadeMux
    port map (
            O => \N__9939\,
            I => \N__9933\
        );

    \I__1119\ : CascadeMux
    port map (
            O => \N__9936\,
            I => \N__9930\
        );

    \I__1118\ : CascadeBuf
    port map (
            O => \N__9933\,
            I => \N__9927\
        );

    \I__1117\ : CascadeBuf
    port map (
            O => \N__9930\,
            I => \N__9924\
        );

    \I__1116\ : CascadeMux
    port map (
            O => \N__9927\,
            I => \N__9921\
        );

    \I__1115\ : CascadeMux
    port map (
            O => \N__9924\,
            I => \N__9918\
        );

    \I__1114\ : CascadeBuf
    port map (
            O => \N__9921\,
            I => \N__9915\
        );

    \I__1113\ : CascadeBuf
    port map (
            O => \N__9918\,
            I => \N__9912\
        );

    \I__1112\ : CascadeMux
    port map (
            O => \N__9915\,
            I => \N__9909\
        );

    \I__1111\ : CascadeMux
    port map (
            O => \N__9912\,
            I => \N__9906\
        );

    \I__1110\ : CascadeBuf
    port map (
            O => \N__9909\,
            I => \N__9903\
        );

    \I__1109\ : CascadeBuf
    port map (
            O => \N__9906\,
            I => \N__9900\
        );

    \I__1108\ : CascadeMux
    port map (
            O => \N__9903\,
            I => \N__9897\
        );

    \I__1107\ : CascadeMux
    port map (
            O => \N__9900\,
            I => \N__9894\
        );

    \I__1106\ : CascadeBuf
    port map (
            O => \N__9897\,
            I => \N__9891\
        );

    \I__1105\ : CascadeBuf
    port map (
            O => \N__9894\,
            I => \N__9888\
        );

    \I__1104\ : CascadeMux
    port map (
            O => \N__9891\,
            I => \N__9885\
        );

    \I__1103\ : CascadeMux
    port map (
            O => \N__9888\,
            I => \N__9882\
        );

    \I__1102\ : CascadeBuf
    port map (
            O => \N__9885\,
            I => \N__9879\
        );

    \I__1101\ : CascadeBuf
    port map (
            O => \N__9882\,
            I => \N__9876\
        );

    \I__1100\ : CascadeMux
    port map (
            O => \N__9879\,
            I => \N__9873\
        );

    \I__1099\ : CascadeMux
    port map (
            O => \N__9876\,
            I => \N__9870\
        );

    \I__1098\ : CascadeBuf
    port map (
            O => \N__9873\,
            I => \N__9867\
        );

    \I__1097\ : CascadeBuf
    port map (
            O => \N__9870\,
            I => \N__9864\
        );

    \I__1096\ : CascadeMux
    port map (
            O => \N__9867\,
            I => \N__9861\
        );

    \I__1095\ : CascadeMux
    port map (
            O => \N__9864\,
            I => \N__9858\
        );

    \I__1094\ : CascadeBuf
    port map (
            O => \N__9861\,
            I => \N__9855\
        );

    \I__1093\ : CascadeBuf
    port map (
            O => \N__9858\,
            I => \N__9852\
        );

    \I__1092\ : CascadeMux
    port map (
            O => \N__9855\,
            I => \N__9849\
        );

    \I__1091\ : CascadeMux
    port map (
            O => \N__9852\,
            I => \N__9846\
        );

    \I__1090\ : CascadeBuf
    port map (
            O => \N__9849\,
            I => \N__9843\
        );

    \I__1089\ : CascadeBuf
    port map (
            O => \N__9846\,
            I => \N__9840\
        );

    \I__1088\ : CascadeMux
    port map (
            O => \N__9843\,
            I => \N__9837\
        );

    \I__1087\ : CascadeMux
    port map (
            O => \N__9840\,
            I => \N__9834\
        );

    \I__1086\ : CascadeBuf
    port map (
            O => \N__9837\,
            I => \N__9831\
        );

    \I__1085\ : CascadeBuf
    port map (
            O => \N__9834\,
            I => \N__9828\
        );

    \I__1084\ : CascadeMux
    port map (
            O => \N__9831\,
            I => \N__9825\
        );

    \I__1083\ : CascadeMux
    port map (
            O => \N__9828\,
            I => \N__9822\
        );

    \I__1082\ : CascadeBuf
    port map (
            O => \N__9825\,
            I => \N__9819\
        );

    \I__1081\ : CascadeBuf
    port map (
            O => \N__9822\,
            I => \N__9816\
        );

    \I__1080\ : CascadeMux
    port map (
            O => \N__9819\,
            I => \N__9813\
        );

    \I__1079\ : CascadeMux
    port map (
            O => \N__9816\,
            I => \N__9810\
        );

    \I__1078\ : CascadeBuf
    port map (
            O => \N__9813\,
            I => \N__9807\
        );

    \I__1077\ : CascadeBuf
    port map (
            O => \N__9810\,
            I => \N__9804\
        );

    \I__1076\ : CascadeMux
    port map (
            O => \N__9807\,
            I => \N__9801\
        );

    \I__1075\ : CascadeMux
    port map (
            O => \N__9804\,
            I => \N__9798\
        );

    \I__1074\ : CascadeBuf
    port map (
            O => \N__9801\,
            I => \N__9795\
        );

    \I__1073\ : InMux
    port map (
            O => \N__9798\,
            I => \N__9792\
        );

    \I__1072\ : CascadeMux
    port map (
            O => \N__9795\,
            I => \N__9789\
        );

    \I__1071\ : LocalMux
    port map (
            O => \N__9792\,
            I => \N__9786\
        );

    \I__1070\ : InMux
    port map (
            O => \N__9789\,
            I => \N__9783\
        );

    \I__1069\ : Span12Mux_h
    port map (
            O => \N__9786\,
            I => \N__9780\
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__9783\,
            I => \N__9777\
        );

    \I__1067\ : Odrv12
    port map (
            O => \N__9780\,
            I => n18
        );

    \I__1066\ : Odrv4
    port map (
            O => \N__9777\,
            I => n18
        );

    \I__1065\ : SRMux
    port map (
            O => \N__9772\,
            I => \N__9769\
        );

    \I__1064\ : LocalMux
    port map (
            O => \N__9769\,
            I => \N__9765\
        );

    \I__1063\ : SRMux
    port map (
            O => \N__9768\,
            I => \N__9762\
        );

    \I__1062\ : Span4Mux_v
    port map (
            O => \N__9765\,
            I => \N__9757\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__9762\,
            I => \N__9757\
        );

    \I__1060\ : Span4Mux_h
    port map (
            O => \N__9757\,
            I => \N__9754\
        );

    \I__1059\ : Sp12to4
    port map (
            O => \N__9754\,
            I => \N__9751\
        );

    \I__1058\ : Odrv12
    port map (
            O => \N__9751\,
            I => \receive_module.rx_counter.PULSE_1HZ_N_97\
        );

    \I__1057\ : CascadeMux
    port map (
            O => \N__9748\,
            I => \transmit_module.video_signal_controller.n3935_cascade_\
        );

    \I__1056\ : InMux
    port map (
            O => \N__9745\,
            I => \N__9742\
        );

    \I__1055\ : LocalMux
    port map (
            O => \N__9742\,
            I => \transmit_module.video_signal_controller.n6\
        );

    \I__1054\ : InMux
    port map (
            O => \N__9739\,
            I => \N__9736\
        );

    \I__1053\ : LocalMux
    port map (
            O => \N__9736\,
            I => \transmit_module.Y_DELTA_PATTERN_98\
        );

    \I__1052\ : InMux
    port map (
            O => \N__9733\,
            I => \N__9730\
        );

    \I__1051\ : LocalMux
    port map (
            O => \N__9730\,
            I => \transmit_module.Y_DELTA_PATTERN_76\
        );

    \I__1050\ : InMux
    port map (
            O => \N__9727\,
            I => \N__9724\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__9724\,
            I => \transmit_module.Y_DELTA_PATTERN_73\
        );

    \I__1048\ : InMux
    port map (
            O => \N__9721\,
            I => \N__9718\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__9718\,
            I => \N__9715\
        );

    \I__1046\ : Span4Mux_v
    port map (
            O => \N__9715\,
            I => \N__9712\
        );

    \I__1045\ : Odrv4
    port map (
            O => \N__9712\,
            I => \transmit_module.Y_DELTA_PATTERN_82\
        );

    \I__1044\ : InMux
    port map (
            O => \N__9709\,
            I => \N__9706\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__9706\,
            I => \transmit_module.Y_DELTA_PATTERN_75\
        );

    \I__1042\ : InMux
    port map (
            O => \N__9703\,
            I => \N__9700\
        );

    \I__1041\ : LocalMux
    port map (
            O => \N__9700\,
            I => \transmit_module.Y_DELTA_PATTERN_74\
        );

    \I__1040\ : InMux
    port map (
            O => \N__9697\,
            I => \N__9694\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__9694\,
            I => \transmit_module.Y_DELTA_PATTERN_77\
        );

    \I__1038\ : CascadeMux
    port map (
            O => \N__9691\,
            I => \N__9688\
        );

    \I__1037\ : InMux
    port map (
            O => \N__9688\,
            I => \N__9685\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__9685\,
            I => \N__9682\
        );

    \I__1035\ : Odrv4
    port map (
            O => \N__9682\,
            I => \receive_module.rx_counter.n3979\
        );

    \I__1034\ : InMux
    port map (
            O => \N__9679\,
            I => \receive_module.rx_counter.O_VISIBLE_N_89\
        );

    \I__1033\ : IoInMux
    port map (
            O => \N__9676\,
            I => \N__9673\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__9673\,
            I => \N__9669\
        );

    \I__1031\ : InMux
    port map (
            O => \N__9672\,
            I => \N__9666\
        );

    \I__1030\ : Span4Mux_s1_h
    port map (
            O => \N__9669\,
            I => \N__9663\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__9666\,
            I => \N__9660\
        );

    \I__1028\ : Sp12to4
    port map (
            O => \N__9663\,
            I => \N__9657\
        );

    \I__1027\ : Span4Mux_h
    port map (
            O => \N__9660\,
            I => \N__9654\
        );

    \I__1026\ : Span12Mux_v
    port map (
            O => \N__9657\,
            I => \N__9651\
        );

    \I__1025\ : Sp12to4
    port map (
            O => \N__9654\,
            I => \N__9648\
        );

    \I__1024\ : Odrv12
    port map (
            O => \N__9651\,
            I => \DEBUG_c_6\
        );

    \I__1023\ : Odrv12
    port map (
            O => \N__9648\,
            I => \DEBUG_c_6\
        );

    \I__1022\ : InMux
    port map (
            O => \N__9643\,
            I => \N__9640\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__9640\,
            I => \transmit_module.video_signal_controller.SYNC_BUFF1\
        );

    \I__1020\ : CascadeMux
    port map (
            O => \N__9637\,
            I => \transmit_module.video_signal_controller.n3987_cascade_\
        );

    \I__1019\ : CascadeMux
    port map (
            O => \N__9634\,
            I => \transmit_module.video_signal_controller.n4_cascade_\
        );

    \I__1018\ : InMux
    port map (
            O => \N__9631\,
            I => \N__9628\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__9628\,
            I => \transmit_module.video_signal_controller.n3935\
        );

    \I__1016\ : CascadeMux
    port map (
            O => \N__9625\,
            I => \N__9622\
        );

    \I__1015\ : InMux
    port map (
            O => \N__9622\,
            I => \N__9616\
        );

    \I__1014\ : InMux
    port map (
            O => \N__9621\,
            I => \N__9613\
        );

    \I__1013\ : InMux
    port map (
            O => \N__9620\,
            I => \N__9610\
        );

    \I__1012\ : InMux
    port map (
            O => \N__9619\,
            I => \N__9607\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__9616\,
            I => \receive_module.rx_counter.Y_1\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__9613\,
            I => \receive_module.rx_counter.Y_1\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__9610\,
            I => \receive_module.rx_counter.Y_1\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__9607\,
            I => \receive_module.rx_counter.Y_1\
        );

    \I__1007\ : InMux
    port map (
            O => \N__9598\,
            I => \receive_module.rx_counter.n3711\
        );

    \I__1006\ : CascadeMux
    port map (
            O => \N__9595\,
            I => \N__9589\
        );

    \I__1005\ : InMux
    port map (
            O => \N__9594\,
            I => \N__9586\
        );

    \I__1004\ : InMux
    port map (
            O => \N__9593\,
            I => \N__9583\
        );

    \I__1003\ : InMux
    port map (
            O => \N__9592\,
            I => \N__9580\
        );

    \I__1002\ : InMux
    port map (
            O => \N__9589\,
            I => \N__9577\
        );

    \I__1001\ : LocalMux
    port map (
            O => \N__9586\,
            I => \receive_module.rx_counter.Y_2\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__9583\,
            I => \receive_module.rx_counter.Y_2\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__9580\,
            I => \receive_module.rx_counter.Y_2\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__9577\,
            I => \receive_module.rx_counter.Y_2\
        );

    \I__997\ : InMux
    port map (
            O => \N__9568\,
            I => \receive_module.rx_counter.n3712\
        );

    \I__996\ : InMux
    port map (
            O => \N__9565\,
            I => \N__9559\
        );

    \I__995\ : InMux
    port map (
            O => \N__9564\,
            I => \N__9556\
        );

    \I__994\ : InMux
    port map (
            O => \N__9563\,
            I => \N__9553\
        );

    \I__993\ : InMux
    port map (
            O => \N__9562\,
            I => \N__9550\
        );

    \I__992\ : LocalMux
    port map (
            O => \N__9559\,
            I => \receive_module.rx_counter.Y_3\
        );

    \I__991\ : LocalMux
    port map (
            O => \N__9556\,
            I => \receive_module.rx_counter.Y_3\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__9553\,
            I => \receive_module.rx_counter.Y_3\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__9550\,
            I => \receive_module.rx_counter.Y_3\
        );

    \I__988\ : InMux
    port map (
            O => \N__9541\,
            I => \receive_module.rx_counter.n3713\
        );

    \I__987\ : InMux
    port map (
            O => \N__9538\,
            I => \N__9532\
        );

    \I__986\ : InMux
    port map (
            O => \N__9537\,
            I => \N__9527\
        );

    \I__985\ : InMux
    port map (
            O => \N__9536\,
            I => \N__9527\
        );

    \I__984\ : InMux
    port map (
            O => \N__9535\,
            I => \N__9524\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__9532\,
            I => \receive_module.rx_counter.Y_4\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__9527\,
            I => \receive_module.rx_counter.Y_4\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__9524\,
            I => \receive_module.rx_counter.Y_4\
        );

    \I__980\ : InMux
    port map (
            O => \N__9517\,
            I => \receive_module.rx_counter.n3714\
        );

    \I__979\ : InMux
    port map (
            O => \N__9514\,
            I => \N__9509\
        );

    \I__978\ : InMux
    port map (
            O => \N__9513\,
            I => \N__9506\
        );

    \I__977\ : InMux
    port map (
            O => \N__9512\,
            I => \N__9503\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__9509\,
            I => \receive_module.rx_counter.Y_5\
        );

    \I__975\ : LocalMux
    port map (
            O => \N__9506\,
            I => \receive_module.rx_counter.Y_5\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__9503\,
            I => \receive_module.rx_counter.Y_5\
        );

    \I__973\ : InMux
    port map (
            O => \N__9496\,
            I => \receive_module.rx_counter.n3715\
        );

    \I__972\ : CascadeMux
    port map (
            O => \N__9493\,
            I => \N__9489\
        );

    \I__971\ : InMux
    port map (
            O => \N__9492\,
            I => \N__9485\
        );

    \I__970\ : InMux
    port map (
            O => \N__9489\,
            I => \N__9482\
        );

    \I__969\ : InMux
    port map (
            O => \N__9488\,
            I => \N__9479\
        );

    \I__968\ : LocalMux
    port map (
            O => \N__9485\,
            I => \receive_module.rx_counter.Y_6\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__9482\,
            I => \receive_module.rx_counter.Y_6\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__9479\,
            I => \receive_module.rx_counter.Y_6\
        );

    \I__965\ : InMux
    port map (
            O => \N__9472\,
            I => \receive_module.rx_counter.n3716\
        );

    \I__964\ : InMux
    port map (
            O => \N__9469\,
            I => \N__9463\
        );

    \I__963\ : InMux
    port map (
            O => \N__9468\,
            I => \N__9458\
        );

    \I__962\ : InMux
    port map (
            O => \N__9467\,
            I => \N__9458\
        );

    \I__961\ : InMux
    port map (
            O => \N__9466\,
            I => \N__9455\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__9463\,
            I => \receive_module.rx_counter.Y_7\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__9458\,
            I => \receive_module.rx_counter.Y_7\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__9455\,
            I => \receive_module.rx_counter.Y_7\
        );

    \I__957\ : InMux
    port map (
            O => \N__9448\,
            I => \receive_module.rx_counter.n3717\
        );

    \I__956\ : InMux
    port map (
            O => \N__9445\,
            I => \N__9439\
        );

    \I__955\ : InMux
    port map (
            O => \N__9444\,
            I => \N__9436\
        );

    \I__954\ : InMux
    port map (
            O => \N__9443\,
            I => \N__9433\
        );

    \I__953\ : InMux
    port map (
            O => \N__9442\,
            I => \N__9430\
        );

    \I__952\ : LocalMux
    port map (
            O => \N__9439\,
            I => \receive_module.rx_counter.Y_8\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__9436\,
            I => \receive_module.rx_counter.Y_8\
        );

    \I__950\ : LocalMux
    port map (
            O => \N__9433\,
            I => \receive_module.rx_counter.Y_8\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__9430\,
            I => \receive_module.rx_counter.Y_8\
        );

    \I__948\ : InMux
    port map (
            O => \N__9421\,
            I => \N__9418\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__9418\,
            I => \transmit_module.Y_DELTA_PATTERN_89\
        );

    \I__946\ : InMux
    port map (
            O => \N__9415\,
            I => \N__9412\
        );

    \I__945\ : LocalMux
    port map (
            O => \N__9412\,
            I => \transmit_module.Y_DELTA_PATTERN_88\
        );

    \I__944\ : InMux
    port map (
            O => \N__9409\,
            I => \N__9406\
        );

    \I__943\ : LocalMux
    port map (
            O => \N__9406\,
            I => \transmit_module.Y_DELTA_PATTERN_87\
        );

    \I__942\ : InMux
    port map (
            O => \N__9403\,
            I => \N__9400\
        );

    \I__941\ : LocalMux
    port map (
            O => \N__9400\,
            I => \transmit_module.Y_DELTA_PATTERN_92\
        );

    \I__940\ : InMux
    port map (
            O => \N__9397\,
            I => \N__9394\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__9394\,
            I => \transmit_module.Y_DELTA_PATTERN_91\
        );

    \I__938\ : InMux
    port map (
            O => \N__9391\,
            I => \N__9388\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__9388\,
            I => \transmit_module.Y_DELTA_PATTERN_86\
        );

    \I__936\ : InMux
    port map (
            O => \N__9385\,
            I => \N__9382\
        );

    \I__935\ : LocalMux
    port map (
            O => \N__9382\,
            I => \N__9379\
        );

    \I__934\ : Odrv4
    port map (
            O => \N__9379\,
            I => \transmit_module.Y_DELTA_PATTERN_85\
        );

    \I__933\ : InMux
    port map (
            O => \N__9376\,
            I => \N__9373\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__9373\,
            I => \transmit_module.Y_DELTA_PATTERN_94\
        );

    \I__931\ : InMux
    port map (
            O => \N__9370\,
            I => \N__9367\
        );

    \I__930\ : LocalMux
    port map (
            O => \N__9367\,
            I => \transmit_module.Y_DELTA_PATTERN_93\
        );

    \I__929\ : InMux
    port map (
            O => \N__9364\,
            I => \N__9361\
        );

    \I__928\ : LocalMux
    port map (
            O => \N__9361\,
            I => \transmit_module.Y_DELTA_PATTERN_96\
        );

    \I__927\ : InMux
    port map (
            O => \N__9358\,
            I => \N__9355\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__9355\,
            I => \transmit_module.Y_DELTA_PATTERN_97\
        );

    \I__925\ : InMux
    port map (
            O => \N__9352\,
            I => \N__9349\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__9349\,
            I => \N__9346\
        );

    \I__923\ : Odrv4
    port map (
            O => \N__9346\,
            I => \line_buffer.n624\
        );

    \I__922\ : InMux
    port map (
            O => \N__9343\,
            I => \N__9340\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__9340\,
            I => \line_buffer.n4122\
        );

    \I__920\ : CascadeMux
    port map (
            O => \N__9337\,
            I => \N__9334\
        );

    \I__919\ : InMux
    port map (
            O => \N__9334\,
            I => \N__9331\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__9331\,
            I => \N__9328\
        );

    \I__917\ : Span4Mux_h
    port map (
            O => \N__9328\,
            I => \N__9325\
        );

    \I__916\ : Span4Mux_h
    port map (
            O => \N__9325\,
            I => \N__9322\
        );

    \I__915\ : Sp12to4
    port map (
            O => \N__9322\,
            I => \N__9319\
        );

    \I__914\ : Span12Mux_v
    port map (
            O => \N__9319\,
            I => \N__9316\
        );

    \I__913\ : Span12Mux_v
    port map (
            O => \N__9316\,
            I => \N__9313\
        );

    \I__912\ : Odrv12
    port map (
            O => \N__9313\,
            I => \line_buffer.n616\
        );

    \I__911\ : InMux
    port map (
            O => \N__9310\,
            I => \N__9304\
        );

    \I__910\ : InMux
    port map (
            O => \N__9309\,
            I => \N__9301\
        );

    \I__909\ : InMux
    port map (
            O => \N__9308\,
            I => \N__9298\
        );

    \I__908\ : InMux
    port map (
            O => \N__9307\,
            I => \N__9295\
        );

    \I__907\ : LocalMux
    port map (
            O => \N__9304\,
            I => \receive_module.rx_counter.Y_0\
        );

    \I__906\ : LocalMux
    port map (
            O => \N__9301\,
            I => \receive_module.rx_counter.Y_0\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__9298\,
            I => \receive_module.rx_counter.Y_0\
        );

    \I__904\ : LocalMux
    port map (
            O => \N__9295\,
            I => \receive_module.rx_counter.Y_0\
        );

    \I__903\ : InMux
    port map (
            O => \N__9286\,
            I => \bfn_11_9_0_\
        );

    \I__902\ : InMux
    port map (
            O => \N__9283\,
            I => \receive_module.rx_counter.n3674\
        );

    \I__901\ : InMux
    port map (
            O => \N__9280\,
            I => \receive_module.rx_counter.n3675\
        );

    \I__900\ : InMux
    port map (
            O => \N__9277\,
            I => \bfn_10_10_0_\
        );

    \I__899\ : InMux
    port map (
            O => \N__9274\,
            I => \N__9271\
        );

    \I__898\ : LocalMux
    port map (
            O => \N__9271\,
            I => \transmit_module.Y_DELTA_PATTERN_84\
        );

    \I__897\ : InMux
    port map (
            O => \N__9268\,
            I => \N__9265\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__9265\,
            I => \transmit_module.Y_DELTA_PATTERN_83\
        );

    \I__895\ : InMux
    port map (
            O => \N__9262\,
            I => \N__9259\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__9259\,
            I => \transmit_module.Y_DELTA_PATTERN_90\
        );

    \I__893\ : InMux
    port map (
            O => \N__9256\,
            I => \N__9253\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__9253\,
            I => \transmit_module.Y_DELTA_PATTERN_95\
        );

    \I__891\ : InMux
    port map (
            O => \N__9250\,
            I => \N__9247\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__9247\,
            I => \N__9244\
        );

    \I__889\ : Span4Mux_v
    port map (
            O => \N__9244\,
            I => \N__9241\
        );

    \I__888\ : Odrv4
    port map (
            O => \N__9241\,
            I => \line_buffer.n680\
        );

    \I__887\ : CascadeMux
    port map (
            O => \N__9238\,
            I => \N__9235\
        );

    \I__886\ : InMux
    port map (
            O => \N__9235\,
            I => \N__9232\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__9232\,
            I => \N__9229\
        );

    \I__884\ : Span4Mux_h
    port map (
            O => \N__9229\,
            I => \N__9226\
        );

    \I__883\ : Odrv4
    port map (
            O => \N__9226\,
            I => \line_buffer.n688\
        );

    \I__882\ : InMux
    port map (
            O => \N__9223\,
            I => \bfn_10_9_0_\
        );

    \I__881\ : InMux
    port map (
            O => \N__9220\,
            I => \receive_module.rx_counter.n3669\
        );

    \I__880\ : InMux
    port map (
            O => \N__9217\,
            I => \receive_module.rx_counter.n3670\
        );

    \I__879\ : InMux
    port map (
            O => \N__9214\,
            I => \receive_module.rx_counter.n3671\
        );

    \I__878\ : InMux
    port map (
            O => \N__9211\,
            I => \receive_module.rx_counter.n3672\
        );

    \I__877\ : InMux
    port map (
            O => \N__9208\,
            I => \receive_module.rx_counter.n3673\
        );

    \I__876\ : CascadeMux
    port map (
            O => \N__9205\,
            I => \receive_module.rx_counter.n3176_cascade_\
        );

    \I__875\ : InMux
    port map (
            O => \N__9202\,
            I => \N__9199\
        );

    \I__874\ : LocalMux
    port map (
            O => \N__9199\,
            I => \receive_module.rx_counter.n3208\
        );

    \I__873\ : InMux
    port map (
            O => \N__9196\,
            I => \N__9193\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__9193\,
            I => \N__9190\
        );

    \I__871\ : Span4Mux_v
    port map (
            O => \N__9190\,
            I => \N__9187\
        );

    \I__870\ : Sp12to4
    port map (
            O => \N__9187\,
            I => \N__9184\
        );

    \I__869\ : Span12Mux_h
    port map (
            O => \N__9184\,
            I => \N__9181\
        );

    \I__868\ : Span12Mux_v
    port map (
            O => \N__9181\,
            I => \N__9178\
        );

    \I__867\ : Odrv12
    port map (
            O => \N__9178\,
            I => \line_buffer.n675\
        );

    \I__866\ : InMux
    port map (
            O => \N__9175\,
            I => \N__9172\
        );

    \I__865\ : LocalMux
    port map (
            O => \N__9172\,
            I => \N__9169\
        );

    \I__864\ : Odrv4
    port map (
            O => \N__9169\,
            I => \line_buffer.n683\
        );

    \I__863\ : InMux
    port map (
            O => \N__9166\,
            I => \N__9163\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__9163\,
            I => \N__9160\
        );

    \I__861\ : Span4Mux_v
    port map (
            O => \N__9160\,
            I => \N__9157\
        );

    \I__860\ : Span4Mux_h
    port map (
            O => \N__9157\,
            I => \N__9154\
        );

    \I__859\ : Sp12to4
    port map (
            O => \N__9154\,
            I => \N__9151\
        );

    \I__858\ : Span12Mux_h
    port map (
            O => \N__9151\,
            I => \N__9148\
        );

    \I__857\ : Odrv12
    port map (
            O => \N__9148\,
            I => \line_buffer.n611\
        );

    \I__856\ : CascadeMux
    port map (
            O => \N__9145\,
            I => \line_buffer.n4170_cascade_\
        );

    \I__855\ : InMux
    port map (
            O => \N__9142\,
            I => \N__9139\
        );

    \I__854\ : LocalMux
    port map (
            O => \N__9139\,
            I => \N__9136\
        );

    \I__853\ : Span4Mux_v
    port map (
            O => \N__9136\,
            I => \N__9133\
        );

    \I__852\ : Span4Mux_v
    port map (
            O => \N__9133\,
            I => \N__9130\
        );

    \I__851\ : Odrv4
    port map (
            O => \N__9130\,
            I => \line_buffer.n619\
        );

    \I__850\ : InMux
    port map (
            O => \N__9127\,
            I => \N__9124\
        );

    \I__849\ : LocalMux
    port map (
            O => \N__9124\,
            I => \N__9121\
        );

    \I__848\ : Span4Mux_v
    port map (
            O => \N__9121\,
            I => \N__9118\
        );

    \I__847\ : Sp12to4
    port map (
            O => \N__9118\,
            I => \N__9115\
        );

    \I__846\ : Span12Mux_h
    port map (
            O => \N__9115\,
            I => \N__9112\
        );

    \I__845\ : Odrv12
    port map (
            O => \N__9112\,
            I => \line_buffer.n643\
        );

    \I__844\ : CascadeMux
    port map (
            O => \N__9109\,
            I => \N__9106\
        );

    \I__843\ : InMux
    port map (
            O => \N__9106\,
            I => \N__9103\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__9103\,
            I => \N__9100\
        );

    \I__841\ : Span4Mux_v
    port map (
            O => \N__9100\,
            I => \N__9097\
        );

    \I__840\ : Odrv4
    port map (
            O => \N__9097\,
            I => \line_buffer.n651\
        );

    \I__839\ : InMux
    port map (
            O => \N__9094\,
            I => \N__9091\
        );

    \I__838\ : LocalMux
    port map (
            O => \N__9091\,
            I => \N__9088\
        );

    \I__837\ : Span4Mux_v
    port map (
            O => \N__9088\,
            I => \N__9085\
        );

    \I__836\ : Span4Mux_v
    port map (
            O => \N__9085\,
            I => \N__9082\
        );

    \I__835\ : Odrv4
    port map (
            O => \N__9082\,
            I => \line_buffer.n687\
        );

    \I__834\ : InMux
    port map (
            O => \N__9079\,
            I => \N__9076\
        );

    \I__833\ : LocalMux
    port map (
            O => \N__9076\,
            I => \line_buffer.n679\
        );

    \I__832\ : InMux
    port map (
            O => \N__9073\,
            I => \N__9070\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__9070\,
            I => \line_buffer.n4152\
        );

    \I__830\ : InMux
    port map (
            O => \N__9067\,
            I => \N__9064\
        );

    \I__829\ : LocalMux
    port map (
            O => \N__9064\,
            I => \N__9061\
        );

    \I__828\ : Span4Mux_h
    port map (
            O => \N__9061\,
            I => \N__9058\
        );

    \I__827\ : Sp12to4
    port map (
            O => \N__9058\,
            I => \N__9055\
        );

    \I__826\ : Span12Mux_v
    port map (
            O => \N__9055\,
            I => \N__9052\
        );

    \I__825\ : Span12Mux_h
    port map (
            O => \N__9052\,
            I => \N__9049\
        );

    \I__824\ : Odrv12
    port map (
            O => \N__9049\,
            I => \line_buffer.n554\
        );

    \I__823\ : CascadeMux
    port map (
            O => \N__9046\,
            I => \N__9043\
        );

    \I__822\ : InMux
    port map (
            O => \N__9043\,
            I => \N__9040\
        );

    \I__821\ : LocalMux
    port map (
            O => \N__9040\,
            I => \N__9037\
        );

    \I__820\ : Span4Mux_h
    port map (
            O => \N__9037\,
            I => \N__9034\
        );

    \I__819\ : Sp12to4
    port map (
            O => \N__9034\,
            I => \N__9031\
        );

    \I__818\ : Span12Mux_v
    port map (
            O => \N__9031\,
            I => \N__9028\
        );

    \I__817\ : Odrv12
    port map (
            O => \N__9028\,
            I => \line_buffer.n546\
        );

    \I__816\ : CascadeMux
    port map (
            O => \N__9025\,
            I => \line_buffer.n4155_cascade_\
        );

    \I__815\ : InMux
    port map (
            O => \N__9022\,
            I => \N__9019\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__9019\,
            I => \line_buffer.n4173\
        );

    \I__813\ : InMux
    port map (
            O => \N__9016\,
            I => \N__9013\
        );

    \I__812\ : LocalMux
    port map (
            O => \N__9013\,
            I => \N__9010\
        );

    \I__811\ : Span4Mux_s2_v
    port map (
            O => \N__9010\,
            I => \N__9006\
        );

    \I__810\ : InMux
    port map (
            O => \N__9009\,
            I => \N__9003\
        );

    \I__809\ : Span4Mux_v
    port map (
            O => \N__9006\,
            I => \N__8998\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__9003\,
            I => \N__8998\
        );

    \I__807\ : Span4Mux_v
    port map (
            O => \N__8998\,
            I => \N__8994\
        );

    \I__806\ : InMux
    port map (
            O => \N__8997\,
            I => \N__8991\
        );

    \I__805\ : Span4Mux_v
    port map (
            O => \N__8994\,
            I => \N__8985\
        );

    \I__804\ : LocalMux
    port map (
            O => \N__8991\,
            I => \N__8985\
        );

    \I__803\ : InMux
    port map (
            O => \N__8990\,
            I => \N__8982\
        );

    \I__802\ : Span4Mux_v
    port map (
            O => \N__8985\,
            I => \N__8979\
        );

    \I__801\ : LocalMux
    port map (
            O => \N__8982\,
            I => \N__8976\
        );

    \I__800\ : Span4Mux_v
    port map (
            O => \N__8979\,
            I => \N__8969\
        );

    \I__799\ : Span4Mux_v
    port map (
            O => \N__8976\,
            I => \N__8969\
        );

    \I__798\ : InMux
    port map (
            O => \N__8975\,
            I => \N__8966\
        );

    \I__797\ : InMux
    port map (
            O => \N__8974\,
            I => \N__8963\
        );

    \I__796\ : Span4Mux_v
    port map (
            O => \N__8969\,
            I => \N__8958\
        );

    \I__795\ : LocalMux
    port map (
            O => \N__8966\,
            I => \N__8958\
        );

    \I__794\ : LocalMux
    port map (
            O => \N__8963\,
            I => \N__8955\
        );

    \I__793\ : Span4Mux_h
    port map (
            O => \N__8958\,
            I => \N__8951\
        );

    \I__792\ : Span4Mux_h
    port map (
            O => \N__8955\,
            I => \N__8948\
        );

    \I__791\ : InMux
    port map (
            O => \N__8954\,
            I => \N__8945\
        );

    \I__790\ : Span4Mux_h
    port map (
            O => \N__8951\,
            I => \N__8942\
        );

    \I__789\ : Span4Mux_v
    port map (
            O => \N__8948\,
            I => \N__8938\
        );

    \I__788\ : LocalMux
    port map (
            O => \N__8945\,
            I => \N__8935\
        );

    \I__787\ : Span4Mux_h
    port map (
            O => \N__8942\,
            I => \N__8932\
        );

    \I__786\ : InMux
    port map (
            O => \N__8941\,
            I => \N__8929\
        );

    \I__785\ : Span4Mux_v
    port map (
            O => \N__8938\,
            I => \N__8924\
        );

    \I__784\ : Span4Mux_h
    port map (
            O => \N__8935\,
            I => \N__8924\
        );

    \I__783\ : Span4Mux_h
    port map (
            O => \N__8932\,
            I => \N__8919\
        );

    \I__782\ : LocalMux
    port map (
            O => \N__8929\,
            I => \N__8919\
        );

    \I__781\ : Span4Mux_v
    port map (
            O => \N__8924\,
            I => \N__8916\
        );

    \I__780\ : Span4Mux_h
    port map (
            O => \N__8919\,
            I => \N__8913\
        );

    \I__779\ : Span4Mux_v
    port map (
            O => \N__8916\,
            I => \N__8910\
        );

    \I__778\ : Span4Mux_v
    port map (
            O => \N__8913\,
            I => \N__8907\
        );

    \I__777\ : Odrv4
    port map (
            O => \N__8910\,
            I => \TVP_VIDEO_c_2\
        );

    \I__776\ : Odrv4
    port map (
            O => \N__8907\,
            I => \TVP_VIDEO_c_2\
        );

    \I__775\ : CascadeMux
    port map (
            O => \N__8902\,
            I => \receive_module.rx_counter.n12_cascade_\
        );

    \I__774\ : CascadeMux
    port map (
            O => \N__8899\,
            I => \receive_module.rx_counter.n3938_cascade_\
        );

    \I__773\ : InMux
    port map (
            O => \N__8896\,
            I => \N__8893\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__8893\,
            I => \receive_module.rx_counter.n3938\
        );

    \I__771\ : InMux
    port map (
            O => \N__8890\,
            I => \N__8887\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__8887\,
            I => \receive_module.rx_counter.n13\
        );

    \I__769\ : InMux
    port map (
            O => \N__8884\,
            I => \N__8880\
        );

    \I__768\ : InMux
    port map (
            O => \N__8883\,
            I => \N__8877\
        );

    \I__767\ : LocalMux
    port map (
            O => \N__8880\,
            I => \N__8870\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__8877\,
            I => \N__8870\
        );

    \I__765\ : InMux
    port map (
            O => \N__8876\,
            I => \N__8867\
        );

    \I__764\ : InMux
    port map (
            O => \N__8875\,
            I => \N__8864\
        );

    \I__763\ : Span4Mux_v
    port map (
            O => \N__8870\,
            I => \N__8857\
        );

    \I__762\ : LocalMux
    port map (
            O => \N__8867\,
            I => \N__8857\
        );

    \I__761\ : LocalMux
    port map (
            O => \N__8864\,
            I => \N__8857\
        );

    \I__760\ : Span4Mux_v
    port map (
            O => \N__8857\,
            I => \N__8852\
        );

    \I__759\ : InMux
    port map (
            O => \N__8856\,
            I => \N__8849\
        );

    \I__758\ : InMux
    port map (
            O => \N__8855\,
            I => \N__8846\
        );

    \I__757\ : Span4Mux_v
    port map (
            O => \N__8852\,
            I => \N__8841\
        );

    \I__756\ : LocalMux
    port map (
            O => \N__8849\,
            I => \N__8841\
        );

    \I__755\ : LocalMux
    port map (
            O => \N__8846\,
            I => \N__8836\
        );

    \I__754\ : Span4Mux_h
    port map (
            O => \N__8841\,
            I => \N__8833\
        );

    \I__753\ : InMux
    port map (
            O => \N__8840\,
            I => \N__8830\
        );

    \I__752\ : InMux
    port map (
            O => \N__8839\,
            I => \N__8827\
        );

    \I__751\ : Span4Mux_v
    port map (
            O => \N__8836\,
            I => \N__8824\
        );

    \I__750\ : Span4Mux_h
    port map (
            O => \N__8833\,
            I => \N__8821\
        );

    \I__749\ : LocalMux
    port map (
            O => \N__8830\,
            I => \N__8818\
        );

    \I__748\ : LocalMux
    port map (
            O => \N__8827\,
            I => \N__8815\
        );

    \I__747\ : Sp12to4
    port map (
            O => \N__8824\,
            I => \N__8812\
        );

    \I__746\ : Span4Mux_v
    port map (
            O => \N__8821\,
            I => \N__8809\
        );

    \I__745\ : Span4Mux_h
    port map (
            O => \N__8818\,
            I => \N__8806\
        );

    \I__744\ : Span4Mux_h
    port map (
            O => \N__8815\,
            I => \N__8803\
        );

    \I__743\ : Span12Mux_h
    port map (
            O => \N__8812\,
            I => \N__8800\
        );

    \I__742\ : Span4Mux_v
    port map (
            O => \N__8809\,
            I => \N__8797\
        );

    \I__741\ : Span4Mux_h
    port map (
            O => \N__8806\,
            I => \N__8794\
        );

    \I__740\ : Span4Mux_h
    port map (
            O => \N__8803\,
            I => \N__8791\
        );

    \I__739\ : Span12Mux_v
    port map (
            O => \N__8800\,
            I => \N__8788\
        );

    \I__738\ : Span4Mux_v
    port map (
            O => \N__8797\,
            I => \N__8783\
        );

    \I__737\ : Span4Mux_h
    port map (
            O => \N__8794\,
            I => \N__8783\
        );

    \I__736\ : Span4Mux_h
    port map (
            O => \N__8791\,
            I => \N__8780\
        );

    \I__735\ : Odrv12
    port map (
            O => \N__8788\,
            I => \TVP_VIDEO_c_8\
        );

    \I__734\ : Odrv4
    port map (
            O => \N__8783\,
            I => \TVP_VIDEO_c_8\
        );

    \I__733\ : Odrv4
    port map (
            O => \N__8780\,
            I => \TVP_VIDEO_c_8\
        );

    \I__732\ : InMux
    port map (
            O => \N__8773\,
            I => \N__8769\
        );

    \I__731\ : InMux
    port map (
            O => \N__8772\,
            I => \N__8766\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__8769\,
            I => \N__8760\
        );

    \I__729\ : LocalMux
    port map (
            O => \N__8766\,
            I => \N__8760\
        );

    \I__728\ : InMux
    port map (
            O => \N__8765\,
            I => \N__8757\
        );

    \I__727\ : Span4Mux_v
    port map (
            O => \N__8760\,
            I => \N__8752\
        );

    \I__726\ : LocalMux
    port map (
            O => \N__8757\,
            I => \N__8752\
        );

    \I__725\ : Span4Mux_v
    port map (
            O => \N__8752\,
            I => \N__8747\
        );

    \I__724\ : InMux
    port map (
            O => \N__8751\,
            I => \N__8744\
        );

    \I__723\ : InMux
    port map (
            O => \N__8750\,
            I => \N__8740\
        );

    \I__722\ : Span4Mux_v
    port map (
            O => \N__8747\,
            I => \N__8735\
        );

    \I__721\ : LocalMux
    port map (
            O => \N__8744\,
            I => \N__8735\
        );

    \I__720\ : InMux
    port map (
            O => \N__8743\,
            I => \N__8732\
        );

    \I__719\ : LocalMux
    port map (
            O => \N__8740\,
            I => \N__8729\
        );

    \I__718\ : Span4Mux_h
    port map (
            O => \N__8735\,
            I => \N__8726\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__8732\,
            I => \N__8723\
        );

    \I__716\ : Span12Mux_s11_h
    port map (
            O => \N__8729\,
            I => \N__8719\
        );

    \I__715\ : Sp12to4
    port map (
            O => \N__8726\,
            I => \N__8716\
        );

    \I__714\ : Span12Mux_s8_h
    port map (
            O => \N__8723\,
            I => \N__8713\
        );

    \I__713\ : InMux
    port map (
            O => \N__8722\,
            I => \N__8710\
        );

    \I__712\ : Span12Mux_h
    port map (
            O => \N__8719\,
            I => \N__8707\
        );

    \I__711\ : Span12Mux_v
    port map (
            O => \N__8716\,
            I => \N__8704\
        );

    \I__710\ : Span12Mux_v
    port map (
            O => \N__8713\,
            I => \N__8701\
        );

    \I__709\ : LocalMux
    port map (
            O => \N__8710\,
            I => \N__8698\
        );

    \I__708\ : Span12Mux_v
    port map (
            O => \N__8707\,
            I => \N__8694\
        );

    \I__707\ : Span12Mux_h
    port map (
            O => \N__8704\,
            I => \N__8691\
        );

    \I__706\ : Span12Mux_v
    port map (
            O => \N__8701\,
            I => \N__8688\
        );

    \I__705\ : Span4Mux_h
    port map (
            O => \N__8698\,
            I => \N__8685\
        );

    \I__704\ : InMux
    port map (
            O => \N__8697\,
            I => \N__8682\
        );

    \I__703\ : Odrv12
    port map (
            O => \N__8694\,
            I => \TVP_VIDEO_c_9\
        );

    \I__702\ : Odrv12
    port map (
            O => \N__8691\,
            I => \TVP_VIDEO_c_9\
        );

    \I__701\ : Odrv12
    port map (
            O => \N__8688\,
            I => \TVP_VIDEO_c_9\
        );

    \I__700\ : Odrv4
    port map (
            O => \N__8685\,
            I => \TVP_VIDEO_c_9\
        );

    \I__699\ : LocalMux
    port map (
            O => \N__8682\,
            I => \TVP_VIDEO_c_9\
        );

    \I__698\ : InMux
    port map (
            O => \N__8671\,
            I => \N__8668\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__8668\,
            I => \N__8662\
        );

    \I__696\ : InMux
    port map (
            O => \N__8667\,
            I => \N__8659\
        );

    \I__695\ : InMux
    port map (
            O => \N__8666\,
            I => \N__8656\
        );

    \I__694\ : InMux
    port map (
            O => \N__8665\,
            I => \N__8653\
        );

    \I__693\ : Span4Mux_h
    port map (
            O => \N__8662\,
            I => \N__8650\
        );

    \I__692\ : LocalMux
    port map (
            O => \N__8659\,
            I => \N__8646\
        );

    \I__691\ : LocalMux
    port map (
            O => \N__8656\,
            I => \N__8643\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__8653\,
            I => \N__8639\
        );

    \I__689\ : Span4Mux_h
    port map (
            O => \N__8650\,
            I => \N__8636\
        );

    \I__688\ : InMux
    port map (
            O => \N__8649\,
            I => \N__8633\
        );

    \I__687\ : Span4Mux_h
    port map (
            O => \N__8646\,
            I => \N__8630\
        );

    \I__686\ : Span4Mux_v
    port map (
            O => \N__8643\,
            I => \N__8627\
        );

    \I__685\ : InMux
    port map (
            O => \N__8642\,
            I => \N__8622\
        );

    \I__684\ : Span12Mux_h
    port map (
            O => \N__8639\,
            I => \N__8619\
        );

    \I__683\ : Sp12to4
    port map (
            O => \N__8636\,
            I => \N__8616\
        );

    \I__682\ : LocalMux
    port map (
            O => \N__8633\,
            I => \N__8613\
        );

    \I__681\ : Span4Mux_h
    port map (
            O => \N__8630\,
            I => \N__8610\
        );

    \I__680\ : Span4Mux_v
    port map (
            O => \N__8627\,
            I => \N__8607\
        );

    \I__679\ : InMux
    port map (
            O => \N__8626\,
            I => \N__8604\
        );

    \I__678\ : InMux
    port map (
            O => \N__8625\,
            I => \N__8601\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__8622\,
            I => \N__8598\
        );

    \I__676\ : Span12Mux_v
    port map (
            O => \N__8619\,
            I => \N__8595\
        );

    \I__675\ : Span12Mux_v
    port map (
            O => \N__8616\,
            I => \N__8588\
        );

    \I__674\ : Span12Mux_h
    port map (
            O => \N__8613\,
            I => \N__8588\
        );

    \I__673\ : Sp12to4
    port map (
            O => \N__8610\,
            I => \N__8588\
        );

    \I__672\ : Sp12to4
    port map (
            O => \N__8607\,
            I => \N__8583\
        );

    \I__671\ : LocalMux
    port map (
            O => \N__8604\,
            I => \N__8583\
        );

    \I__670\ : LocalMux
    port map (
            O => \N__8601\,
            I => \N__8580\
        );

    \I__669\ : Span4Mux_h
    port map (
            O => \N__8598\,
            I => \N__8577\
        );

    \I__668\ : Span12Mux_v
    port map (
            O => \N__8595\,
            I => \N__8574\
        );

    \I__667\ : Span12Mux_v
    port map (
            O => \N__8588\,
            I => \N__8567\
        );

    \I__666\ : Span12Mux_h
    port map (
            O => \N__8583\,
            I => \N__8567\
        );

    \I__665\ : Span12Mux_h
    port map (
            O => \N__8580\,
            I => \N__8567\
        );

    \I__664\ : Span4Mux_h
    port map (
            O => \N__8577\,
            I => \N__8564\
        );

    \I__663\ : Odrv12
    port map (
            O => \N__8574\,
            I => \TVP_VIDEO_c_7\
        );

    \I__662\ : Odrv12
    port map (
            O => \N__8567\,
            I => \TVP_VIDEO_c_7\
        );

    \I__661\ : Odrv4
    port map (
            O => \N__8564\,
            I => \TVP_VIDEO_c_7\
        );

    \I__660\ : InMux
    port map (
            O => \N__8557\,
            I => \N__8553\
        );

    \I__659\ : InMux
    port map (
            O => \N__8556\,
            I => \N__8550\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__8553\,
            I => \N__8547\
        );

    \I__657\ : LocalMux
    port map (
            O => \N__8550\,
            I => \N__8543\
        );

    \I__656\ : Span4Mux_v
    port map (
            O => \N__8547\,
            I => \N__8540\
        );

    \I__655\ : InMux
    port map (
            O => \N__8546\,
            I => \N__8537\
        );

    \I__654\ : Span4Mux_v
    port map (
            O => \N__8543\,
            I => \N__8533\
        );

    \I__653\ : Span4Mux_v
    port map (
            O => \N__8540\,
            I => \N__8528\
        );

    \I__652\ : LocalMux
    port map (
            O => \N__8537\,
            I => \N__8528\
        );

    \I__651\ : InMux
    port map (
            O => \N__8536\,
            I => \N__8525\
        );

    \I__650\ : Span4Mux_v
    port map (
            O => \N__8533\,
            I => \N__8522\
        );

    \I__649\ : Span4Mux_v
    port map (
            O => \N__8528\,
            I => \N__8516\
        );

    \I__648\ : LocalMux
    port map (
            O => \N__8525\,
            I => \N__8516\
        );

    \I__647\ : Span4Mux_v
    port map (
            O => \N__8522\,
            I => \N__8512\
        );

    \I__646\ : InMux
    port map (
            O => \N__8521\,
            I => \N__8509\
        );

    \I__645\ : Span4Mux_v
    port map (
            O => \N__8516\,
            I => \N__8505\
        );

    \I__644\ : InMux
    port map (
            O => \N__8515\,
            I => \N__8502\
        );

    \I__643\ : Span4Mux_v
    port map (
            O => \N__8512\,
            I => \N__8497\
        );

    \I__642\ : LocalMux
    port map (
            O => \N__8509\,
            I => \N__8497\
        );

    \I__641\ : InMux
    port map (
            O => \N__8508\,
            I => \N__8494\
        );

    \I__640\ : Span4Mux_v
    port map (
            O => \N__8505\,
            I => \N__8489\
        );

    \I__639\ : LocalMux
    port map (
            O => \N__8502\,
            I => \N__8489\
        );

    \I__638\ : Span4Mux_v
    port map (
            O => \N__8497\,
            I => \N__8484\
        );

    \I__637\ : LocalMux
    port map (
            O => \N__8494\,
            I => \N__8484\
        );

    \I__636\ : Span4Mux_v
    port map (
            O => \N__8489\,
            I => \N__8480\
        );

    \I__635\ : Span4Mux_v
    port map (
            O => \N__8484\,
            I => \N__8477\
        );

    \I__634\ : InMux
    port map (
            O => \N__8483\,
            I => \N__8474\
        );

    \I__633\ : Sp12to4
    port map (
            O => \N__8480\,
            I => \N__8471\
        );

    \I__632\ : Span4Mux_v
    port map (
            O => \N__8477\,
            I => \N__8466\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__8474\,
            I => \N__8466\
        );

    \I__630\ : Span12Mux_h
    port map (
            O => \N__8471\,
            I => \N__8463\
        );

    \I__629\ : Span4Mux_h
    port map (
            O => \N__8466\,
            I => \N__8460\
        );

    \I__628\ : Odrv12
    port map (
            O => \N__8463\,
            I => \TVP_VIDEO_c_6\
        );

    \I__627\ : Odrv4
    port map (
            O => \N__8460\,
            I => \TVP_VIDEO_c_6\
        );

    \I__626\ : InMux
    port map (
            O => \N__8455\,
            I => \N__8452\
        );

    \I__625\ : LocalMux
    port map (
            O => \N__8452\,
            I => \N__8448\
        );

    \I__624\ : InMux
    port map (
            O => \N__8451\,
            I => \N__8444\
        );

    \I__623\ : Span4Mux_v
    port map (
            O => \N__8448\,
            I => \N__8441\
        );

    \I__622\ : InMux
    port map (
            O => \N__8447\,
            I => \N__8437\
        );

    \I__621\ : LocalMux
    port map (
            O => \N__8444\,
            I => \N__8434\
        );

    \I__620\ : Span4Mux_v
    port map (
            O => \N__8441\,
            I => \N__8430\
        );

    \I__619\ : InMux
    port map (
            O => \N__8440\,
            I => \N__8427\
        );

    \I__618\ : LocalMux
    port map (
            O => \N__8437\,
            I => \N__8424\
        );

    \I__617\ : Span4Mux_v
    port map (
            O => \N__8434\,
            I => \N__8421\
        );

    \I__616\ : InMux
    port map (
            O => \N__8433\,
            I => \N__8418\
        );

    \I__615\ : Span4Mux_v
    port map (
            O => \N__8430\,
            I => \N__8412\
        );

    \I__614\ : LocalMux
    port map (
            O => \N__8427\,
            I => \N__8412\
        );

    \I__613\ : Span4Mux_h
    port map (
            O => \N__8424\,
            I => \N__8408\
        );

    \I__612\ : Span4Mux_v
    port map (
            O => \N__8421\,
            I => \N__8403\
        );

    \I__611\ : LocalMux
    port map (
            O => \N__8418\,
            I => \N__8403\
        );

    \I__610\ : InMux
    port map (
            O => \N__8417\,
            I => \N__8400\
        );

    \I__609\ : Span4Mux_v
    port map (
            O => \N__8412\,
            I => \N__8397\
        );

    \I__608\ : InMux
    port map (
            O => \N__8411\,
            I => \N__8394\
        );

    \I__607\ : Sp12to4
    port map (
            O => \N__8408\,
            I => \N__8391\
        );

    \I__606\ : Span4Mux_v
    port map (
            O => \N__8403\,
            I => \N__8386\
        );

    \I__605\ : LocalMux
    port map (
            O => \N__8400\,
            I => \N__8386\
        );

    \I__604\ : Span4Mux_v
    port map (
            O => \N__8397\,
            I => \N__8381\
        );

    \I__603\ : LocalMux
    port map (
            O => \N__8394\,
            I => \N__8381\
        );

    \I__602\ : Span12Mux_v
    port map (
            O => \N__8391\,
            I => \N__8377\
        );

    \I__601\ : Span4Mux_v
    port map (
            O => \N__8386\,
            I => \N__8374\
        );

    \I__600\ : Span4Mux_v
    port map (
            O => \N__8381\,
            I => \N__8371\
        );

    \I__599\ : InMux
    port map (
            O => \N__8380\,
            I => \N__8368\
        );

    \I__598\ : Span12Mux_v
    port map (
            O => \N__8377\,
            I => \N__8363\
        );

    \I__597\ : Sp12to4
    port map (
            O => \N__8374\,
            I => \N__8363\
        );

    \I__596\ : Span4Mux_v
    port map (
            O => \N__8371\,
            I => \N__8358\
        );

    \I__595\ : LocalMux
    port map (
            O => \N__8368\,
            I => \N__8358\
        );

    \I__594\ : Span12Mux_h
    port map (
            O => \N__8363\,
            I => \N__8355\
        );

    \I__593\ : Span4Mux_h
    port map (
            O => \N__8358\,
            I => \N__8352\
        );

    \I__592\ : Odrv12
    port map (
            O => \N__8355\,
            I => \TVP_VIDEO_c_5\
        );

    \I__591\ : Odrv4
    port map (
            O => \N__8352\,
            I => \TVP_VIDEO_c_5\
        );

    \I__590\ : InMux
    port map (
            O => \N__8347\,
            I => \N__8343\
        );

    \I__589\ : InMux
    port map (
            O => \N__8346\,
            I => \N__8340\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__8343\,
            I => \N__8337\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__8340\,
            I => \N__8332\
        );

    \I__586\ : Span4Mux_v
    port map (
            O => \N__8337\,
            I => \N__8329\
        );

    \I__585\ : InMux
    port map (
            O => \N__8336\,
            I => \N__8326\
        );

    \I__584\ : InMux
    port map (
            O => \N__8335\,
            I => \N__8322\
        );

    \I__583\ : Span4Mux_s1_v
    port map (
            O => \N__8332\,
            I => \N__8318\
        );

    \I__582\ : Span4Mux_v
    port map (
            O => \N__8329\,
            I => \N__8313\
        );

    \I__581\ : LocalMux
    port map (
            O => \N__8326\,
            I => \N__8313\
        );

    \I__580\ : InMux
    port map (
            O => \N__8325\,
            I => \N__8310\
        );

    \I__579\ : LocalMux
    port map (
            O => \N__8322\,
            I => \N__8307\
        );

    \I__578\ : InMux
    port map (
            O => \N__8321\,
            I => \N__8304\
        );

    \I__577\ : Span4Mux_h
    port map (
            O => \N__8318\,
            I => \N__8301\
        );

    \I__576\ : Span4Mux_v
    port map (
            O => \N__8313\,
            I => \N__8296\
        );

    \I__575\ : LocalMux
    port map (
            O => \N__8310\,
            I => \N__8296\
        );

    \I__574\ : Span4Mux_h
    port map (
            O => \N__8307\,
            I => \N__8293\
        );

    \I__573\ : LocalMux
    port map (
            O => \N__8304\,
            I => \N__8290\
        );

    \I__572\ : Span4Mux_v
    port map (
            O => \N__8301\,
            I => \N__8286\
        );

    \I__571\ : Span4Mux_v
    port map (
            O => \N__8296\,
            I => \N__8283\
        );

    \I__570\ : Span4Mux_h
    port map (
            O => \N__8293\,
            I => \N__8280\
        );

    \I__569\ : Span4Mux_h
    port map (
            O => \N__8290\,
            I => \N__8277\
        );

    \I__568\ : InMux
    port map (
            O => \N__8289\,
            I => \N__8274\
        );

    \I__567\ : Sp12to4
    port map (
            O => \N__8286\,
            I => \N__8271\
        );

    \I__566\ : Span4Mux_h
    port map (
            O => \N__8283\,
            I => \N__8268\
        );

    \I__565\ : Span4Mux_h
    port map (
            O => \N__8280\,
            I => \N__8265\
        );

    \I__564\ : Span4Mux_v
    port map (
            O => \N__8277\,
            I => \N__8262\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__8274\,
            I => \N__8259\
        );

    \I__562\ : Span12Mux_h
    port map (
            O => \N__8271\,
            I => \N__8255\
        );

    \I__561\ : Sp12to4
    port map (
            O => \N__8268\,
            I => \N__8252\
        );

    \I__560\ : Span4Mux_h
    port map (
            O => \N__8265\,
            I => \N__8245\
        );

    \I__559\ : Span4Mux_v
    port map (
            O => \N__8262\,
            I => \N__8245\
        );

    \I__558\ : Span4Mux_h
    port map (
            O => \N__8259\,
            I => \N__8245\
        );

    \I__557\ : InMux
    port map (
            O => \N__8258\,
            I => \N__8242\
        );

    \I__556\ : Span12Mux_v
    port map (
            O => \N__8255\,
            I => \N__8237\
        );

    \I__555\ : Span12Mux_h
    port map (
            O => \N__8252\,
            I => \N__8237\
        );

    \I__554\ : Span4Mux_v
    port map (
            O => \N__8245\,
            I => \N__8234\
        );

    \I__553\ : LocalMux
    port map (
            O => \N__8242\,
            I => \N__8231\
        );

    \I__552\ : Span12Mux_v
    port map (
            O => \N__8237\,
            I => \N__8228\
        );

    \I__551\ : Span4Mux_v
    port map (
            O => \N__8234\,
            I => \N__8225\
        );

    \I__550\ : Span4Mux_h
    port map (
            O => \N__8231\,
            I => \N__8222\
        );

    \I__549\ : Odrv12
    port map (
            O => \N__8228\,
            I => \TVP_VIDEO_c_4\
        );

    \I__548\ : Odrv4
    port map (
            O => \N__8225\,
            I => \TVP_VIDEO_c_4\
        );

    \I__547\ : Odrv4
    port map (
            O => \N__8222\,
            I => \TVP_VIDEO_c_4\
        );

    \I__546\ : InMux
    port map (
            O => \N__8215\,
            I => \N__8211\
        );

    \I__545\ : InMux
    port map (
            O => \N__8214\,
            I => \N__8208\
        );

    \I__544\ : LocalMux
    port map (
            O => \N__8211\,
            I => \N__8203\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__8208\,
            I => \N__8200\
        );

    \I__542\ : InMux
    port map (
            O => \N__8207\,
            I => \N__8197\
        );

    \I__541\ : InMux
    port map (
            O => \N__8206\,
            I => \N__8194\
        );

    \I__540\ : Sp12to4
    port map (
            O => \N__8203\,
            I => \N__8190\
        );

    \I__539\ : Span4Mux_h
    port map (
            O => \N__8200\,
            I => \N__8187\
        );

    \I__538\ : LocalMux
    port map (
            O => \N__8197\,
            I => \N__8184\
        );

    \I__537\ : LocalMux
    port map (
            O => \N__8194\,
            I => \N__8179\
        );

    \I__536\ : InMux
    port map (
            O => \N__8193\,
            I => \N__8176\
        );

    \I__535\ : Span12Mux_h
    port map (
            O => \N__8190\,
            I => \N__8172\
        );

    \I__534\ : Span4Mux_h
    port map (
            O => \N__8187\,
            I => \N__8169\
        );

    \I__533\ : Span4Mux_v
    port map (
            O => \N__8184\,
            I => \N__8166\
        );

    \I__532\ : InMux
    port map (
            O => \N__8183\,
            I => \N__8163\
        );

    \I__531\ : InMux
    port map (
            O => \N__8182\,
            I => \N__8160\
        );

    \I__530\ : Span12Mux_h
    port map (
            O => \N__8179\,
            I => \N__8157\
        );

    \I__529\ : LocalMux
    port map (
            O => \N__8176\,
            I => \N__8154\
        );

    \I__528\ : InMux
    port map (
            O => \N__8175\,
            I => \N__8151\
        );

    \I__527\ : Span12Mux_v
    port map (
            O => \N__8172\,
            I => \N__8146\
        );

    \I__526\ : Sp12to4
    port map (
            O => \N__8169\,
            I => \N__8146\
        );

    \I__525\ : Sp12to4
    port map (
            O => \N__8166\,
            I => \N__8143\
        );

    \I__524\ : LocalMux
    port map (
            O => \N__8163\,
            I => \N__8140\
        );

    \I__523\ : LocalMux
    port map (
            O => \N__8160\,
            I => \N__8137\
        );

    \I__522\ : Span12Mux_v
    port map (
            O => \N__8157\,
            I => \N__8130\
        );

    \I__521\ : Span12Mux_h
    port map (
            O => \N__8154\,
            I => \N__8130\
        );

    \I__520\ : LocalMux
    port map (
            O => \N__8151\,
            I => \N__8130\
        );

    \I__519\ : Span12Mux_v
    port map (
            O => \N__8146\,
            I => \N__8125\
        );

    \I__518\ : Span12Mux_h
    port map (
            O => \N__8143\,
            I => \N__8125\
        );

    \I__517\ : Span12Mux_h
    port map (
            O => \N__8140\,
            I => \N__8122\
        );

    \I__516\ : Span4Mux_h
    port map (
            O => \N__8137\,
            I => \N__8119\
        );

    \I__515\ : Span12Mux_h
    port map (
            O => \N__8130\,
            I => \N__8116\
        );

    \I__514\ : Span12Mux_h
    port map (
            O => \N__8125\,
            I => \N__8109\
        );

    \I__513\ : Span12Mux_v
    port map (
            O => \N__8122\,
            I => \N__8109\
        );

    \I__512\ : Sp12to4
    port map (
            O => \N__8119\,
            I => \N__8109\
        );

    \I__511\ : Odrv12
    port map (
            O => \N__8116\,
            I => \TVP_VIDEO_c_3\
        );

    \I__510\ : Odrv12
    port map (
            O => \N__8109\,
            I => \TVP_VIDEO_c_3\
        );

    \INVADV_R__i2C\ : INV
    port map (
            O => \INVADV_R__i2C_net\,
            I => \N__22547\
        );

    \INVdb5.NEXT_COUNTER__i3C\ : INV
    port map (
            O => \INVdb5.NEXT_COUNTER__i3C_net\,
            I => \N__19340\
        );

    \INVADV_R__i1C\ : INV
    port map (
            O => \INVADV_R__i1C_net\,
            I => \N__22535\
        );

    \IN_MUX_bfv_12_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_16_0_\
        );

    \IN_MUX_bfv_12_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \transmit_module.video_signal_controller.n3684\,
            carryinitout => \bfn_12_17_0_\
        );

    \IN_MUX_bfv_13_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_15_0_\
        );

    \IN_MUX_bfv_13_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \transmit_module.video_signal_controller.n3695\,
            carryinitout => \bfn_13_16_0_\
        );

    \IN_MUX_bfv_15_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_17_0_\
        );

    \IN_MUX_bfv_15_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \transmit_module.n3663\,
            carryinitout => \bfn_15_18_0_\
        );

    \IN_MUX_bfv_13_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_10_0_\
        );

    \IN_MUX_bfv_11_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_9_0_\
        );

    \IN_MUX_bfv_11_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \receive_module.rx_counter.n3718\,
            carryinitout => \bfn_11_10_0_\
        );

    \IN_MUX_bfv_10_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_9_0_\
        );

    \IN_MUX_bfv_10_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \receive_module.rx_counter.n3676\,
            carryinitout => \bfn_10_10_0_\
        );

    \IN_MUX_bfv_14_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_9_0_\
        );

    \IN_MUX_bfv_14_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \receive_module.rx_counter.n3727\,
            carryinitout => \bfn_14_10_0_\
        );

    \IN_MUX_bfv_15_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_8_0_\
        );

    \IN_MUX_bfv_13_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_11_0_\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \receive_module.rx_counter.i4_2_lut_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9444\,
            in2 => \_gnd_net_\,
            in3 => \N__9565\,
            lcout => OPEN,
            ltout => \receive_module.rx_counter.n12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.SYNC_45_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__8890\,
            in1 => \N__9594\,
            in2 => \N__8902\,
            in3 => \N__9310\,
            lcout => \DEBUG_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19342\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1_2_lut_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9488\,
            in2 => \_gnd_net_\,
            in3 => \N__9513\,
            lcout => \receive_module.rx_counter.n3938\,
            ltout => \receive_module.rx_counter.n3938_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i2_4_lut_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__9467\,
            in1 => \N__9442\,
            in2 => \N__8899\,
            in3 => \N__9202\,
            lcout => \receive_module.rx_counter.n3979\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i5_4_lut_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__8896\,
            in1 => \N__9537\,
            in2 => \N__9625\,
            in3 => \N__9468\,
            lcout => \receive_module.rx_counter.n13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1803_2_lut_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9620\,
            in2 => \_gnd_net_\,
            in3 => \N__9308\,
            lcout => OPEN,
            ltout => \receive_module.rx_counter.n3176_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1835_4_lut_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101000"
        )
    port map (
            in0 => \N__9536\,
            in1 => \N__9563\,
            in2 => \N__9205\,
            in3 => \N__9592\,
            lcout => \receive_module.rx_counter.n3208\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_2693_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000111000"
        )
    port map (
            in0 => \N__9196\,
            in1 => \N__23838\,
            in2 => \N__23613\,
            in3 => \N__9175\,
            lcout => OPEN,
            ltout => \line_buffer.n4170_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n4170_bdd_4_lut_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__23839\,
            in1 => \N__9166\,
            in2 => \N__9145\,
            in3 => \N__9142\,
            lcout => \line_buffer.n4173\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_2678_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__9127\,
            in1 => \N__23837\,
            in2 => \N__9109\,
            in3 => \N__23604\,
            lcout => \line_buffer.n4152\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2598_3_lut_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__23603\,
            in1 => \N__9094\,
            in2 => \_gnd_net_\,
            in3 => \N__9079\,
            lcout => \line_buffer.n4072\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n4152_bdd_4_lut_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011011000"
        )
    port map (
            in0 => \N__9073\,
            in1 => \N__9067\,
            in2 => \N__9046\,
            in3 => \N__23863\,
            lcout => OPEN,
            ltout => \line_buffer.n4155_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i2_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22846\,
            in2 => \N__9025\,
            in3 => \N__9022\,
            lcout => \TX_DATA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22650\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.Y_DELTA_PATTERN_i90_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9397\,
            lcout => \transmit_module.Y_DELTA_PATTERN_90\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22581\,
            ce => \N__16039\,
            sr => \N__21279\
        );

    \transmit_module.Y_DELTA_PATTERN_i94_LC_9_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9256\,
            lcout => \transmit_module.Y_DELTA_PATTERN_94\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22563\,
            ce => \N__16037\,
            sr => \N__21151\
        );

    \transmit_module.Y_DELTA_PATTERN_i95_LC_9_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9364\,
            lcout => \transmit_module.Y_DELTA_PATTERN_95\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22563\,
            ce => \N__16037\,
            sr => \N__21151\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_2668_LC_9_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__9250\,
            in1 => \N__23844\,
            in2 => \N__9238\,
            in3 => \N__23543\,
            lcout => \line_buffer.n4122\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.Y__i0_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9309\,
            in2 => \_gnd_net_\,
            in3 => \N__9223\,
            lcout => \receive_module.rx_counter.Y_0\,
            ltout => OPEN,
            carryin => \bfn_10_9_0_\,
            carryout => \receive_module.rx_counter.n3669\,
            clk => \N__19334\,
            ce => \N__11691\,
            sr => \N__9768\
        );

    \receive_module.rx_counter.Y__i1_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9621\,
            in2 => \_gnd_net_\,
            in3 => \N__9220\,
            lcout => \receive_module.rx_counter.Y_1\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3669\,
            carryout => \receive_module.rx_counter.n3670\,
            clk => \N__19334\,
            ce => \N__11691\,
            sr => \N__9768\
        );

    \receive_module.rx_counter.Y__i2_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9593\,
            in2 => \_gnd_net_\,
            in3 => \N__9217\,
            lcout => \receive_module.rx_counter.Y_2\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3670\,
            carryout => \receive_module.rx_counter.n3671\,
            clk => \N__19334\,
            ce => \N__11691\,
            sr => \N__9768\
        );

    \receive_module.rx_counter.Y__i3_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9564\,
            in2 => \_gnd_net_\,
            in3 => \N__9214\,
            lcout => \receive_module.rx_counter.Y_3\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3671\,
            carryout => \receive_module.rx_counter.n3672\,
            clk => \N__19334\,
            ce => \N__11691\,
            sr => \N__9768\
        );

    \receive_module.rx_counter.Y__i4_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9538\,
            in2 => \_gnd_net_\,
            in3 => \N__9211\,
            lcout => \receive_module.rx_counter.Y_4\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3672\,
            carryout => \receive_module.rx_counter.n3673\,
            clk => \N__19334\,
            ce => \N__11691\,
            sr => \N__9768\
        );

    \receive_module.rx_counter.Y__i5_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9514\,
            in2 => \_gnd_net_\,
            in3 => \N__9208\,
            lcout => \receive_module.rx_counter.Y_5\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3673\,
            carryout => \receive_module.rx_counter.n3674\,
            clk => \N__19334\,
            ce => \N__11691\,
            sr => \N__9768\
        );

    \receive_module.rx_counter.Y__i6_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9492\,
            in2 => \_gnd_net_\,
            in3 => \N__9283\,
            lcout => \receive_module.rx_counter.Y_6\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3674\,
            carryout => \receive_module.rx_counter.n3675\,
            clk => \N__19334\,
            ce => \N__11691\,
            sr => \N__9768\
        );

    \receive_module.rx_counter.Y__i7_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9469\,
            in2 => \_gnd_net_\,
            in3 => \N__9280\,
            lcout => \receive_module.rx_counter.Y_7\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3675\,
            carryout => \receive_module.rx_counter.n3676\,
            clk => \N__19334\,
            ce => \N__11691\,
            sr => \N__9768\
        );

    \receive_module.rx_counter.Y__i8_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9445\,
            in2 => \_gnd_net_\,
            in3 => \N__9277\,
            lcout => \receive_module.rx_counter.Y_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19338\,
            ce => \N__11692\,
            sr => \N__9772\
        );

    \transmit_module.Y_DELTA_PATTERN_i84_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9385\,
            lcout => \transmit_module.Y_DELTA_PATTERN_84\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22537\,
            ce => \N__16036\,
            sr => \N__21056\
        );

    \transmit_module.Y_DELTA_PATTERN_i83_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9274\,
            lcout => \transmit_module.Y_DELTA_PATTERN_83\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22537\,
            ce => \N__16036\,
            sr => \N__21056\
        );

    \transmit_module.Y_DELTA_PATTERN_i82_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__9268\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.Y_DELTA_PATTERN_82\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22649\,
            ce => \N__21457\,
            sr => \N__20955\
        );

    \transmit_module.Y_DELTA_PATTERN_i87_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9415\,
            lcout => \transmit_module.Y_DELTA_PATTERN_87\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22578\,
            ce => \N__16029\,
            sr => \N__21321\
        );

    \transmit_module.Y_DELTA_PATTERN_i92_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9370\,
            lcout => \transmit_module.Y_DELTA_PATTERN_92\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22578\,
            ce => \N__16029\,
            sr => \N__21321\
        );

    \transmit_module.Y_DELTA_PATTERN_i89_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9262\,
            lcout => \transmit_module.Y_DELTA_PATTERN_89\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22578\,
            ce => \N__16029\,
            sr => \N__21321\
        );

    \transmit_module.Y_DELTA_PATTERN_i88_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9421\,
            lcout => \transmit_module.Y_DELTA_PATTERN_88\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22578\,
            ce => \N__16029\,
            sr => \N__21321\
        );

    \transmit_module.Y_DELTA_PATTERN_i86_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9409\,
            lcout => \transmit_module.Y_DELTA_PATTERN_86\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22578\,
            ce => \N__16029\,
            sr => \N__21321\
        );

    \transmit_module.Y_DELTA_PATTERN_i91_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9403\,
            lcout => \transmit_module.Y_DELTA_PATTERN_91\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22578\,
            ce => \N__16029\,
            sr => \N__21321\
        );

    \transmit_module.Y_DELTA_PATTERN_i85_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9391\,
            lcout => \transmit_module.Y_DELTA_PATTERN_85\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22578\,
            ce => \N__16029\,
            sr => \N__21321\
        );

    \transmit_module.Y_DELTA_PATTERN_i93_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9376\,
            lcout => \transmit_module.Y_DELTA_PATTERN_93\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22564\,
            ce => \N__20596\,
            sr => \N__21251\
        );

    \transmit_module.Y_DELTA_PATTERN_i96_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9358\,
            lcout => \transmit_module.Y_DELTA_PATTERN_96\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22435\,
            ce => \N__21480\,
            sr => \N__21055\
        );

    \transmit_module.Y_DELTA_PATTERN_i97_LC_10_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9739\,
            lcout => \transmit_module.Y_DELTA_PATTERN_97\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22435\,
            ce => \N__21480\,
            sr => \N__21055\
        );

    \line_buffer.n4122_bdd_4_lut_LC_10_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__9352\,
            in1 => \N__9343\,
            in2 => \N__9337\,
            in3 => \N__23845\,
            lcout => \line_buffer.n4125\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.sub_23_add_2_2_lut_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9307\,
            in2 => \_gnd_net_\,
            in3 => \N__9286\,
            lcout => \receive_module.O_Y_0\,
            ltout => OPEN,
            carryin => \bfn_11_9_0_\,
            carryout => \receive_module.rx_counter.n3711\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.sub_23_add_2_3_lut_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9619\,
            in2 => \N__23307\,
            in3 => \N__9598\,
            lcout => \receive_module.O_Y_1\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3711\,
            carryout => \receive_module.rx_counter.n3712\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.sub_23_add_2_4_lut_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23252\,
            in2 => \N__9595\,
            in3 => \N__9568\,
            lcout => \receive_module.O_Y_2\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3712\,
            carryout => \receive_module.rx_counter.n3713\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.sub_23_add_2_5_lut_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9562\,
            in2 => \_gnd_net_\,
            in3 => \N__9541\,
            lcout => \receive_module.O_Y_3\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3713\,
            carryout => \receive_module.rx_counter.n3714\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.sub_23_add_2_6_lut_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9535\,
            in2 => \_gnd_net_\,
            in3 => \N__9517\,
            lcout => \receive_module.O_Y_4\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3714\,
            carryout => \receive_module.rx_counter.n3715\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.sub_23_add_2_7_lut_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9512\,
            in2 => \N__23308\,
            in3 => \N__9496\,
            lcout => \receive_module.O_Y_5\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3715\,
            carryout => \receive_module.rx_counter.n3716\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.sub_23_add_2_8_lut_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23256\,
            in2 => \N__9493\,
            in3 => \N__9472\,
            lcout => \receive_module.O_Y_6\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3716\,
            carryout => \receive_module.rx_counter.n3717\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.sub_23_add_2_9_lut_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9466\,
            in2 => \N__23309\,
            in3 => \N__9448\,
            lcout => \receive_module.O_Y_7\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3717\,
            carryout => \receive_module.rx_counter.n3718\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.sub_23_add_2_10_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9443\,
            in2 => \N__23306\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_10_0_\,
            carryout => \receive_module.rx_counter.O_VISIBLE_N_89\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i3_4_lut_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__10126\,
            in1 => \N__17386\,
            in2 => \N__9691\,
            in3 => \N__9679\,
            lcout => \DEBUG_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.SYNC_BUFF1_57_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9672\,
            lcout => \transmit_module.video_signal_controller.SYNC_BUFF1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22580\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.SYNC_BUFF2_58_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9643\,
            lcout => \transmit_module.video_signal_controller.SYNC_BUFF2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22580\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i3_4_lut_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__10560\,
            in1 => \N__10402\,
            in2 => \N__10527\,
            in3 => \N__10495\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n3987_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.VGA_VS_61_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10444\,
            in2 => \N__9637\,
            in3 => \N__10428\,
            lcout => \ADV_VSYNC_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22438\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_3_lut_4_lut_adj_17_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__10400\,
            in1 => \N__10516\,
            in2 => \N__10429\,
            in3 => \N__10555\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_4_lut_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__10350\,
            in1 => \N__9631\,
            in2 => \N__9634\,
            in3 => \N__10371\,
            lcout => \transmit_module.video_signal_controller.n3936\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_2_lut_3_lut_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111110"
        )
    port map (
            in0 => \N__10901\,
            in1 => \N__10349\,
            in2 => \N__10924\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.video_signal_controller.n6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_2_lut_rep_24_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10423\,
            in2 => \_gnd_net_\,
            in3 => \N__10399\,
            lcout => \transmit_module.video_signal_controller.n4215\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_2_lut_adj_12_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10623\,
            in2 => \_gnd_net_\,
            in3 => \N__10608\,
            lcout => \transmit_module.video_signal_controller.n3935\,
            ltout => \transmit_module.video_signal_controller.n3935_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i4_4_lut_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__10481\,
            in1 => \N__10370\,
            in2 => \N__9748\,
            in3 => \N__9745\,
            lcout => \transmit_module.video_signal_controller.n3892\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.Y_DELTA_PATTERN_i98_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19603\,
            lcout => \transmit_module.Y_DELTA_PATTERN_98\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22437\,
            ce => \N__16038\,
            sr => \N__21252\
        );

    \transmit_module.Y_DELTA_PATTERN_i76_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9697\,
            lcout => \transmit_module.Y_DELTA_PATTERN_76\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22437\,
            ce => \N__16038\,
            sr => \N__21252\
        );

    \transmit_module.Y_DELTA_PATTERN_i72_LC_11_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9727\,
            lcout => \transmit_module.Y_DELTA_PATTERN_72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22437\,
            ce => \N__16038\,
            sr => \N__21252\
        );

    \transmit_module.Y_DELTA_PATTERN_i75_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9733\,
            lcout => \transmit_module.Y_DELTA_PATTERN_75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22434\,
            ce => \N__21463\,
            sr => \N__21093\
        );

    \transmit_module.Y_DELTA_PATTERN_i73_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9703\,
            lcout => \transmit_module.Y_DELTA_PATTERN_73\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22434\,
            ce => \N__21463\,
            sr => \N__21093\
        );

    \transmit_module.Y_DELTA_PATTERN_i81_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9721\,
            lcout => \transmit_module.Y_DELTA_PATTERN_81\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22434\,
            ce => \N__21463\,
            sr => \N__21093\
        );

    \transmit_module.Y_DELTA_PATTERN_i74_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9709\,
            lcout => \transmit_module.Y_DELTA_PATTERN_74\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22434\,
            ce => \N__21463\,
            sr => \N__21093\
        );

    \transmit_module.Y_DELTA_PATTERN_i77_LC_11_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__10969\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.Y_DELTA_PATTERN_77\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22434\,
            ce => \N__21463\,
            sr => \N__21093\
        );

    \ADV_R__i1_LC_11_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22960\,
            lcout => n1996,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADV_R__i1C_net\,
            ce => 'H',
            sr => \N__14604\
        );

    \transmit_module.Y_DELTA_PATTERN_i63_LC_11_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10636\,
            lcout => \transmit_module.Y_DELTA_PATTERN_63\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22439\,
            ce => \N__21458\,
            sr => \N__21092\
        );

    \transmit_module.Y_DELTA_PATTERN_i70_LC_11_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9991\,
            lcout => \transmit_module.Y_DELTA_PATTERN_70\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22439\,
            ce => \N__21458\,
            sr => \N__21092\
        );

    \transmit_module.Y_DELTA_PATTERN_i69_LC_11_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10006\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.Y_DELTA_PATTERN_69\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22439\,
            ce => \N__21458\,
            sr => \N__21092\
        );

    \transmit_module.Y_DELTA_PATTERN_i71_LC_11_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10000\,
            lcout => \transmit_module.Y_DELTA_PATTERN_71\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22439\,
            ce => \N__21458\,
            sr => \N__21092\
        );

    \transmit_module.Y_DELTA_PATTERN_i62_LC_11_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9985\,
            lcout => \transmit_module.Y_DELTA_PATTERN_62\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22439\,
            ce => \N__21458\,
            sr => \N__21092\
        );

    \transmit_module.i1773_4_lut_LC_11_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__11713\,
            in1 => \N__11725\,
            in2 => \N__21335\,
            in3 => \N__20245\,
            lcout => n18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i29_1_lut_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__17110\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \receive_module.rx_counter.PULSE_1HZ_N_97\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.i667_3_lut_4_lut_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__12236\,
            in1 => \N__11987\,
            in2 => \N__12516\,
            in3 => \N__12545\,
            lcout => \receive_module.n5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.i1_2_lut_rep_21_3_lut_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__12512\,
            in1 => \N__11986\,
            in2 => \_gnd_net_\,
            in3 => \N__12237\,
            lcout => OPEN,
            ltout => \receive_module.n4212_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.i681_4_lut_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__13221\,
            in1 => \N__12963\,
            in2 => \N__10132\,
            in3 => \N__12547\,
            lcout => \receive_module.n3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.i1_2_lut_rep_22_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12506\,
            in2 => \_gnd_net_\,
            in3 => \N__12235\,
            lcout => OPEN,
            ltout => \receive_module.n4213_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.i674_3_lut_4_lut_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__13220\,
            in1 => \N__11988\,
            in2 => \N__10129\,
            in3 => \N__12546\,
            lcout => \receive_module.n4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.i660_3_lut_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__12544\,
            in1 => \N__12508\,
            in2 => \_gnd_net_\,
            in3 => \N__12234\,
            lcout => \receive_module.n6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.i652_2_lut_org_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__12507\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12543\,
            lcout => \receive_module.n7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1831_4_lut_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010001000"
        )
    port map (
            in0 => \N__17476\,
            in1 => \N__17503\,
            in2 => \N__12529\,
            in3 => \N__17416\,
            lcout => \receive_module.rx_counter.n3204\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1_2_lut_4_lut_adj_18_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__15760\,
            in1 => \N__15928\,
            in2 => \N__15807\,
            in3 => \N__15886\,
            lcout => n659,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \db5.i2_2_lut_rep_30_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__13426\,
            in1 => \_gnd_net_\,
            in2 => \N__13393\,
            in3 => \_gnd_net_\,
            lcout => \db5.n4221\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \db5.CLK_EN_13_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__13326\,
            in1 => \N__13388\,
            in2 => \N__13363\,
            in3 => \N__13425\,
            lcout => \DEBUG_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19335\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \db5.COUNTER_i2_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13389\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \db5.COUNTER_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19335\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1_2_lut_4_lut_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15759\,
            in1 => \N__15927\,
            in2 => \N__15806\,
            in3 => \N__15885\,
            lcout => n691,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \db5.COUNTER_i0_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13327\,
            lcout => \db5.COUNTER_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19335\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1_2_lut_3_lut_4_lut_adj_11_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__15887\,
            in1 => \N__15795\,
            in2 => \N__15931\,
            in3 => \N__15758\,
            lcout => \line_buffer.n626\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \db5.COUNTER_i1_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13356\,
            lcout => \db5.COUNTER_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19339\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1_3_lut_4_lut_adj_10_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__15929\,
            in1 => \N__15892\,
            in2 => \N__15848\,
            in3 => \N__15762\,
            lcout => \line_buffer.n561\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_2_lut_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13630\,
            in2 => \_gnd_net_\,
            in3 => \N__13603\,
            lcout => \transmit_module.video_signal_controller.n3917\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i3_4_lut_adj_14_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__13583\,
            in1 => \N__13559\,
            in2 => \N__13303\,
            in3 => \N__13604\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n3978_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i2578_3_lut_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10450\,
            in2 => \N__10135\,
            in3 => \N__13536\,
            lcout => \transmit_module.video_signal_controller.n4052\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_2_lut_rep_25_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__13560\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13537\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n4216_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.VGA_HS_60_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011101111"
        )
    port map (
            in0 => \N__13513\,
            in1 => \N__10333\,
            in2 => \N__10327\,
            in3 => \N__10324\,
            lcout => \ADV_HSYNC_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22620\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i570_3_lut_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__13605\,
            in1 => \N__13633\,
            in2 => \_gnd_net_\,
            in3 => \N__13584\,
            lcout => \transmit_module.video_signal_controller.n12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1859_4_lut_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001000"
        )
    port map (
            in0 => \N__13837\,
            in1 => \N__13811\,
            in2 => \N__10309\,
            in3 => \N__13784\,
            lcout => \transmit_module.video_signal_controller.n2274\,
            ltout => \transmit_module.video_signal_controller.n2274_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1227_2_lut_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10318\,
            in3 => \N__10315\,
            lcout => \transmit_module.video_signal_controller.n2594\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1853_4_lut_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100000000000"
        )
    port map (
            in0 => \N__10291\,
            in1 => \N__13294\,
            in2 => \N__10300\,
            in3 => \N__13508\,
            lcout => \transmit_module.video_signal_controller.n3226\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i560_2_lut_rep_26_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13654\,
            in2 => \_gnd_net_\,
            in3 => \N__13681\,
            lcout => \transmit_module.video_signal_controller.n4217\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_2_lut_3_lut_adj_15_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__13582\,
            in1 => \N__13558\,
            in2 => \_gnd_net_\,
            in3 => \N__13534\,
            lcout => \transmit_module.video_signal_controller.n2260\,
            ltout => \transmit_module.video_signal_controller.n2260_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i557_4_lut_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010100000"
        )
    port map (
            in0 => \N__13507\,
            in1 => \N__10290\,
            in2 => \N__10282\,
            in3 => \N__10279\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i2_4_lut_4_lut_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110110"
        )
    port map (
            in0 => \N__13835\,
            in1 => \N__13807\,
            in2 => \N__10453\,
            in3 => \N__13783\,
            lcout => \transmit_module.n3910\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i2_3_lut_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__13785\,
            in1 => \_gnd_net_\,
            in2 => \N__13813\,
            in3 => \N__13836\,
            lcout => \transmit_module.video_signal_controller.n2219\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.VGA_Y_i0_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10443\,
            in2 => \_gnd_net_\,
            in3 => \N__10432\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_0\,
            ltout => OPEN,
            carryin => \bfn_12_16_0_\,
            carryout => \transmit_module.video_signal_controller.n3677\,
            clk => \N__22561\,
            ce => \N__13761\,
            sr => \N__10584\
        );

    \transmit_module.video_signal_controller.VGA_Y_i1_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10427\,
            in2 => \_gnd_net_\,
            in3 => \N__10405\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_1\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3677\,
            carryout => \transmit_module.video_signal_controller.n3678\,
            clk => \N__22561\,
            ce => \N__13761\,
            sr => \N__10584\
        );

    \transmit_module.video_signal_controller.VGA_Y_i2_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10401\,
            in2 => \_gnd_net_\,
            in3 => \N__10381\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_2\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3678\,
            carryout => \transmit_module.video_signal_controller.n3679\,
            clk => \N__22561\,
            ce => \N__13761\,
            sr => \N__10584\
        );

    \transmit_module.video_signal_controller.VGA_Y_i3_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10559\,
            in2 => \_gnd_net_\,
            in3 => \N__10378\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_3\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3679\,
            carryout => \transmit_module.video_signal_controller.n3680\,
            clk => \N__22561\,
            ce => \N__13761\,
            sr => \N__10584\
        );

    \transmit_module.video_signal_controller.VGA_Y_i4_LC_12_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10520\,
            in2 => \_gnd_net_\,
            in3 => \N__10375\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_4\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3680\,
            carryout => \transmit_module.video_signal_controller.n3681\,
            clk => \N__22561\,
            ce => \N__13761\,
            sr => \N__10584\
        );

    \transmit_module.video_signal_controller.VGA_Y_i5_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10372\,
            in2 => \_gnd_net_\,
            in3 => \N__10354\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_5\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3681\,
            carryout => \transmit_module.video_signal_controller.n3682\,
            clk => \N__22561\,
            ce => \N__13761\,
            sr => \N__10584\
        );

    \transmit_module.video_signal_controller.VGA_Y_i6_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10351\,
            in2 => \_gnd_net_\,
            in3 => \N__10336\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_6\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3682\,
            carryout => \transmit_module.video_signal_controller.n3683\,
            clk => \N__22561\,
            ce => \N__13761\,
            sr => \N__10584\
        );

    \transmit_module.video_signal_controller.VGA_Y_i7_LC_12_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10624\,
            in2 => \_gnd_net_\,
            in3 => \N__10612\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_7\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3683\,
            carryout => \transmit_module.video_signal_controller.n3684\,
            clk => \N__22561\,
            ce => \N__13761\,
            sr => \N__10584\
        );

    \transmit_module.video_signal_controller.VGA_Y_i8_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10609\,
            in2 => \_gnd_net_\,
            in3 => \N__10597\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_8\,
            ltout => OPEN,
            carryin => \bfn_12_17_0_\,
            carryout => \transmit_module.video_signal_controller.n3685\,
            clk => \N__22499\,
            ce => \N__13768\,
            sr => \N__10585\
        );

    \transmit_module.video_signal_controller.VGA_Y_i9_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10483\,
            in2 => \_gnd_net_\,
            in3 => \N__10594\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_9\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3685\,
            carryout => \transmit_module.video_signal_controller.n3686\,
            clk => \N__22499\,
            ce => \N__13768\,
            sr => \N__10585\
        );

    \transmit_module.video_signal_controller.VGA_Y_i10_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10903\,
            in2 => \_gnd_net_\,
            in3 => \N__10591\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_10\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3686\,
            carryout => \transmit_module.video_signal_controller.n3687\,
            clk => \N__22499\,
            ce => \N__13768\,
            sr => \N__10585\
        );

    \transmit_module.video_signal_controller.VGA_Y_i11_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10923\,
            in2 => \_gnd_net_\,
            in3 => \N__10588\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22499\,
            ce => \N__13768\,
            sr => \N__10585\
        );

    \transmit_module.video_signal_controller.i1_4_lut_adj_13_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111100000"
        )
    port map (
            in0 => \N__10561\,
            in1 => \N__10534\,
            in2 => \N__10528\,
            in3 => \N__10494\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.VGA_VISIBLE_Y_N_553_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i2_4_lut_adj_16_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000001010000"
        )
    port map (
            in0 => \N__10885\,
            in1 => \N__10482\,
            in2 => \N__10465\,
            in3 => \N__10462\,
            lcout => \transmit_module.n3926\,
            ltout => \transmit_module.n3926_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.mux_14_i3_3_lut_4_lut_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110011001100"
        )
    port map (
            in0 => \N__17797\,
            in1 => \N__17822\,
            in2 => \N__10456\,
            in3 => \N__19100\,
            lcout => \transmit_module.n217\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_2_lut_rep_27_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10922\,
            in2 => \_gnd_net_\,
            in3 => \N__10902\,
            lcout => \transmit_module.video_signal_controller.n4218\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1211_1_lut_2_lut_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19095\,
            in2 => \_gnd_net_\,
            in3 => \N__19467\,
            lcout => n2587,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.mux_14_i1_3_lut_4_lut_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__18420\,
            in1 => \N__19099\,
            in2 => \N__17521\,
            in3 => \N__19468\,
            lcout => \transmit_module.n219\,
            ltout => \transmit_module.n219_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1757_4_lut_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__20167\,
            in1 => \N__21036\,
            in2 => \N__10879\,
            in3 => \N__17839\,
            lcout => n28,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_2_lut_rep_19_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__19469\,
            in1 => \_gnd_net_\,
            in2 => \N__19121\,
            in3 => \_gnd_net_\,
            lcout => n4210,
            ltout => \n4210_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1762_4_lut_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111100"
        )
    port map (
            in0 => \N__19716\,
            in1 => \N__21037\,
            in2 => \N__10639\,
            in3 => \N__20166\,
            lcout => \transmit_module.n2277\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i13_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__22793\,
            in1 => \N__19150\,
            in2 => \_gnd_net_\,
            in3 => \N__19397\,
            lcout => \DEBUG_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22534\,
            ce => 'H',
            sr => \N__21167\
        );

    \transmit_module.Y_DELTA_PATTERN_i64_LC_12_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10948\,
            lcout => \transmit_module.Y_DELTA_PATTERN_64\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22348\,
            ce => \N__21456\,
            sr => \N__21306\
        );

    \transmit_module.Y_DELTA_PATTERN_i66_LC_12_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10630\,
            lcout => \transmit_module.Y_DELTA_PATTERN_66\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22348\,
            ce => \N__21456\,
            sr => \N__21306\
        );

    \transmit_module.Y_DELTA_PATTERN_i67_LC_12_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10975\,
            lcout => \transmit_module.Y_DELTA_PATTERN_67\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22348\,
            ce => \N__21456\,
            sr => \N__21306\
        );

    \transmit_module.Y_DELTA_PATTERN_i80_LC_12_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10993\,
            lcout => \transmit_module.Y_DELTA_PATTERN_80\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22348\,
            ce => \N__21456\,
            sr => \N__21306\
        );

    \transmit_module.Y_DELTA_PATTERN_i68_LC_12_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__10981\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.Y_DELTA_PATTERN_68\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22348\,
            ce => \N__21456\,
            sr => \N__21306\
        );

    \transmit_module.Y_DELTA_PATTERN_i78_LC_12_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10936\,
            lcout => \transmit_module.Y_DELTA_PATTERN_78\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22315\,
            ce => \N__21489\,
            sr => \N__21278\
        );

    \transmit_module.Y_DELTA_PATTERN_i61_LC_12_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10960\,
            lcout => \transmit_module.Y_DELTA_PATTERN_61\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22315\,
            ce => \N__21489\,
            sr => \N__21278\
        );

    \transmit_module.Y_DELTA_PATTERN_i51_LC_12_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14545\,
            lcout => \transmit_module.Y_DELTA_PATTERN_51\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22315\,
            ce => \N__21489\,
            sr => \N__21278\
        );

    \transmit_module.Y_DELTA_PATTERN_i65_LC_12_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10954\,
            lcout => \transmit_module.Y_DELTA_PATTERN_65\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22315\,
            ce => \N__21489\,
            sr => \N__21278\
        );

    \transmit_module.Y_DELTA_PATTERN_i79_LC_12_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10942\,
            lcout => \transmit_module.Y_DELTA_PATTERN_79\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22315\,
            ce => \N__21489\,
            sr => \N__21278\
        );

    \transmit_module.Y_DELTA_PATTERN_i56_LC_12_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10930\,
            lcout => \transmit_module.Y_DELTA_PATTERN_56\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21958\,
            ce => \N__21493\,
            sr => \N__21288\
        );

    \transmit_module.Y_DELTA_PATTERN_i57_LC_12_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14656\,
            lcout => \transmit_module.Y_DELTA_PATTERN_57\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__21958\,
            ce => \N__21493\,
            sr => \N__21288\
        );

    \transmit_module.ADDR_Y_COMPONENT__i10_LC_12_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17951\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22230\,
            ce => \N__19881\,
            sr => \N__21325\
        );

    \transmit_module.mux_12_i11_3_lut_LC_12_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__19717\,
            in1 => \N__11731\,
            in2 => \_gnd_net_\,
            in3 => \N__17944\,
            lcout => \transmit_module.n178\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.mux_14_i11_3_lut_4_lut_LC_12_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__17920\,
            in1 => \N__19129\,
            in2 => \N__17955\,
            in3 => \N__19520\,
            lcout => \transmit_module.n209\,
            ltout => \transmit_module.n209_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i10_LC_12_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__11709\,
            in1 => \N__21268\,
            in2 => \N__11695\,
            in3 => \N__20239\,
            lcout => \transmit_module.TX_ADDR_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22229\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i284_3_lut_3_lut_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101010101"
        )
    port map (
            in0 => \N__17106\,
            in1 => \N__15441\,
            in2 => \_gnd_net_\,
            in3 => \N__11668\,
            lcout => n2283,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.old_HS_50_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15442\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \old_HS\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19329\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.sub_29_add_2_2_lut_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17026\,
            in2 => \_gnd_net_\,
            in3 => \N__11434\,
            lcout => \RX_ADDR_3\,
            ltout => OPEN,
            carryin => \bfn_13_10_0_\,
            carryout => \receive_module.rx_counter.n3650\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.sub_29_add_2_3_lut_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17047\,
            in2 => \N__23303\,
            in3 => \N__11212\,
            lcout => \RX_ADDR_4\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3650\,
            carryout => \receive_module.rx_counter.n3651\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.sub_29_add_2_4_lut_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23238\,
            in2 => \N__17074\,
            in3 => \N__10996\,
            lcout => \RX_ADDR_5\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3651\,
            carryout => \receive_module.rx_counter.n3652\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.sub_29_add_2_5_lut_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17407\,
            in2 => \N__23304\,
            in3 => \N__12559\,
            lcout => \receive_module.O_X_6\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3652\,
            carryout => \receive_module.rx_counter.n3653\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.sub_29_add_2_6_lut_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17437\,
            in2 => \_gnd_net_\,
            in3 => \N__12556\,
            lcout => \receive_module.O_X_7\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3653\,
            carryout => \receive_module.rx_counter.n3654\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.sub_29_add_2_7_lut_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17497\,
            in2 => \N__23305\,
            in3 => \N__12553\,
            lcout => \receive_module.O_X_8\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3654\,
            carryout => \receive_module.rx_counter.n3655\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.sub_29_add_2_8_lut_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__17470\,
            in1 => \N__23245\,
            in2 => \_gnd_net_\,
            in3 => \N__12550\,
            lcout => \receive_module.O_X_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1_2_lut_4_lut_adj_19_LC_13_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__17027\,
            in1 => \N__17071\,
            in2 => \N__17443\,
            in3 => \N__17048\,
            lcout => \receive_module.rx_counter.n4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_629_2_lut_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12520\,
            in2 => \N__12484\,
            in3 => \_gnd_net_\,
            lcout => \RX_ADDR_6\,
            ltout => OPEN,
            carryin => \bfn_13_11_0_\,
            carryout => \receive_module.n3699\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_629_3_lut_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12250\,
            in2 => \N__12244\,
            in3 => \N__11998\,
            lcout => \RX_ADDR_7\,
            ltout => OPEN,
            carryin => \receive_module.n3699\,
            carryout => \receive_module.n3700\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_629_4_lut_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11995\,
            in2 => \N__11968\,
            in3 => \N__11734\,
            lcout => \RX_ADDR_8\,
            ltout => OPEN,
            carryin => \receive_module.n3700\,
            carryout => \receive_module.n3701\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_629_5_lut_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13237\,
            in2 => \N__13231\,
            in3 => \N__12982\,
            lcout => \RX_ADDR_9\,
            ltout => OPEN,
            carryin => \receive_module.n3701\,
            carryout => \receive_module.n3702\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_629_6_lut_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12979\,
            in2 => \N__12973\,
            in3 => \N__12730\,
            lcout => \RX_ADDR_10\,
            ltout => OPEN,
            carryin => \receive_module.n3702\,
            carryout => \receive_module.n3703\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_629_7_lut_LC_13_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12727\,
            in2 => \N__12721\,
            in3 => \N__12706\,
            lcout => \RX_ADDR_11\,
            ltout => OPEN,
            carryin => \receive_module.n3703\,
            carryout => \receive_module.n3704\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_629_8_lut_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12703\,
            in2 => \N__12697\,
            in3 => \N__12682\,
            lcout => \RX_ADDR_12\,
            ltout => OPEN,
            carryin => \receive_module.n3704\,
            carryout => \receive_module.n3705\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_629_9_lut_LC_13_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__12679\,
            in1 => \N__12673\,
            in2 => \_gnd_net_\,
            in3 => \N__12661\,
            lcout => \DEBUG_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1_2_lut_3_lut_4_lut_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__15923\,
            in1 => \N__15889\,
            in2 => \N__15843\,
            in3 => \N__15755\,
            lcout => \line_buffer.n627\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1_3_lut_4_lut_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__15922\,
            in1 => \N__15890\,
            in2 => \N__15844\,
            in3 => \N__15756\,
            lcout => \line_buffer.n562\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \db5.COUNTER_i3_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13424\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \db5.COUNTER_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19336\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1_2_lut_4_lut_adj_22_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__15921\,
            in1 => \N__15888\,
            in2 => \N__15842\,
            in3 => \N__15757\,
            lcout => n690,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \db5.NEXT_COUNTER__i3_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__13345\,
            in1 => \N__13408\,
            in2 => \N__13435\,
            in3 => \N__13375\,
            lcout => \db5.NEXT_COUNTER_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVdb5.NEXT_COUNTER__i3C_net\,
            ce => 'H',
            sr => \N__13315\
        );

    \db5.NEXT_COUNTER__i2_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__13374\,
            in1 => \N__13407\,
            in2 => \_gnd_net_\,
            in3 => \N__13344\,
            lcout => \db5.NEXT_COUNTER_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVdb5.NEXT_COUNTER__i3C_net\,
            ce => 'H',
            sr => \N__13315\
        );

    \db5.NEXT_COUNTER__i1_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__13343\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13373\,
            lcout => \db5.NEXT_COUNTER_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVdb5.NEXT_COUNTER__i3C_net\,
            ce => 'H',
            sr => \N__13315\
        );

    \db5.NEXT_COUNTER__i0_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13342\,
            lcout => \db5.NEXT_COUNTER_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVdb5.NEXT_COUNTER__i3C_net\,
            ce => 'H',
            sr => \N__13315\
        );

    \transmit_module.video_signal_controller.i2_4_lut_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010000000"
        )
    port map (
            in0 => \N__13683\,
            in1 => \N__13631\,
            in2 => \N__13660\,
            in3 => \N__13254\,
            lcout => \transmit_module.video_signal_controller.n3997\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1823_2_lut_3_lut_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__13253\,
            in1 => \N__13655\,
            in2 => \_gnd_net_\,
            in3 => \N__13682\,
            lcout => \transmit_module.video_signal_controller.n3196\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2628_3_lut_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__13288\,
            in1 => \N__13270\,
            in2 => \_gnd_net_\,
            in3 => \N__23591\,
            lcout => \line_buffer.n4102\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.VGA_X_i0_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13255\,
            in2 => \_gnd_net_\,
            in3 => \N__13240\,
            lcout => \transmit_module.video_signal_controller.VGA_X_0\,
            ltout => OPEN,
            carryin => \bfn_13_15_0_\,
            carryout => \transmit_module.video_signal_controller.n3688\,
            clk => \N__22422\,
            ce => 'H',
            sr => \N__13753\
        );

    \transmit_module.video_signal_controller.VGA_X_i1_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13684\,
            in2 => \_gnd_net_\,
            in3 => \N__13663\,
            lcout => \transmit_module.video_signal_controller.VGA_X_1\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3688\,
            carryout => \transmit_module.video_signal_controller.n3689\,
            clk => \N__22422\,
            ce => 'H',
            sr => \N__13753\
        );

    \transmit_module.video_signal_controller.VGA_X_i2_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13659\,
            in2 => \_gnd_net_\,
            in3 => \N__13636\,
            lcout => \transmit_module.video_signal_controller.VGA_X_2\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3689\,
            carryout => \transmit_module.video_signal_controller.n3690\,
            clk => \N__22422\,
            ce => 'H',
            sr => \N__13753\
        );

    \transmit_module.video_signal_controller.VGA_X_i3_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13632\,
            in2 => \_gnd_net_\,
            in3 => \N__13609\,
            lcout => \transmit_module.video_signal_controller.VGA_X_3\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3690\,
            carryout => \transmit_module.video_signal_controller.n3691\,
            clk => \N__22422\,
            ce => 'H',
            sr => \N__13753\
        );

    \transmit_module.video_signal_controller.VGA_X_i4_LC_13_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13606\,
            in2 => \_gnd_net_\,
            in3 => \N__13588\,
            lcout => \transmit_module.video_signal_controller.VGA_X_4\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3691\,
            carryout => \transmit_module.video_signal_controller.n3692\,
            clk => \N__22422\,
            ce => 'H',
            sr => \N__13753\
        );

    \transmit_module.video_signal_controller.VGA_X_i5_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13585\,
            in2 => \_gnd_net_\,
            in3 => \N__13564\,
            lcout => \transmit_module.video_signal_controller.VGA_X_5\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3692\,
            carryout => \transmit_module.video_signal_controller.n3693\,
            clk => \N__22422\,
            ce => 'H',
            sr => \N__13753\
        );

    \transmit_module.video_signal_controller.VGA_X_i6_LC_13_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13561\,
            in2 => \_gnd_net_\,
            in3 => \N__13540\,
            lcout => \transmit_module.video_signal_controller.VGA_X_6\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3693\,
            carryout => \transmit_module.video_signal_controller.n3694\,
            clk => \N__22422\,
            ce => 'H',
            sr => \N__13753\
        );

    \transmit_module.video_signal_controller.VGA_X_i7_LC_13_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13535\,
            in2 => \_gnd_net_\,
            in3 => \N__13516\,
            lcout => \transmit_module.video_signal_controller.VGA_X_7\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3694\,
            carryout => \transmit_module.video_signal_controller.n3695\,
            clk => \N__22422\,
            ce => 'H',
            sr => \N__13753\
        );

    \transmit_module.video_signal_controller.VGA_X_i8_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13509\,
            in2 => \_gnd_net_\,
            in3 => \N__13489\,
            lcout => \transmit_module.video_signal_controller.VGA_X_8\,
            ltout => OPEN,
            carryin => \bfn_13_16_0_\,
            carryout => \transmit_module.video_signal_controller.n3696\,
            clk => \N__22609\,
            ce => 'H',
            sr => \N__13754\
        );

    \transmit_module.video_signal_controller.VGA_X_i9_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13834\,
            in2 => \_gnd_net_\,
            in3 => \N__13816\,
            lcout => \transmit_module.video_signal_controller.VGA_X_9\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3696\,
            carryout => \transmit_module.video_signal_controller.n3697\,
            clk => \N__22609\,
            ce => 'H',
            sr => \N__13754\
        );

    \transmit_module.video_signal_controller.VGA_X_i10_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13812\,
            in2 => \_gnd_net_\,
            in3 => \N__13792\,
            lcout => \transmit_module.video_signal_controller.VGA_X_10\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3697\,
            carryout => \transmit_module.video_signal_controller.n3698\,
            clk => \N__22609\,
            ce => 'H',
            sr => \N__13754\
        );

    \transmit_module.video_signal_controller.VGA_X_i11_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13786\,
            in2 => \_gnd_net_\,
            in3 => \N__13789\,
            lcout => \transmit_module.video_signal_controller.VGA_X_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22609\,
            ce => 'H',
            sr => \N__13754\
        );

    \transmit_module.video_signal_controller.mux_14_i7_3_lut_4_lut_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__17725\,
            in1 => \N__19101\,
            in2 => \N__17756\,
            in3 => \N__19500\,
            lcout => \transmit_module.n213\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i2_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__14122\,
            in1 => \N__14107\,
            in2 => \N__21259\,
            in3 => \N__20215\,
            lcout => \transmit_module.TX_ADDR_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22533\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i6_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__13726\,
            in1 => \N__22829\,
            in2 => \N__15670\,
            in3 => \N__16051\,
            lcout => \TX_DATA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22533\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i143_2_lut_3_lut_4_lut_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__19501\,
            in1 => \N__16762\,
            in2 => \N__21219\,
            in3 => \N__16705\,
            lcout => \transmit_module.n2361\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_2703_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__13717\,
            in1 => \N__23807\,
            in2 => \N__13702\,
            in3 => \N__23576\,
            lcout => \line_buffer.n4182\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.mux_14_i9_3_lut_4_lut_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__17668\,
            in1 => \N__19103\,
            in2 => \N__17893\,
            in3 => \N__19494\,
            lcout => \transmit_module.n211\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.mux_14_i8_3_lut_4_lut_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__19493\,
            in1 => \N__17683\,
            in2 => \N__17712\,
            in3 => \N__19104\,
            lcout => \transmit_module.n212\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i3_3_lut_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__19714\,
            in1 => \N__16366\,
            in2 => \_gnd_net_\,
            in3 => \N__17821\,
            lcout => \transmit_module.n186\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_3_lut_4_lut_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__19496\,
            in1 => \N__19715\,
            in2 => \N__21196\,
            in3 => \N__19572\,
            lcout => \transmit_module.n2305\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.mux_14_i10_3_lut_4_lut_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011110000"
        )
    port map (
            in0 => \N__17653\,
            in1 => \N__19102\,
            in2 => \N__18465\,
            in3 => \N__19492\,
            lcout => \transmit_module.n210\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i143_2_lut_3_lut_4_lut_rep_34_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__19495\,
            in1 => \N__16761\,
            in2 => \N__21195\,
            in3 => \N__16717\,
            lcout => \transmit_module.n4225\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i9_3_lut_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__17886\,
            in1 => \N__19692\,
            in2 => \_gnd_net_\,
            in3 => \N__17866\,
            lcout => \transmit_module.n180\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_2_lut_rep_20_3_lut_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__16712\,
            in1 => \N__16756\,
            in2 => \_gnd_net_\,
            in3 => \N__19470\,
            lcout => \transmit_module.n4211\,
            ltout => \transmit_module.n4211_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1765_4_lut_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__21035\,
            in1 => \N__14121\,
            in2 => \N__14110\,
            in3 => \N__14106\,
            lcout => n26,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.mux_14_i4_3_lut_4_lut_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__18375\,
            in1 => \N__19122\,
            in2 => \N__17782\,
            in3 => \N__19471\,
            lcout => \transmit_module.n216\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n4182_bdd_4_lut_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__13876\,
            in1 => \N__13861\,
            in2 => \N__13852\,
            in3 => \N__23855\,
            lcout => OPEN,
            ltout => \line_buffer.n4185_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i7_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22764\,
            in2 => \N__14539\,
            in3 => \N__14536\,
            lcout => \TX_DATA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22266\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.old_VGA_HS_34_LC_13_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16713\,
            lcout => \transmit_module.old_VGA_HS\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22266\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADV_R__i2_LC_13_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20404\,
            lcout => n1995,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADV_R__i2C_net\,
            ce => 'H',
            sr => \N__14605\
        );

    \ADV_R__i3_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14479\,
            lcout => n1994,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADV_R__i2C_net\,
            ce => 'H',
            sr => \N__14605\
        );

    \ADV_R__i4_LC_13_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21580\,
            lcout => n1993,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADV_R__i2C_net\,
            ce => 'H',
            sr => \N__14605\
        );

    \ADV_R__i5_LC_13_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22708\,
            lcout => n1992,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADV_R__i2C_net\,
            ce => 'H',
            sr => \N__14605\
        );

    \ADV_R__i6_LC_13_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17971\,
            lcout => n1991,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADV_R__i2C_net\,
            ce => 'H',
            sr => \N__14605\
        );

    \ADV_R__i7_LC_13_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__14254\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n1990,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADV_R__i2C_net\,
            ce => 'H',
            sr => \N__14605\
        );

    \ADV_R__i8_LC_13_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14188\,
            lcout => \ADV_B_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADV_R__i2C_net\,
            ce => 'H',
            sr => \N__14605\
        );

    \transmit_module.Y_DELTA_PATTERN_i42_LC_13_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14587\,
            lcout => \transmit_module.Y_DELTA_PATTERN_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22486\,
            ce => \N__21436\,
            sr => \N__21344\
        );

    \transmit_module.Y_DELTA_PATTERN_i43_LC_13_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14581\,
            lcout => \transmit_module.Y_DELTA_PATTERN_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22486\,
            ce => \N__21436\,
            sr => \N__21344\
        );

    \transmit_module.Y_DELTA_PATTERN_i46_LC_13_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14563\,
            lcout => \transmit_module.Y_DELTA_PATTERN_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22486\,
            ce => \N__21436\,
            sr => \N__21344\
        );

    \transmit_module.Y_DELTA_PATTERN_i44_LC_13_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14569\,
            lcout => \transmit_module.Y_DELTA_PATTERN_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22486\,
            ce => \N__21436\,
            sr => \N__21344\
        );

    \transmit_module.Y_DELTA_PATTERN_i45_LC_13_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14575\,
            lcout => \transmit_module.Y_DELTA_PATTERN_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22486\,
            ce => \N__21436\,
            sr => \N__21344\
        );

    \transmit_module.Y_DELTA_PATTERN_i47_LC_13_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14557\,
            lcout => \transmit_module.Y_DELTA_PATTERN_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22486\,
            ce => \N__21436\,
            sr => \N__21344\
        );

    \transmit_module.Y_DELTA_PATTERN_i53_LC_13_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14692\,
            lcout => \transmit_module.Y_DELTA_PATTERN_53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22322\,
            ce => \N__21464\,
            sr => \N__21166\
        );

    \transmit_module.Y_DELTA_PATTERN_i48_LC_13_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14698\,
            lcout => \transmit_module.Y_DELTA_PATTERN_48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22322\,
            ce => \N__21464\,
            sr => \N__21166\
        );

    \transmit_module.Y_DELTA_PATTERN_i52_LC_13_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14551\,
            lcout => \transmit_module.Y_DELTA_PATTERN_52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22322\,
            ce => \N__21464\,
            sr => \N__21166\
        );

    \transmit_module.Y_DELTA_PATTERN_i49_LC_13_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14680\,
            lcout => \transmit_module.Y_DELTA_PATTERN_49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22322\,
            ce => \N__21464\,
            sr => \N__21166\
        );

    \transmit_module.Y_DELTA_PATTERN_i54_LC_13_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__14668\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.Y_DELTA_PATTERN_54\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22322\,
            ce => \N__21464\,
            sr => \N__21166\
        );

    \transmit_module.Y_DELTA_PATTERN_i50_LC_13_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14686\,
            lcout => \transmit_module.Y_DELTA_PATTERN_50\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22322\,
            ce => \N__21464\,
            sr => \N__21166\
        );

    \transmit_module.Y_DELTA_PATTERN_i59_LC_13_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14644\,
            lcout => \transmit_module.Y_DELTA_PATTERN_59\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22409\,
            ce => \N__21437\,
            sr => \N__21345\
        );

    \transmit_module.Y_DELTA_PATTERN_i55_LC_13_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14674\,
            lcout => \transmit_module.Y_DELTA_PATTERN_55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22409\,
            ce => \N__21437\,
            sr => \N__21345\
        );

    \transmit_module.Y_DELTA_PATTERN_i58_LC_13_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14662\,
            lcout => \transmit_module.Y_DELTA_PATTERN_58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22409\,
            ce => \N__21437\,
            sr => \N__21345\
        );

    \transmit_module.Y_DELTA_PATTERN_i60_LC_13_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14650\,
            lcout => \transmit_module.Y_DELTA_PATTERN_60\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22409\,
            ce => \N__21437\,
            sr => \N__21345\
        );

    \transmit_module.ADDR_Y_COMPONENT__i6_LC_13_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17758\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22282\,
            ce => \N__19882\,
            sr => \N__21269\
        );

    \line_buffer.i2627_3_lut_LC_13_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__14638\,
            in1 => \N__14620\,
            in2 => \_gnd_net_\,
            in3 => \N__23553\,
            lcout => \line_buffer.n4101\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1769_4_lut_LC_13_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__16414\,
            in1 => \N__16345\,
            in2 => \N__21346\,
            in3 => \N__20241\,
            lcout => n22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1_2_lut_adj_25_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17157\,
            in2 => \_gnd_net_\,
            in3 => \N__17187\,
            lcout => OPEN,
            ltout => \receive_module.rx_counter.n5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i3_4_lut_adj_26_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111111111"
        )
    port map (
            in0 => \N__16392\,
            in1 => \N__17139\,
            in2 => \N__15445\,
            in3 => \N__15403\,
            lcout => \receive_module.rx_counter.n11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i28_1_lut_rep_23_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15440\,
            lcout => n4214,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1_2_lut_adj_24_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16377\,
            in2 => \_gnd_net_\,
            in3 => \N__17172\,
            lcout => \receive_module.rx_counter.n4_adj_576\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.X_277__i1_LC_14_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15185\,
            in2 => \_gnd_net_\,
            in3 => \N__15166\,
            lcout => \RX_ADDR_0\,
            ltout => OPEN,
            carryin => \bfn_14_9_0_\,
            carryout => \receive_module.rx_counter.n3720\,
            clk => \N__19326\,
            ce => 'H',
            sr => \N__15952\
        );

    \receive_module.rx_counter.X_277__i2_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14954\,
            in2 => \_gnd_net_\,
            in3 => \N__14932\,
            lcout => \RX_ADDR_1\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3720\,
            carryout => \receive_module.rx_counter.n3721\,
            clk => \N__19326\,
            ce => 'H',
            sr => \N__15952\
        );

    \receive_module.rx_counter.X_277__i3_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14723\,
            in2 => \_gnd_net_\,
            in3 => \N__14701\,
            lcout => \RX_ADDR_2\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3721\,
            carryout => \receive_module.rx_counter.n3722\,
            clk => \N__19326\,
            ce => 'H',
            sr => \N__15952\
        );

    \receive_module.rx_counter.X_277__i4_LC_14_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17029\,
            in2 => \_gnd_net_\,
            in3 => \N__15973\,
            lcout => \receive_module.rx_counter.X_3\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3722\,
            carryout => \receive_module.rx_counter.n3723\,
            clk => \N__19326\,
            ce => 'H',
            sr => \N__15952\
        );

    \receive_module.rx_counter.X_277__i5_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17050\,
            in2 => \_gnd_net_\,
            in3 => \N__15970\,
            lcout => \receive_module.rx_counter.X_4\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3723\,
            carryout => \receive_module.rx_counter.n3724\,
            clk => \N__19326\,
            ce => 'H',
            sr => \N__15952\
        );

    \receive_module.rx_counter.X_277__i6_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17073\,
            in2 => \_gnd_net_\,
            in3 => \N__15967\,
            lcout => \receive_module.rx_counter.X_5\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3724\,
            carryout => \receive_module.rx_counter.n3725\,
            clk => \N__19326\,
            ce => 'H',
            sr => \N__15952\
        );

    \receive_module.rx_counter.X_277__i7_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17412\,
            in2 => \_gnd_net_\,
            in3 => \N__15964\,
            lcout => \receive_module.rx_counter.X_6\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3725\,
            carryout => \receive_module.rx_counter.n3726\,
            clk => \N__19326\,
            ce => 'H',
            sr => \N__15952\
        );

    \receive_module.rx_counter.X_277__i8_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17442\,
            in2 => \_gnd_net_\,
            in3 => \N__15961\,
            lcout => \receive_module.rx_counter.X_7\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3726\,
            carryout => \receive_module.rx_counter.n3727\,
            clk => \N__19326\,
            ce => 'H',
            sr => \N__15952\
        );

    \receive_module.rx_counter.X_277__i9_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17502\,
            in2 => \_gnd_net_\,
            in3 => \N__15958\,
            lcout => \receive_module.rx_counter.X_8\,
            ltout => OPEN,
            carryin => \bfn_14_10_0_\,
            carryout => \receive_module.rx_counter.n3728\,
            clk => \N__19330\,
            ce => 'H',
            sr => \N__15948\
        );

    \receive_module.rx_counter.X_277__i10_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17475\,
            in2 => \_gnd_net_\,
            in3 => \N__15955\,
            lcout => \receive_module.rx_counter.X_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19330\,
            ce => 'H',
            sr => \N__15948\
        );

    \receive_module.rx_counter.i1_2_lut_4_lut_adj_27_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__15930\,
            in1 => \N__15891\,
            in2 => \N__15852\,
            in3 => \N__15761\,
            lcout => n658,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.X_DELTA_PATTERN_i9_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16066\,
            lcout => \transmit_module.X_DELTA_PATTERN_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22619\,
            ce => \N__17578\,
            sr => \N__20565\
        );

    \transmit_module.X_DELTA_PATTERN_i12_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16090\,
            lcout => \transmit_module.X_DELTA_PATTERN_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22619\,
            ce => \N__17578\,
            sr => \N__20565\
        );

    \transmit_module.X_DELTA_PATTERN_i13_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17629\,
            lcout => \transmit_module.X_DELTA_PATTERN_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22619\,
            ce => \N__17578\,
            sr => \N__20565\
        );

    \transmit_module.X_DELTA_PATTERN_i8_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16084\,
            lcout => \transmit_module.X_DELTA_PATTERN_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22619\,
            ce => \N__17578\,
            sr => \N__20565\
        );

    \transmit_module.X_DELTA_PATTERN_i11_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16078\,
            lcout => \transmit_module.X_DELTA_PATTERN_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22619\,
            ce => \N__17578\,
            sr => \N__20565\
        );

    \transmit_module.X_DELTA_PATTERN_i10_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16072\,
            lcout => \transmit_module.X_DELTA_PATTERN_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22619\,
            ce => \N__17578\,
            sr => \N__20565\
        );

    \line_buffer.TX_ADDR_12__bdd_4_lut_2663_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111110100000"
        )
    port map (
            in0 => \N__17281\,
            in1 => \N__16060\,
            in2 => \N__22858\,
            in3 => \N__23836\,
            lcout => \line_buffer.n4134\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i2_4_lut_LC_14_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011110000"
        )
    port map (
            in0 => \N__19583\,
            in1 => \N__19120\,
            in2 => \N__21194\,
            in3 => \N__19525\,
            lcout => \transmit_module.n2315\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.X_DELTA_PATTERN_i0_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17614\,
            lcout => \transmit_module.X_DELTA_PATTERN_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22560\,
            ce => \N__17583\,
            sr => \N__16025\
        );

    \transmit_module.ADDR_Y_COMPONENT__i4_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18991\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22498\,
            ce => \N__19876\,
            sr => \N__21317\
        );

    \transmit_module.ADDR_Y_COMPONENT__i2_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17824\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22498\,
            ce => \N__19876\,
            sr => \N__21317\
        );

    \transmit_module.BRAM_ADDR__i8_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011100100"
        )
    port map (
            in0 => \N__20195\,
            in1 => \N__16987\,
            in2 => \N__17008\,
            in3 => \N__21209\,
            lcout => \transmit_module.TX_ADDR_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22470\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i0_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__17838\,
            in1 => \N__16360\,
            in2 => \N__21292\,
            in3 => \N__20191\,
            lcout => \transmit_module.TX_ADDR_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22470\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i10_3_lut_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__19697\,
            in1 => \N__18433\,
            in2 => \_gnd_net_\,
            in3 => \N__18457\,
            lcout => \transmit_module.n179\,
            ltout => \transmit_module.n179_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i9_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001000100"
        )
    port map (
            in0 => \N__21198\,
            in1 => \N__16321\,
            in2 => \N__16348\,
            in3 => \N__20196\,
            lcout => \transmit_module.TX_ADDR_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22470\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i7_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__20194\,
            in1 => \N__21199\,
            in2 => \N__16663\,
            in3 => \N__16654\,
            lcout => \transmit_module.TX_ADDR_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22470\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i6_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__16413\,
            in1 => \N__16341\,
            in2 => \N__21294\,
            in3 => \N__20193\,
            lcout => \transmit_module.TX_ADDR_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22470\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i143_2_lut_3_lut_4_lut_rep_33_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101100"
        )
    port map (
            in0 => \N__16760\,
            in1 => \N__21197\,
            in2 => \N__19533\,
            in3 => \N__16719\,
            lcout => \transmit_module.n4224\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i3_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__20274\,
            in1 => \N__20259\,
            in2 => \N__21293\,
            in3 => \N__20192\,
            lcout => \transmit_module.TX_ADDR_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22470\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1772_4_lut_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__16327\,
            in1 => \N__16320\,
            in2 => \N__21180\,
            in3 => \N__20170\,
            lcout => n19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1771_4_lut_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__20169\,
            in1 => \N__21034\,
            in2 => \N__17004\,
            in3 => \N__16986\,
            lcout => n20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_2_lut_rep_29_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16755\,
            in2 => \_gnd_net_\,
            in3 => \N__16718\,
            lcout => \transmit_module.n4220\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i8_3_lut_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__19701\,
            in1 => \N__16429\,
            in2 => \_gnd_net_\,
            in3 => \N__17708\,
            lcout => \transmit_module.n181\,
            ltout => \transmit_module.n181_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1770_4_lut_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001000100"
        )
    port map (
            in0 => \N__21033\,
            in1 => \N__16653\,
            in2 => \N__16642\,
            in3 => \N__20168\,
            lcout => n21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.ADDR_Y_COMPONENT__i7_LC_14_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17713\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22347\,
            ce => \N__19869\,
            sr => \N__21307\
        );

    \transmit_module.ADDR_Y_COMPONENT__i1_LC_14_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18322\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22314\,
            ce => \N__19875\,
            sr => \N__21340\
        );

    \transmit_module.mux_12_i7_3_lut_LC_14_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__19713\,
            in1 => \N__16420\,
            in2 => \_gnd_net_\,
            in3 => \N__17757\,
            lcout => \transmit_module.n182\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.FRAME_COUNTER_278__i0_LC_15_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16393\,
            in2 => \_gnd_net_\,
            in3 => \N__16381\,
            lcout => \receive_module.rx_counter.FRAME_COUNTER_0\,
            ltout => OPEN,
            carryin => \bfn_15_8_0_\,
            carryout => \receive_module.rx_counter.n3706\,
            clk => \N__19322\,
            ce => \N__17332\,
            sr => \N__17128\
        );

    \receive_module.rx_counter.FRAME_COUNTER_278__i1_LC_15_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16378\,
            in2 => \_gnd_net_\,
            in3 => \N__17191\,
            lcout => \receive_module.rx_counter.FRAME_COUNTER_1\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3706\,
            carryout => \receive_module.rx_counter.n3707\,
            clk => \N__19322\,
            ce => \N__17332\,
            sr => \N__17128\
        );

    \receive_module.rx_counter.FRAME_COUNTER_278__i2_LC_15_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17188\,
            in2 => \_gnd_net_\,
            in3 => \N__17176\,
            lcout => \receive_module.rx_counter.FRAME_COUNTER_2\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3707\,
            carryout => \receive_module.rx_counter.n3708\,
            clk => \N__19322\,
            ce => \N__17332\,
            sr => \N__17128\
        );

    \receive_module.rx_counter.FRAME_COUNTER_278__i3_LC_15_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17173\,
            in2 => \_gnd_net_\,
            in3 => \N__17161\,
            lcout => \receive_module.rx_counter.FRAME_COUNTER_3\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3708\,
            carryout => \receive_module.rx_counter.n3709\,
            clk => \N__19322\,
            ce => \N__17332\,
            sr => \N__17128\
        );

    \receive_module.rx_counter.FRAME_COUNTER_278__i4_LC_15_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17158\,
            in2 => \_gnd_net_\,
            in3 => \N__17146\,
            lcout => \receive_module.rx_counter.FRAME_COUNTER_4\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3709\,
            carryout => \receive_module.rx_counter.n3710\,
            clk => \N__19322\,
            ce => \N__17332\,
            sr => \N__17128\
        );

    \receive_module.rx_counter.FRAME_COUNTER_278__i5_LC_15_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17140\,
            in2 => \_gnd_net_\,
            in3 => \N__17143\,
            lcout => \receive_module.rx_counter.FRAME_COUNTER_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19322\,
            ce => \N__17332\,
            sr => \N__17128\
        );

    \receive_module.rx_counter.old_VS_51_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17099\,
            lcout => \receive_module.rx_counter.old_VS\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19324\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1360_2_lut_3_lut_LC_15_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__17097\,
            in1 => \N__17118\,
            in2 => \_gnd_net_\,
            in3 => \N__17370\,
            lcout => \receive_module.rx_counter.n2605\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i150_2_lut_rep_31_LC_15_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__17119\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17098\,
            lcout => \receive_module.rx_counter.n4222\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i2_3_lut_rep_28_LC_15_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__17072\,
            in1 => \N__17049\,
            in2 => \_gnd_net_\,
            in3 => \N__17028\,
            lcout => \receive_module.rx_counter.n4219\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1_2_lut_adj_20_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17498\,
            in2 => \_gnd_net_\,
            in3 => \N__17471\,
            lcout => OPEN,
            ltout => \receive_module.rx_counter.n4_adj_575_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i2_4_lut_adj_21_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111000"
        )
    port map (
            in0 => \N__17449\,
            in1 => \N__17441\,
            in2 => \N__17419\,
            in3 => \N__17408\,
            lcout => \receive_module.rx_counter.O_VISIBLE_N_86\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.PULSE_1HZ_48_LC_15_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__17374\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17343\,
            lcout => \LED_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19327\,
            ce => \N__17331\,
            sr => \_gnd_net_\
        );

    \line_buffer.i2597_3_lut_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__23492\,
            in1 => \N__17320\,
            in2 => \_gnd_net_\,
            in3 => \N__17302\,
            lcout => \line_buffer.n4071\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_2698_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__17272\,
            in1 => \N__23846\,
            in2 => \N__17260\,
            in3 => \N__23493\,
            lcout => OPEN,
            ltout => \line_buffer.n4176_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n4176_bdd_4_lut_LC_15_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__23847\,
            in1 => \N__17239\,
            in2 => \N__17218\,
            in3 => \N__17215\,
            lcout => \line_buffer.n4179\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.X_DELTA_PATTERN_i7_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__17197\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.X_DELTA_PATTERN_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22514\,
            ce => \N__17582\,
            sr => \N__20587\
        );

    \transmit_module.X_DELTA_PATTERN_i5_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17635\,
            lcout => \transmit_module.X_DELTA_PATTERN_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22513\,
            ce => \N__17571\,
            sr => \N__20583\
        );

    \transmit_module.X_DELTA_PATTERN_i6_LC_15_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17641\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.X_DELTA_PATTERN_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22513\,
            ce => \N__17571\,
            sr => \N__20583\
        );

    \transmit_module.X_DELTA_PATTERN_i14_LC_15_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17602\,
            lcout => \transmit_module.X_DELTA_PATTERN_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22248\,
            ce => \N__17584\,
            sr => \N__20550\
        );

    \transmit_module.X_DELTA_PATTERN_i2_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17608\,
            lcout => \transmit_module.X_DELTA_PATTERN_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22248\,
            ce => \N__17584\,
            sr => \N__20550\
        );

    \transmit_module.X_DELTA_PATTERN_i1_LC_15_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17620\,
            lcout => \transmit_module.X_DELTA_PATTERN_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22248\,
            ce => \N__17584\,
            sr => \N__20550\
        );

    \transmit_module.X_DELTA_PATTERN_i3_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17590\,
            lcout => \transmit_module.X_DELTA_PATTERN_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22248\,
            ce => \N__17584\,
            sr => \N__20550\
        );

    \transmit_module.X_DELTA_PATTERN_i15_LC_15_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17535\,
            lcout => \transmit_module.X_DELTA_PATTERN_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22248\,
            ce => \N__17584\,
            sr => \N__20550\
        );

    \transmit_module.X_DELTA_PATTERN_i4_LC_15_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__17596\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.X_DELTA_PATTERN_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22248\,
            ce => \N__17584\,
            sr => \N__20550\
        );

    \transmit_module.add_13_2_lut_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18406\,
            in2 => \N__17536\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.n204\,
            ltout => OPEN,
            carryin => \bfn_15_17_0_\,
            carryout => \transmit_module.n3656\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_3_lut_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18320\,
            in2 => \_gnd_net_\,
            in3 => \N__17506\,
            lcout => \transmit_module.n203\,
            ltout => OPEN,
            carryin => \transmit_module.n3656\,
            carryout => \transmit_module.n3657\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_4_lut_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17823\,
            in2 => \_gnd_net_\,
            in3 => \N__17785\,
            lcout => \transmit_module.n202\,
            ltout => OPEN,
            carryin => \transmit_module.n3657\,
            carryout => \transmit_module.n3658\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_5_lut_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18373\,
            in2 => \_gnd_net_\,
            in3 => \N__17767\,
            lcout => \transmit_module.n201\,
            ltout => OPEN,
            carryin => \transmit_module.n3658\,
            carryout => \transmit_module.n3659\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_6_lut_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18987\,
            in3 => \N__17764\,
            lcout => \transmit_module.n200\,
            ltout => OPEN,
            carryin => \transmit_module.n3659\,
            carryout => \transmit_module.n3660\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_7_lut_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19021\,
            in2 => \_gnd_net_\,
            in3 => \N__17761\,
            lcout => \transmit_module.n199\,
            ltout => OPEN,
            carryin => \transmit_module.n3660\,
            carryout => \transmit_module.n3661\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_8_lut_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17741\,
            in2 => \_gnd_net_\,
            in3 => \N__17716\,
            lcout => \transmit_module.n198\,
            ltout => OPEN,
            carryin => \transmit_module.n3661\,
            carryout => \transmit_module.n3662\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_9_lut_LC_15_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17704\,
            in2 => \_gnd_net_\,
            in3 => \N__17671\,
            lcout => \transmit_module.n197\,
            ltout => OPEN,
            carryin => \transmit_module.n3662\,
            carryout => \transmit_module.n3663\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_10_lut_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17884\,
            in2 => \_gnd_net_\,
            in3 => \N__17656\,
            lcout => \transmit_module.n196\,
            ltout => OPEN,
            carryin => \bfn_15_18_0_\,
            carryout => \transmit_module.n3664\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_11_lut_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18464\,
            in3 => \N__17644\,
            lcout => \transmit_module.n195\,
            ltout => OPEN,
            carryin => \transmit_module.n3664\,
            carryout => \transmit_module.n3665\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_12_lut_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17956\,
            in2 => \_gnd_net_\,
            in3 => \N__17905\,
            lcout => \transmit_module.n194\,
            ltout => OPEN,
            carryin => \transmit_module.n3665\,
            carryout => \transmit_module.n3666\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_13_lut_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23518\,
            in2 => \_gnd_net_\,
            in3 => \N__17902\,
            lcout => \transmit_module.n193\,
            ltout => OPEN,
            carryin => \transmit_module.n3666\,
            carryout => \transmit_module.n3667\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_14_lut_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23806\,
            in3 => \N__17899\,
            lcout => \transmit_module.n192\,
            ltout => OPEN,
            carryin => \transmit_module.n3667\,
            carryout => \transmit_module.n3668\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_15_lut_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__22802\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17896\,
            lcout => \transmit_module.n191\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.ADDR_Y_COMPONENT__i8_LC_15_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__17885\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22445\,
            ce => \N__19853\,
            sr => \N__21210\
        );

    \transmit_module.mux_12_i4_3_lut_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__18352\,
            in1 => \N__19670\,
            in2 => \_gnd_net_\,
            in3 => \N__18374\,
            lcout => \transmit_module.n185\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.mux_14_i2_3_lut_4_lut_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__18319\,
            in1 => \N__19128\,
            in2 => \N__17854\,
            in3 => \N__19521\,
            lcout => \transmit_module.n218\,
            ltout => \transmit_module.n218_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i1_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001010000"
        )
    port map (
            in0 => \N__21179\,
            in1 => \N__18292\,
            in2 => \N__17842\,
            in3 => \N__20209\,
            lcout => \transmit_module.TX_ADDR_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22352\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i1_3_lut_LC_15_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__19691\,
            in1 => \N__18385\,
            in2 => \_gnd_net_\,
            in3 => \N__18407\,
            lcout => \transmit_module.n188\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.ADDR_Y_COMPONENT__i0_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18421\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22070\,
            ce => \N__19874\,
            sr => \N__21181\
        );

    \transmit_module.ADDR_Y_COMPONENT__i11_LC_15_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23485\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22070\,
            ce => \N__19874\,
            sr => \N__21181\
        );

    \transmit_module.ADDR_Y_COMPONENT__i3_LC_15_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18379\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22070\,
            ce => \N__19874\,
            sr => \N__21181\
        );

    \transmit_module.BRAM_ADDR__rep_1_i0_LC_15_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__19582\,
            in1 => \N__18346\,
            in2 => \N__18337\,
            in3 => \N__19532\,
            lcout => \TX_ADDR_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22062\,
            ce => \N__19410\,
            sr => \N__21338\
        );

    \transmit_module.mux_12_i2_3_lut_LC_15_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__19693\,
            in1 => \N__18328\,
            in2 => \_gnd_net_\,
            in3 => \N__18321\,
            lcout => \transmit_module.n187\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1764_4_lut_LC_15_27_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__18291\,
            in1 => \N__18274\,
            in2 => \N__21336\,
            in3 => \N__20240\,
            lcout => n27,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_LC_16_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__18049\,
            in1 => \N__23848\,
            in2 => \N__18031\,
            in3 => \N__23611\,
            lcout => OPEN,
            ltout => \line_buffer.n4188_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n4188_bdd_4_lut_LC_16_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__23849\,
            in1 => \N__18019\,
            in2 => \N__18001\,
            in3 => \N__17998\,
            lcout => OPEN,
            ltout => \line_buffer.n4191_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i5_LC_16_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22856\,
            in2 => \N__17980\,
            in3 => \N__17977\,
            lcout => \TX_DATA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22421\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.Y_DELTA_PATTERN_i18_LC_16_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18481\,
            lcout => \transmit_module.Y_DELTA_PATTERN_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22247\,
            ce => \N__20597\,
            sr => \N__21147\
        );

    \transmit_module.Y_DELTA_PATTERN_i20_LC_16_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18493\,
            lcout => \transmit_module.Y_DELTA_PATTERN_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22247\,
            ce => \N__20597\,
            sr => \N__21147\
        );

    \transmit_module.Y_DELTA_PATTERN_i0_LC_16_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18475\,
            lcout => \transmit_module.Y_DELTA_PATTERN_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22247\,
            ce => \N__20597\,
            sr => \N__21147\
        );

    \transmit_module.Y_DELTA_PATTERN_i17_LC_16_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18499\,
            lcout => \transmit_module.Y_DELTA_PATTERN_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22247\,
            ce => \N__20597\,
            sr => \N__21147\
        );

    \transmit_module.Y_DELTA_PATTERN_i21_LC_16_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20647\,
            lcout => \transmit_module.Y_DELTA_PATTERN_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22247\,
            ce => \N__20597\,
            sr => \N__21147\
        );

    \transmit_module.Y_DELTA_PATTERN_i19_LC_16_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18487\,
            lcout => \transmit_module.Y_DELTA_PATTERN_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22247\,
            ce => \N__20597\,
            sr => \N__21147\
        );

    \transmit_module.Y_DELTA_PATTERN_i1_LC_16_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20656\,
            lcout => \transmit_module.Y_DELTA_PATTERN_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22247\,
            ce => \N__20597\,
            sr => \N__21147\
        );

    \transmit_module.ADDR_Y_COMPONENT__i5_LC_16_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19026\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22243\,
            ce => \N__19877\,
            sr => \N__21341\
        );

    \transmit_module.ADDR_Y_COMPONENT__i9_LC_16_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18469\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22243\,
            ce => \N__19877\,
            sr => \N__21341\
        );

    \transmit_module.video_signal_controller.mux_14_i5_3_lut_4_lut_LC_16_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__18983\,
            in1 => \N__19126\,
            in2 => \N__19174\,
            in3 => \N__19512\,
            lcout => \transmit_module.n215\,
            ltout => \transmit_module.n215_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i4_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001010000"
        )
    port map (
            in0 => \N__21217\,
            in1 => \N__18961\,
            in2 => \N__19165\,
            in3 => \N__20228\,
            lcout => \transmit_module.TX_ADDR_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22444\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i6_3_lut_LC_16_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__19663\,
            in1 => \N__19162\,
            in2 => \_gnd_net_\,
            in3 => \N__19022\,
            lcout => \transmit_module.n183\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.mux_18_i14_3_lut_4_lut_LC_16_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__19513\,
            in1 => \N__19587\,
            in2 => \N__19897\,
            in3 => \N__19156\,
            lcout => \transmit_module.BRAM_ADDR_13_N_258_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.mux_14_i6_3_lut_4_lut_LC_16_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__19511\,
            in1 => \N__19138\,
            in2 => \N__19027\,
            in3 => \N__19127\,
            lcout => \transmit_module.n214\,
            ltout => \transmit_module.n214_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i5_LC_16_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__20229\,
            in1 => \N__21218\,
            in2 => \N__19030\,
            in3 => \N__18732\,
            lcout => \transmit_module.TX_ADDR_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22444\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i5_3_lut_LC_16_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__19662\,
            in1 => \N__19003\,
            in2 => \_gnd_net_\,
            in3 => \N__18982\,
            lcout => \transmit_module.n184\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1767_4_lut_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__18960\,
            in1 => \N__18949\,
            in2 => \N__21280\,
            in3 => \N__20197\,
            lcout => n24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1768_4_lut_LC_16_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__20198\,
            in1 => \N__21172\,
            in2 => \N__18733\,
            in3 => \N__18718\,
            lcout => n23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i12_LC_16_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__19588\,
            in1 => \N__19543\,
            in2 => \N__19906\,
            in3 => \N__19534\,
            lcout => \TX_ADDR_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22069\,
            ce => \N__19411\,
            sr => \N__21260\
        );

    \transmit_module.Y_DELTA_PATTERN_i41_LC_16_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19381\,
            lcout => \transmit_module.Y_DELTA_PATTERN_41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22061\,
            ce => \N__21459\,
            sr => \N__21339\
        );

    \GB_BUFFER_DEBUG_c_1_c_THRU_LUT4_0_LC_16_30_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19372\,
            lcout => \GB_BUFFER_DEBUG_c_1_c_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.Y_DELTA_PATTERN_i5_LC_17_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20350\,
            lcout => \transmit_module.Y_DELTA_PATTERN_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22565\,
            ce => \N__20622\,
            sr => \N__21295\
        );

    \transmit_module.Y_DELTA_PATTERN_i28_LC_17_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19192\,
            lcout => \transmit_module.Y_DELTA_PATTERN_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22420\,
            ce => \N__20599\,
            sr => \N__21266\
        );

    \transmit_module.Y_DELTA_PATTERN_i31_LC_17_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19762\,
            lcout => \transmit_module.Y_DELTA_PATTERN_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22420\,
            ce => \N__20599\,
            sr => \N__21266\
        );

    \transmit_module.Y_DELTA_PATTERN_i29_LC_17_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19180\,
            lcout => \transmit_module.Y_DELTA_PATTERN_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22420\,
            ce => \N__20599\,
            sr => \N__21266\
        );

    \transmit_module.Y_DELTA_PATTERN_i30_LC_17_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19186\,
            lcout => \transmit_module.Y_DELTA_PATTERN_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22420\,
            ce => \N__20599\,
            sr => \N__21266\
        );

    \transmit_module.Y_DELTA_PATTERN_i12_LC_17_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19756\,
            lcout => \transmit_module.Y_DELTA_PATTERN_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22548\,
            ce => \N__20614\,
            sr => \N__21324\
        );

    \transmit_module.Y_DELTA_PATTERN_i11_LC_17_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19768\,
            lcout => \transmit_module.Y_DELTA_PATTERN_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22548\,
            ce => \N__20614\,
            sr => \N__21324\
        );

    \transmit_module.Y_DELTA_PATTERN_i32_LC_17_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21523\,
            lcout => \transmit_module.Y_DELTA_PATTERN_32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22548\,
            ce => \N__20614\,
            sr => \N__21324\
        );

    \transmit_module.Y_DELTA_PATTERN_i13_LC_17_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19750\,
            lcout => \transmit_module.Y_DELTA_PATTERN_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22548\,
            ce => \N__20614\,
            sr => \N__21324\
        );

    \transmit_module.Y_DELTA_PATTERN_i14_LC_17_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20308\,
            lcout => \transmit_module.Y_DELTA_PATTERN_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22548\,
            ce => \N__20614\,
            sr => \N__21324\
        );

    \transmit_module.Y_DELTA_PATTERN_i26_LC_17_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19723\,
            lcout => \transmit_module.Y_DELTA_PATTERN_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22573\,
            ce => \N__20598\,
            sr => \N__21343\
        );

    \transmit_module.Y_DELTA_PATTERN_i24_LC_17_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19738\,
            lcout => \transmit_module.Y_DELTA_PATTERN_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22573\,
            ce => \N__20598\,
            sr => \N__21343\
        );

    \transmit_module.Y_DELTA_PATTERN_i25_LC_17_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19744\,
            lcout => \transmit_module.Y_DELTA_PATTERN_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22573\,
            ce => \N__20598\,
            sr => \N__21343\
        );

    \transmit_module.Y_DELTA_PATTERN_i27_LC_17_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19732\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.Y_DELTA_PATTERN_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22573\,
            ce => \N__20598\,
            sr => \N__21343\
        );

    \transmit_module.Y_DELTA_PATTERN_i99_LC_17_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19661\,
            lcout => \transmit_module.Y_DELTA_PATTERN_99\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22573\,
            ce => \N__20598\,
            sr => \N__21343\
        );

    \transmit_module.Y_DELTA_PATTERN_i37_LC_17_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20281\,
            lcout => \transmit_module.Y_DELTA_PATTERN_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22466\,
            ce => \N__21473\,
            sr => \N__21262\
        );

    \transmit_module.Y_DELTA_PATTERN_i35_LC_17_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20287\,
            lcout => \transmit_module.Y_DELTA_PATTERN_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22466\,
            ce => \N__21473\,
            sr => \N__21262\
        );

    \transmit_module.Y_DELTA_PATTERN_i36_LC_17_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20293\,
            lcout => \transmit_module.Y_DELTA_PATTERN_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22466\,
            ce => \N__21473\,
            sr => \N__21262\
        );

    \transmit_module.Y_DELTA_PATTERN_i38_LC_17_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__19789\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.Y_DELTA_PATTERN_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22466\,
            ce => \N__21473\,
            sr => \N__21262\
        );

    \transmit_module.i1766_4_lut_LC_17_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__20275\,
            in1 => \N__20260\,
            in2 => \N__21281\,
            in3 => \N__20216\,
            lcout => n25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.ADDR_Y_COMPONENT__i12_LC_17_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23741\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22440\,
            ce => \N__19870\,
            sr => \N__21261\
        );

    \transmit_module.ADDR_Y_COMPONENT__i13_LC_17_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22818\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22440\,
            ce => \N__19870\,
            sr => \N__21261\
        );

    \transmit_module.Y_DELTA_PATTERN_i39_LC_17_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19774\,
            lcout => \transmit_module.Y_DELTA_PATTERN_39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22340\,
            ce => \N__21487\,
            sr => \N__21337\
        );

    \transmit_module.Y_DELTA_PATTERN_i40_LC_17_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19780\,
            lcout => \transmit_module.Y_DELTA_PATTERN_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22340\,
            ce => \N__21487\,
            sr => \N__21337\
        );

    \line_buffer.i2591_3_lut_LC_18_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__20377\,
            in1 => \N__20359\,
            in2 => \_gnd_net_\,
            in3 => \N__23535\,
            lcout => \line_buffer.n4065\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.Y_DELTA_PATTERN_i6_LC_18_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20338\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.Y_DELTA_PATTERN_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22572\,
            ce => \N__20623\,
            sr => \N__21296\
        );

    \transmit_module.Y_DELTA_PATTERN_i4_LC_18_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20344\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.Y_DELTA_PATTERN_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22572\,
            ce => \N__20623\,
            sr => \N__21296\
        );

    \transmit_module.Y_DELTA_PATTERN_i9_LC_18_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20326\,
            lcout => \transmit_module.Y_DELTA_PATTERN_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22419\,
            ce => \N__20618\,
            sr => \N__21323\
        );

    \transmit_module.Y_DELTA_PATTERN_i7_LC_18_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20314\,
            lcout => \transmit_module.Y_DELTA_PATTERN_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22419\,
            ce => \N__20618\,
            sr => \N__21323\
        );

    \transmit_module.Y_DELTA_PATTERN_i10_LC_18_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__20332\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.Y_DELTA_PATTERN_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22419\,
            ce => \N__20618\,
            sr => \N__21323\
        );

    \transmit_module.Y_DELTA_PATTERN_i8_LC_18_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20320\,
            lcout => \transmit_module.Y_DELTA_PATTERN_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22419\,
            ce => \N__20618\,
            sr => \N__21323\
        );

    \transmit_module.Y_DELTA_PATTERN_i15_LC_18_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20668\,
            lcout => \transmit_module.Y_DELTA_PATTERN_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22562\,
            ce => \N__20607\,
            sr => \N__21267\
        );

    \transmit_module.Y_DELTA_PATTERN_i3_LC_18_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20302\,
            lcout => \transmit_module.Y_DELTA_PATTERN_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22562\,
            ce => \N__20607\,
            sr => \N__21267\
        );

    \transmit_module.Y_DELTA_PATTERN_i16_LC_18_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20677\,
            lcout => \transmit_module.Y_DELTA_PATTERN_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22562\,
            ce => \N__20607\,
            sr => \N__21267\
        );

    \transmit_module.Y_DELTA_PATTERN_i2_LC_18_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20662\,
            lcout => \transmit_module.Y_DELTA_PATTERN_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22562\,
            ce => \N__20607\,
            sr => \N__21267\
        );

    \transmit_module.Y_DELTA_PATTERN_i22_LC_18_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20629\,
            lcout => \transmit_module.Y_DELTA_PATTERN_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22512\,
            ce => \N__20606\,
            sr => \N__21342\
        );

    \transmit_module.Y_DELTA_PATTERN_i23_LC_18_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20635\,
            lcout => \transmit_module.Y_DELTA_PATTERN_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22512\,
            ce => \N__20606\,
            sr => \N__21342\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_2688_LC_18_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__23602\,
            in1 => \N__20485\,
            in2 => \N__20470\,
            in3 => \N__23842\,
            lcout => OPEN,
            ltout => \line_buffer.n4164_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n4164_bdd_4_lut_LC_18_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__23843\,
            in1 => \N__20449\,
            in2 => \N__20428\,
            in3 => \N__20425\,
            lcout => OPEN,
            ltout => \line_buffer.n4167_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i1_LC_18_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22835\,
            in2 => \N__20407\,
            in3 => \N__20683\,
            lcout => \TX_DATA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22474\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_12__bdd_4_lut_2658_LC_18_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111110100000"
        )
    port map (
            in0 => \N__20389\,
            in1 => \N__21628\,
            in2 => \N__22857\,
            in3 => \N__23829\,
            lcout => \line_buffer.n4128\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2592_3_lut_LC_18_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21664\,
            in1 => \N__21646\,
            in2 => \_gnd_net_\,
            in3 => \N__23598\,
            lcout => \line_buffer.n4066\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2600_3_lut_LC_18_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__23600\,
            in1 => \N__21622\,
            in2 => \_gnd_net_\,
            in3 => \N__21607\,
            lcout => OPEN,
            ltout => \line_buffer.n4074_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i3_LC_18_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__22819\,
            in1 => \N__21529\,
            in2 => \N__21589\,
            in3 => \N__21586\,
            lcout => \TX_DATA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22465\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2601_3_lut_LC_18_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__23599\,
            in1 => \N__21571\,
            in2 => \_gnd_net_\,
            in3 => \N__21547\,
            lcout => \line_buffer.n4075\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.Y_DELTA_PATTERN_i33_LC_19_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21499\,
            lcout => \transmit_module.Y_DELTA_PATTERN_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22574\,
            ce => \N__21488\,
            sr => \N__21322\
        );

    \transmit_module.Y_DELTA_PATTERN_i34_LC_19_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21511\,
            lcout => \transmit_module.Y_DELTA_PATTERN_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22574\,
            ce => \N__21488\,
            sr => \N__21322\
        );

    \line_buffer.n4146_bdd_4_lut_LC_19_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__20761\,
            in1 => \N__22972\,
            in2 => \N__20746\,
            in3 => \N__23841\,
            lcout => \line_buffer.n4149\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n4158_bdd_4_lut_LC_19_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001000100"
        )
    port map (
            in0 => \N__23840\,
            in1 => \N__20725\,
            in2 => \N__20707\,
            in3 => \N__23659\,
            lcout => \line_buffer.n4161\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_2673_LC_19_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__23011\,
            in1 => \N__23828\,
            in2 => \N__22990\,
            in3 => \N__23601\,
            lcout => \line_buffer.n4146\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i0_LC_19_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__22842\,
            in1 => \N__21670\,
            in2 => \_gnd_net_\,
            in3 => \N__22966\,
            lcout => \TX_DATA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22487\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2588_3_lut_LC_20_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22945\,
            in1 => \N__22933\,
            in2 => \_gnd_net_\,
            in3 => \N__23536\,
            lcout => \line_buffer.n4062\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2604_3_lut_LC_20_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22918\,
            in1 => \N__22906\,
            in2 => \_gnd_net_\,
            in3 => \N__23614\,
            lcout => \line_buffer.n4078\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_12__bdd_4_lut_LC_20_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111111000000"
        )
    port map (
            in0 => \N__23401\,
            in1 => \N__22891\,
            in2 => \N__22869\,
            in3 => \N__23859\,
            lcout => \line_buffer.n4140\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i4_LC_20_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__22882\,
            in1 => \N__22865\,
            in2 => \N__23893\,
            in3 => \N__22714\,
            lcout => \TX_DATA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22621\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_2649_LC_20_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__21739\,
            in1 => \N__23850\,
            in2 => \N__21724\,
            in3 => \N__23577\,
            lcout => \line_buffer.n4116\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n4116_bdd_4_lut_LC_20_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__21709\,
            in1 => \N__21694\,
            in2 => \N__21688\,
            in3 => \N__23851\,
            lcout => \line_buffer.n4119\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2603_3_lut_LC_20_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__23590\,
            in1 => \N__23923\,
            in2 => \_gnd_net_\,
            in3 => \N__23908\,
            lcout => \line_buffer.n4077\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_2683_LC_20_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__23881\,
            in1 => \N__23818\,
            in2 => \N__23674\,
            in3 => \N__23586\,
            lcout => \line_buffer.n4158\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2589_3_lut_LC_21_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__23653\,
            in1 => \N__23635\,
            in2 => \_gnd_net_\,
            in3 => \N__23612\,
            lcout => \line_buffer.n4063\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_24_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
