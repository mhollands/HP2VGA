-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     Oct 7 2018 19:46:25

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "main" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of main
entity main is
port (
    TVP_VIDEO : in std_logic_vector(9 downto 0);
    ADV_B : out std_logic_vector(7 downto 0);
    ADV_G : out std_logic_vector(7 downto 0);
    ADV_R : out std_logic_vector(7 downto 0);
    DEBUG : inout std_logic_vector(7 downto 0);
    TVP_CLK : in std_logic;
    ADV_CLK : out std_logic;
    TVP_HSYNC : in std_logic;
    ADV_HSYNC : out std_logic;
    TVP_VSYNC : in std_logic;
    ADV_VSYNC : out std_logic;
    ADV_BLANK_N : out std_logic;
    LED : out std_logic;
    ADV_SYNC_N : out std_logic);
end main;

-- Architecture of main
-- View name is \INTERFACE\
architecture \INTERFACE\ of main is

signal \N__25265\ : std_logic;
signal \N__25264\ : std_logic;
signal \N__25263\ : std_logic;
signal \N__25254\ : std_logic;
signal \N__25253\ : std_logic;
signal \N__25252\ : std_logic;
signal \N__25245\ : std_logic;
signal \N__25244\ : std_logic;
signal \N__25243\ : std_logic;
signal \N__25236\ : std_logic;
signal \N__25235\ : std_logic;
signal \N__25234\ : std_logic;
signal \N__25227\ : std_logic;
signal \N__25226\ : std_logic;
signal \N__25225\ : std_logic;
signal \N__25218\ : std_logic;
signal \N__25217\ : std_logic;
signal \N__25216\ : std_logic;
signal \N__25209\ : std_logic;
signal \N__25208\ : std_logic;
signal \N__25207\ : std_logic;
signal \N__25200\ : std_logic;
signal \N__25199\ : std_logic;
signal \N__25198\ : std_logic;
signal \N__25191\ : std_logic;
signal \N__25190\ : std_logic;
signal \N__25189\ : std_logic;
signal \N__25182\ : std_logic;
signal \N__25181\ : std_logic;
signal \N__25180\ : std_logic;
signal \N__25173\ : std_logic;
signal \N__25172\ : std_logic;
signal \N__25171\ : std_logic;
signal \N__25164\ : std_logic;
signal \N__25163\ : std_logic;
signal \N__25162\ : std_logic;
signal \N__25155\ : std_logic;
signal \N__25154\ : std_logic;
signal \N__25153\ : std_logic;
signal \N__25146\ : std_logic;
signal \N__25145\ : std_logic;
signal \N__25144\ : std_logic;
signal \N__25137\ : std_logic;
signal \N__25136\ : std_logic;
signal \N__25135\ : std_logic;
signal \N__25128\ : std_logic;
signal \N__25127\ : std_logic;
signal \N__25126\ : std_logic;
signal \N__25119\ : std_logic;
signal \N__25118\ : std_logic;
signal \N__25117\ : std_logic;
signal \N__25110\ : std_logic;
signal \N__25109\ : std_logic;
signal \N__25108\ : std_logic;
signal \N__25101\ : std_logic;
signal \N__25100\ : std_logic;
signal \N__25099\ : std_logic;
signal \N__25092\ : std_logic;
signal \N__25091\ : std_logic;
signal \N__25090\ : std_logic;
signal \N__25083\ : std_logic;
signal \N__25082\ : std_logic;
signal \N__25081\ : std_logic;
signal \N__25074\ : std_logic;
signal \N__25073\ : std_logic;
signal \N__25072\ : std_logic;
signal \N__25065\ : std_logic;
signal \N__25064\ : std_logic;
signal \N__25063\ : std_logic;
signal \N__25056\ : std_logic;
signal \N__25055\ : std_logic;
signal \N__25054\ : std_logic;
signal \N__25047\ : std_logic;
signal \N__25046\ : std_logic;
signal \N__25045\ : std_logic;
signal \N__25038\ : std_logic;
signal \N__25037\ : std_logic;
signal \N__25036\ : std_logic;
signal \N__25029\ : std_logic;
signal \N__25028\ : std_logic;
signal \N__25027\ : std_logic;
signal \N__25020\ : std_logic;
signal \N__25019\ : std_logic;
signal \N__25018\ : std_logic;
signal \N__25011\ : std_logic;
signal \N__25010\ : std_logic;
signal \N__25009\ : std_logic;
signal \N__25002\ : std_logic;
signal \N__25001\ : std_logic;
signal \N__25000\ : std_logic;
signal \N__24993\ : std_logic;
signal \N__24992\ : std_logic;
signal \N__24991\ : std_logic;
signal \N__24984\ : std_logic;
signal \N__24983\ : std_logic;
signal \N__24982\ : std_logic;
signal \N__24975\ : std_logic;
signal \N__24974\ : std_logic;
signal \N__24973\ : std_logic;
signal \N__24966\ : std_logic;
signal \N__24965\ : std_logic;
signal \N__24964\ : std_logic;
signal \N__24957\ : std_logic;
signal \N__24956\ : std_logic;
signal \N__24955\ : std_logic;
signal \N__24948\ : std_logic;
signal \N__24947\ : std_logic;
signal \N__24946\ : std_logic;
signal \N__24939\ : std_logic;
signal \N__24938\ : std_logic;
signal \N__24937\ : std_logic;
signal \N__24930\ : std_logic;
signal \N__24929\ : std_logic;
signal \N__24928\ : std_logic;
signal \N__24921\ : std_logic;
signal \N__24920\ : std_logic;
signal \N__24919\ : std_logic;
signal \N__24912\ : std_logic;
signal \N__24911\ : std_logic;
signal \N__24910\ : std_logic;
signal \N__24903\ : std_logic;
signal \N__24902\ : std_logic;
signal \N__24901\ : std_logic;
signal \N__24894\ : std_logic;
signal \N__24893\ : std_logic;
signal \N__24892\ : std_logic;
signal \N__24885\ : std_logic;
signal \N__24884\ : std_logic;
signal \N__24883\ : std_logic;
signal \N__24876\ : std_logic;
signal \N__24875\ : std_logic;
signal \N__24874\ : std_logic;
signal \N__24867\ : std_logic;
signal \N__24866\ : std_logic;
signal \N__24865\ : std_logic;
signal \N__24858\ : std_logic;
signal \N__24857\ : std_logic;
signal \N__24856\ : std_logic;
signal \N__24849\ : std_logic;
signal \N__24848\ : std_logic;
signal \N__24847\ : std_logic;
signal \N__24840\ : std_logic;
signal \N__24839\ : std_logic;
signal \N__24838\ : std_logic;
signal \N__24831\ : std_logic;
signal \N__24830\ : std_logic;
signal \N__24829\ : std_logic;
signal \N__24812\ : std_logic;
signal \N__24809\ : std_logic;
signal \N__24806\ : std_logic;
signal \N__24803\ : std_logic;
signal \N__24800\ : std_logic;
signal \N__24799\ : std_logic;
signal \N__24798\ : std_logic;
signal \N__24797\ : std_logic;
signal \N__24796\ : std_logic;
signal \N__24795\ : std_logic;
signal \N__24794\ : std_logic;
signal \N__24793\ : std_logic;
signal \N__24790\ : std_logic;
signal \N__24787\ : std_logic;
signal \N__24786\ : std_logic;
signal \N__24785\ : std_logic;
signal \N__24784\ : std_logic;
signal \N__24781\ : std_logic;
signal \N__24780\ : std_logic;
signal \N__24779\ : std_logic;
signal \N__24776\ : std_logic;
signal \N__24773\ : std_logic;
signal \N__24772\ : std_logic;
signal \N__24769\ : std_logic;
signal \N__24766\ : std_logic;
signal \N__24765\ : std_logic;
signal \N__24764\ : std_logic;
signal \N__24763\ : std_logic;
signal \N__24760\ : std_logic;
signal \N__24757\ : std_logic;
signal \N__24754\ : std_logic;
signal \N__24749\ : std_logic;
signal \N__24746\ : std_logic;
signal \N__24745\ : std_logic;
signal \N__24744\ : std_logic;
signal \N__24743\ : std_logic;
signal \N__24740\ : std_logic;
signal \N__24737\ : std_logic;
signal \N__24734\ : std_logic;
signal \N__24733\ : std_logic;
signal \N__24732\ : std_logic;
signal \N__24727\ : std_logic;
signal \N__24724\ : std_logic;
signal \N__24719\ : std_logic;
signal \N__24716\ : std_logic;
signal \N__24715\ : std_logic;
signal \N__24714\ : std_logic;
signal \N__24711\ : std_logic;
signal \N__24708\ : std_logic;
signal \N__24705\ : std_logic;
signal \N__24696\ : std_logic;
signal \N__24693\ : std_logic;
signal \N__24690\ : std_logic;
signal \N__24687\ : std_logic;
signal \N__24686\ : std_logic;
signal \N__24681\ : std_logic;
signal \N__24678\ : std_logic;
signal \N__24675\ : std_logic;
signal \N__24672\ : std_logic;
signal \N__24669\ : std_logic;
signal \N__24666\ : std_logic;
signal \N__24663\ : std_logic;
signal \N__24660\ : std_logic;
signal \N__24657\ : std_logic;
signal \N__24654\ : std_logic;
signal \N__24651\ : std_logic;
signal \N__24642\ : std_logic;
signal \N__24641\ : std_logic;
signal \N__24636\ : std_logic;
signal \N__24633\ : std_logic;
signal \N__24630\ : std_logic;
signal \N__24625\ : std_logic;
signal \N__24618\ : std_logic;
signal \N__24613\ : std_logic;
signal \N__24606\ : std_logic;
signal \N__24603\ : std_logic;
signal \N__24600\ : std_logic;
signal \N__24597\ : std_logic;
signal \N__24594\ : std_logic;
signal \N__24585\ : std_logic;
signal \N__24582\ : std_logic;
signal \N__24579\ : std_logic;
signal \N__24566\ : std_logic;
signal \N__24563\ : std_logic;
signal \N__24560\ : std_logic;
signal \N__24557\ : std_logic;
signal \N__24554\ : std_logic;
signal \N__24551\ : std_logic;
signal \N__24548\ : std_logic;
signal \N__24545\ : std_logic;
signal \N__24542\ : std_logic;
signal \N__24539\ : std_logic;
signal \N__24536\ : std_logic;
signal \N__24533\ : std_logic;
signal \N__24530\ : std_logic;
signal \N__24527\ : std_logic;
signal \N__24524\ : std_logic;
signal \N__24523\ : std_logic;
signal \N__24522\ : std_logic;
signal \N__24521\ : std_logic;
signal \N__24518\ : std_logic;
signal \N__24515\ : std_logic;
signal \N__24514\ : std_logic;
signal \N__24513\ : std_logic;
signal \N__24512\ : std_logic;
signal \N__24509\ : std_logic;
signal \N__24506\ : std_logic;
signal \N__24505\ : std_logic;
signal \N__24500\ : std_logic;
signal \N__24497\ : std_logic;
signal \N__24496\ : std_logic;
signal \N__24493\ : std_logic;
signal \N__24490\ : std_logic;
signal \N__24489\ : std_logic;
signal \N__24488\ : std_logic;
signal \N__24485\ : std_logic;
signal \N__24482\ : std_logic;
signal \N__24479\ : std_logic;
signal \N__24474\ : std_logic;
signal \N__24471\ : std_logic;
signal \N__24470\ : std_logic;
signal \N__24469\ : std_logic;
signal \N__24468\ : std_logic;
signal \N__24463\ : std_logic;
signal \N__24462\ : std_logic;
signal \N__24459\ : std_logic;
signal \N__24456\ : std_logic;
signal \N__24455\ : std_logic;
signal \N__24454\ : std_logic;
signal \N__24447\ : std_logic;
signal \N__24442\ : std_logic;
signal \N__24439\ : std_logic;
signal \N__24436\ : std_logic;
signal \N__24435\ : std_logic;
signal \N__24432\ : std_logic;
signal \N__24429\ : std_logic;
signal \N__24426\ : std_logic;
signal \N__24425\ : std_logic;
signal \N__24424\ : std_logic;
signal \N__24419\ : std_logic;
signal \N__24416\ : std_logic;
signal \N__24413\ : std_logic;
signal \N__24412\ : std_logic;
signal \N__24411\ : std_logic;
signal \N__24410\ : std_logic;
signal \N__24409\ : std_logic;
signal \N__24408\ : std_logic;
signal \N__24407\ : std_logic;
signal \N__24404\ : std_logic;
signal \N__24397\ : std_logic;
signal \N__24394\ : std_logic;
signal \N__24391\ : std_logic;
signal \N__24388\ : std_logic;
signal \N__24385\ : std_logic;
signal \N__24382\ : std_logic;
signal \N__24379\ : std_logic;
signal \N__24378\ : std_logic;
signal \N__24377\ : std_logic;
signal \N__24370\ : std_logic;
signal \N__24367\ : std_logic;
signal \N__24364\ : std_logic;
signal \N__24363\ : std_logic;
signal \N__24360\ : std_logic;
signal \N__24357\ : std_logic;
signal \N__24354\ : std_logic;
signal \N__24351\ : std_logic;
signal \N__24344\ : std_logic;
signal \N__24343\ : std_logic;
signal \N__24342\ : std_logic;
signal \N__24339\ : std_logic;
signal \N__24330\ : std_logic;
signal \N__24327\ : std_logic;
signal \N__24324\ : std_logic;
signal \N__24323\ : std_logic;
signal \N__24322\ : std_logic;
signal \N__24315\ : std_logic;
signal \N__24312\ : std_logic;
signal \N__24309\ : std_logic;
signal \N__24306\ : std_logic;
signal \N__24303\ : std_logic;
signal \N__24300\ : std_logic;
signal \N__24297\ : std_logic;
signal \N__24294\ : std_logic;
signal \N__24291\ : std_logic;
signal \N__24288\ : std_logic;
signal \N__24281\ : std_logic;
signal \N__24278\ : std_logic;
signal \N__24275\ : std_logic;
signal \N__24270\ : std_logic;
signal \N__24269\ : std_logic;
signal \N__24266\ : std_logic;
signal \N__24263\ : std_logic;
signal \N__24260\ : std_logic;
signal \N__24257\ : std_logic;
signal \N__24252\ : std_logic;
signal \N__24249\ : std_logic;
signal \N__24246\ : std_logic;
signal \N__24241\ : std_logic;
signal \N__24238\ : std_logic;
signal \N__24235\ : std_logic;
signal \N__24232\ : std_logic;
signal \N__24227\ : std_logic;
signal \N__24220\ : std_logic;
signal \N__24217\ : std_logic;
signal \N__24210\ : std_logic;
signal \N__24205\ : std_logic;
signal \N__24194\ : std_logic;
signal \N__24191\ : std_logic;
signal \N__24188\ : std_logic;
signal \N__24185\ : std_logic;
signal \N__24182\ : std_logic;
signal \N__24179\ : std_logic;
signal \N__24176\ : std_logic;
signal \N__24173\ : std_logic;
signal \N__24170\ : std_logic;
signal \N__24169\ : std_logic;
signal \N__24168\ : std_logic;
signal \N__24167\ : std_logic;
signal \N__24166\ : std_logic;
signal \N__24165\ : std_logic;
signal \N__24164\ : std_logic;
signal \N__24163\ : std_logic;
signal \N__24162\ : std_logic;
signal \N__24161\ : std_logic;
signal \N__24160\ : std_logic;
signal \N__24159\ : std_logic;
signal \N__24158\ : std_logic;
signal \N__24157\ : std_logic;
signal \N__24156\ : std_logic;
signal \N__24155\ : std_logic;
signal \N__24154\ : std_logic;
signal \N__24153\ : std_logic;
signal \N__24152\ : std_logic;
signal \N__24149\ : std_logic;
signal \N__24148\ : std_logic;
signal \N__24147\ : std_logic;
signal \N__24146\ : std_logic;
signal \N__24145\ : std_logic;
signal \N__24144\ : std_logic;
signal \N__24143\ : std_logic;
signal \N__24142\ : std_logic;
signal \N__24141\ : std_logic;
signal \N__24140\ : std_logic;
signal \N__24139\ : std_logic;
signal \N__24138\ : std_logic;
signal \N__24137\ : std_logic;
signal \N__24136\ : std_logic;
signal \N__24135\ : std_logic;
signal \N__24134\ : std_logic;
signal \N__24133\ : std_logic;
signal \N__24132\ : std_logic;
signal \N__24131\ : std_logic;
signal \N__24130\ : std_logic;
signal \N__24129\ : std_logic;
signal \N__24128\ : std_logic;
signal \N__24127\ : std_logic;
signal \N__24126\ : std_logic;
signal \N__24125\ : std_logic;
signal \N__24124\ : std_logic;
signal \N__24123\ : std_logic;
signal \N__24122\ : std_logic;
signal \N__24121\ : std_logic;
signal \N__24120\ : std_logic;
signal \N__24119\ : std_logic;
signal \N__24118\ : std_logic;
signal \N__24117\ : std_logic;
signal \N__24116\ : std_logic;
signal \N__24115\ : std_logic;
signal \N__24114\ : std_logic;
signal \N__24113\ : std_logic;
signal \N__24112\ : std_logic;
signal \N__24111\ : std_logic;
signal \N__24110\ : std_logic;
signal \N__24109\ : std_logic;
signal \N__24108\ : std_logic;
signal \N__24107\ : std_logic;
signal \N__24106\ : std_logic;
signal \N__24105\ : std_logic;
signal \N__24104\ : std_logic;
signal \N__24103\ : std_logic;
signal \N__24102\ : std_logic;
signal \N__24101\ : std_logic;
signal \N__24100\ : std_logic;
signal \N__24099\ : std_logic;
signal \N__24098\ : std_logic;
signal \N__23957\ : std_logic;
signal \N__23954\ : std_logic;
signal \N__23951\ : std_logic;
signal \N__23950\ : std_logic;
signal \N__23949\ : std_logic;
signal \N__23948\ : std_logic;
signal \N__23945\ : std_logic;
signal \N__23944\ : std_logic;
signal \N__23941\ : std_logic;
signal \N__23940\ : std_logic;
signal \N__23939\ : std_logic;
signal \N__23938\ : std_logic;
signal \N__23937\ : std_logic;
signal \N__23934\ : std_logic;
signal \N__23933\ : std_logic;
signal \N__23932\ : std_logic;
signal \N__23929\ : std_logic;
signal \N__23926\ : std_logic;
signal \N__23923\ : std_logic;
signal \N__23920\ : std_logic;
signal \N__23919\ : std_logic;
signal \N__23918\ : std_logic;
signal \N__23917\ : std_logic;
signal \N__23914\ : std_logic;
signal \N__23911\ : std_logic;
signal \N__23908\ : std_logic;
signal \N__23905\ : std_logic;
signal \N__23902\ : std_logic;
signal \N__23899\ : std_logic;
signal \N__23896\ : std_logic;
signal \N__23891\ : std_logic;
signal \N__23886\ : std_logic;
signal \N__23883\ : std_logic;
signal \N__23880\ : std_logic;
signal \N__23877\ : std_logic;
signal \N__23874\ : std_logic;
signal \N__23871\ : std_logic;
signal \N__23864\ : std_logic;
signal \N__23861\ : std_logic;
signal \N__23856\ : std_logic;
signal \N__23853\ : std_logic;
signal \N__23850\ : std_logic;
signal \N__23847\ : std_logic;
signal \N__23844\ : std_logic;
signal \N__23839\ : std_logic;
signal \N__23836\ : std_logic;
signal \N__23827\ : std_logic;
signal \N__23822\ : std_logic;
signal \N__23813\ : std_logic;
signal \N__23810\ : std_logic;
signal \N__23807\ : std_logic;
signal \N__23804\ : std_logic;
signal \N__23801\ : std_logic;
signal \N__23798\ : std_logic;
signal \N__23795\ : std_logic;
signal \N__23792\ : std_logic;
signal \N__23791\ : std_logic;
signal \N__23790\ : std_logic;
signal \N__23787\ : std_logic;
signal \N__23784\ : std_logic;
signal \N__23781\ : std_logic;
signal \N__23778\ : std_logic;
signal \N__23775\ : std_logic;
signal \N__23772\ : std_logic;
signal \N__23769\ : std_logic;
signal \N__23766\ : std_logic;
signal \N__23763\ : std_logic;
signal \N__23760\ : std_logic;
signal \N__23757\ : std_logic;
signal \N__23754\ : std_logic;
signal \N__23751\ : std_logic;
signal \N__23748\ : std_logic;
signal \N__23745\ : std_logic;
signal \N__23738\ : std_logic;
signal \N__23735\ : std_logic;
signal \N__23734\ : std_logic;
signal \N__23731\ : std_logic;
signal \N__23730\ : std_logic;
signal \N__23729\ : std_logic;
signal \N__23728\ : std_logic;
signal \N__23725\ : std_logic;
signal \N__23724\ : std_logic;
signal \N__23723\ : std_logic;
signal \N__23722\ : std_logic;
signal \N__23719\ : std_logic;
signal \N__23716\ : std_logic;
signal \N__23715\ : std_logic;
signal \N__23714\ : std_logic;
signal \N__23711\ : std_logic;
signal \N__23710\ : std_logic;
signal \N__23709\ : std_logic;
signal \N__23708\ : std_logic;
signal \N__23705\ : std_logic;
signal \N__23704\ : std_logic;
signal \N__23703\ : std_logic;
signal \N__23700\ : std_logic;
signal \N__23697\ : std_logic;
signal \N__23696\ : std_logic;
signal \N__23693\ : std_logic;
signal \N__23690\ : std_logic;
signal \N__23689\ : std_logic;
signal \N__23688\ : std_logic;
signal \N__23687\ : std_logic;
signal \N__23686\ : std_logic;
signal \N__23681\ : std_logic;
signal \N__23678\ : std_logic;
signal \N__23677\ : std_logic;
signal \N__23674\ : std_logic;
signal \N__23671\ : std_logic;
signal \N__23668\ : std_logic;
signal \N__23667\ : std_logic;
signal \N__23666\ : std_logic;
signal \N__23663\ : std_logic;
signal \N__23660\ : std_logic;
signal \N__23657\ : std_logic;
signal \N__23656\ : std_logic;
signal \N__23653\ : std_logic;
signal \N__23650\ : std_logic;
signal \N__23649\ : std_logic;
signal \N__23648\ : std_logic;
signal \N__23647\ : std_logic;
signal \N__23646\ : std_logic;
signal \N__23641\ : std_logic;
signal \N__23638\ : std_logic;
signal \N__23637\ : std_logic;
signal \N__23636\ : std_logic;
signal \N__23635\ : std_logic;
signal \N__23634\ : std_logic;
signal \N__23631\ : std_logic;
signal \N__23628\ : std_logic;
signal \N__23625\ : std_logic;
signal \N__23622\ : std_logic;
signal \N__23621\ : std_logic;
signal \N__23620\ : std_logic;
signal \N__23617\ : std_logic;
signal \N__23614\ : std_logic;
signal \N__23613\ : std_logic;
signal \N__23608\ : std_logic;
signal \N__23605\ : std_logic;
signal \N__23604\ : std_logic;
signal \N__23603\ : std_logic;
signal \N__23602\ : std_logic;
signal \N__23601\ : std_logic;
signal \N__23600\ : std_logic;
signal \N__23599\ : std_logic;
signal \N__23598\ : std_logic;
signal \N__23595\ : std_logic;
signal \N__23590\ : std_logic;
signal \N__23587\ : std_logic;
signal \N__23584\ : std_logic;
signal \N__23581\ : std_logic;
signal \N__23578\ : std_logic;
signal \N__23575\ : std_logic;
signal \N__23572\ : std_logic;
signal \N__23571\ : std_logic;
signal \N__23570\ : std_logic;
signal \N__23567\ : std_logic;
signal \N__23564\ : std_logic;
signal \N__23561\ : std_logic;
signal \N__23560\ : std_logic;
signal \N__23557\ : std_logic;
signal \N__23554\ : std_logic;
signal \N__23553\ : std_logic;
signal \N__23552\ : std_logic;
signal \N__23551\ : std_logic;
signal \N__23550\ : std_logic;
signal \N__23547\ : std_logic;
signal \N__23542\ : std_logic;
signal \N__23539\ : std_logic;
signal \N__23536\ : std_logic;
signal \N__23533\ : std_logic;
signal \N__23532\ : std_logic;
signal \N__23531\ : std_logic;
signal \N__23528\ : std_logic;
signal \N__23527\ : std_logic;
signal \N__23520\ : std_logic;
signal \N__23517\ : std_logic;
signal \N__23514\ : std_logic;
signal \N__23511\ : std_logic;
signal \N__23510\ : std_logic;
signal \N__23509\ : std_logic;
signal \N__23506\ : std_logic;
signal \N__23503\ : std_logic;
signal \N__23500\ : std_logic;
signal \N__23495\ : std_logic;
signal \N__23492\ : std_logic;
signal \N__23489\ : std_logic;
signal \N__23488\ : std_logic;
signal \N__23487\ : std_logic;
signal \N__23486\ : std_logic;
signal \N__23483\ : std_logic;
signal \N__23482\ : std_logic;
signal \N__23479\ : std_logic;
signal \N__23478\ : std_logic;
signal \N__23475\ : std_logic;
signal \N__23474\ : std_logic;
signal \N__23471\ : std_logic;
signal \N__23468\ : std_logic;
signal \N__23467\ : std_logic;
signal \N__23466\ : std_logic;
signal \N__23457\ : std_logic;
signal \N__23452\ : std_logic;
signal \N__23447\ : std_logic;
signal \N__23444\ : std_logic;
signal \N__23441\ : std_logic;
signal \N__23440\ : std_logic;
signal \N__23439\ : std_logic;
signal \N__23436\ : std_logic;
signal \N__23431\ : std_logic;
signal \N__23428\ : std_logic;
signal \N__23425\ : std_logic;
signal \N__23422\ : std_logic;
signal \N__23419\ : std_logic;
signal \N__23418\ : std_logic;
signal \N__23417\ : std_logic;
signal \N__23414\ : std_logic;
signal \N__23413\ : std_logic;
signal \N__23410\ : std_logic;
signal \N__23409\ : std_logic;
signal \N__23406\ : std_logic;
signal \N__23405\ : std_logic;
signal \N__23404\ : std_logic;
signal \N__23403\ : std_logic;
signal \N__23400\ : std_logic;
signal \N__23395\ : std_logic;
signal \N__23390\ : std_logic;
signal \N__23387\ : std_logic;
signal \N__23384\ : std_logic;
signal \N__23383\ : std_logic;
signal \N__23380\ : std_logic;
signal \N__23377\ : std_logic;
signal \N__23376\ : std_logic;
signal \N__23375\ : std_logic;
signal \N__23368\ : std_logic;
signal \N__23365\ : std_logic;
signal \N__23362\ : std_logic;
signal \N__23359\ : std_logic;
signal \N__23358\ : std_logic;
signal \N__23357\ : std_logic;
signal \N__23350\ : std_logic;
signal \N__23343\ : std_logic;
signal \N__23340\ : std_logic;
signal \N__23337\ : std_logic;
signal \N__23336\ : std_logic;
signal \N__23335\ : std_logic;
signal \N__23332\ : std_logic;
signal \N__23331\ : std_logic;
signal \N__23328\ : std_logic;
signal \N__23325\ : std_logic;
signal \N__23324\ : std_logic;
signal \N__23321\ : std_logic;
signal \N__23318\ : std_logic;
signal \N__23315\ : std_logic;
signal \N__23312\ : std_logic;
signal \N__23309\ : std_logic;
signal \N__23306\ : std_logic;
signal \N__23303\ : std_logic;
signal \N__23302\ : std_logic;
signal \N__23299\ : std_logic;
signal \N__23298\ : std_logic;
signal \N__23295\ : std_logic;
signal \N__23288\ : std_logic;
signal \N__23285\ : std_logic;
signal \N__23282\ : std_logic;
signal \N__23279\ : std_logic;
signal \N__23278\ : std_logic;
signal \N__23271\ : std_logic;
signal \N__23264\ : std_logic;
signal \N__23261\ : std_logic;
signal \N__23258\ : std_logic;
signal \N__23257\ : std_logic;
signal \N__23254\ : std_logic;
signal \N__23253\ : std_logic;
signal \N__23250\ : std_logic;
signal \N__23249\ : std_logic;
signal \N__23248\ : std_logic;
signal \N__23245\ : std_logic;
signal \N__23242\ : std_logic;
signal \N__23239\ : std_logic;
signal \N__23236\ : std_logic;
signal \N__23233\ : std_logic;
signal \N__23232\ : std_logic;
signal \N__23229\ : std_logic;
signal \N__23228\ : std_logic;
signal \N__23227\ : std_logic;
signal \N__23216\ : std_logic;
signal \N__23213\ : std_logic;
signal \N__23208\ : std_logic;
signal \N__23205\ : std_logic;
signal \N__23202\ : std_logic;
signal \N__23201\ : std_logic;
signal \N__23194\ : std_logic;
signal \N__23191\ : std_logic;
signal \N__23188\ : std_logic;
signal \N__23185\ : std_logic;
signal \N__23184\ : std_logic;
signal \N__23177\ : std_logic;
signal \N__23174\ : std_logic;
signal \N__23171\ : std_logic;
signal \N__23168\ : std_logic;
signal \N__23165\ : std_logic;
signal \N__23162\ : std_logic;
signal \N__23157\ : std_logic;
signal \N__23154\ : std_logic;
signal \N__23149\ : std_logic;
signal \N__23144\ : std_logic;
signal \N__23137\ : std_logic;
signal \N__23134\ : std_logic;
signal \N__23133\ : std_logic;
signal \N__23132\ : std_logic;
signal \N__23129\ : std_logic;
signal \N__23126\ : std_logic;
signal \N__23125\ : std_logic;
signal \N__23118\ : std_logic;
signal \N__23115\ : std_logic;
signal \N__23112\ : std_logic;
signal \N__23109\ : std_logic;
signal \N__23106\ : std_logic;
signal \N__23099\ : std_logic;
signal \N__23096\ : std_logic;
signal \N__23093\ : std_logic;
signal \N__23090\ : std_logic;
signal \N__23087\ : std_logic;
signal \N__23084\ : std_logic;
signal \N__23083\ : std_logic;
signal \N__23080\ : std_logic;
signal \N__23075\ : std_logic;
signal \N__23068\ : std_logic;
signal \N__23065\ : std_logic;
signal \N__23062\ : std_logic;
signal \N__23059\ : std_logic;
signal \N__23056\ : std_logic;
signal \N__23051\ : std_logic;
signal \N__23046\ : std_logic;
signal \N__23043\ : std_logic;
signal \N__23040\ : std_logic;
signal \N__23039\ : std_logic;
signal \N__23038\ : std_logic;
signal \N__23037\ : std_logic;
signal \N__23030\ : std_logic;
signal \N__23027\ : std_logic;
signal \N__23024\ : std_logic;
signal \N__23023\ : std_logic;
signal \N__23020\ : std_logic;
signal \N__23015\ : std_logic;
signal \N__23012\ : std_logic;
signal \N__23003\ : std_logic;
signal \N__22994\ : std_logic;
signal \N__22991\ : std_logic;
signal \N__22988\ : std_logic;
signal \N__22987\ : std_logic;
signal \N__22982\ : std_logic;
signal \N__22979\ : std_logic;
signal \N__22972\ : std_logic;
signal \N__22969\ : std_logic;
signal \N__22964\ : std_logic;
signal \N__22961\ : std_logic;
signal \N__22956\ : std_logic;
signal \N__22955\ : std_logic;
signal \N__22952\ : std_logic;
signal \N__22949\ : std_logic;
signal \N__22946\ : std_logic;
signal \N__22943\ : std_logic;
signal \N__22936\ : std_logic;
signal \N__22931\ : std_logic;
signal \N__22928\ : std_logic;
signal \N__22919\ : std_logic;
signal \N__22916\ : std_logic;
signal \N__22913\ : std_logic;
signal \N__22912\ : std_logic;
signal \N__22909\ : std_logic;
signal \N__22908\ : std_logic;
signal \N__22901\ : std_logic;
signal \N__22898\ : std_logic;
signal \N__22895\ : std_logic;
signal \N__22892\ : std_logic;
signal \N__22887\ : std_logic;
signal \N__22880\ : std_logic;
signal \N__22877\ : std_logic;
signal \N__22876\ : std_logic;
signal \N__22873\ : std_logic;
signal \N__22870\ : std_logic;
signal \N__22869\ : std_logic;
signal \N__22866\ : std_logic;
signal \N__22863\ : std_logic;
signal \N__22858\ : std_logic;
signal \N__22855\ : std_logic;
signal \N__22852\ : std_logic;
signal \N__22847\ : std_logic;
signal \N__22844\ : std_logic;
signal \N__22841\ : std_logic;
signal \N__22830\ : std_logic;
signal \N__22827\ : std_logic;
signal \N__22824\ : std_logic;
signal \N__22821\ : std_logic;
signal \N__22818\ : std_logic;
signal \N__22815\ : std_logic;
signal \N__22812\ : std_logic;
signal \N__22807\ : std_logic;
signal \N__22800\ : std_logic;
signal \N__22797\ : std_logic;
signal \N__22792\ : std_logic;
signal \N__22789\ : std_logic;
signal \N__22786\ : std_logic;
signal \N__22783\ : std_logic;
signal \N__22780\ : std_logic;
signal \N__22777\ : std_logic;
signal \N__22774\ : std_logic;
signal \N__22771\ : std_logic;
signal \N__22768\ : std_logic;
signal \N__22761\ : std_logic;
signal \N__22758\ : std_logic;
signal \N__22753\ : std_logic;
signal \N__22746\ : std_logic;
signal \N__22737\ : std_logic;
signal \N__22732\ : std_logic;
signal \N__22729\ : std_logic;
signal \N__22726\ : std_logic;
signal \N__22723\ : std_logic;
signal \N__22716\ : std_logic;
signal \N__22707\ : std_logic;
signal \N__22694\ : std_logic;
signal \N__22693\ : std_logic;
signal \N__22692\ : std_logic;
signal \N__22689\ : std_logic;
signal \N__22688\ : std_logic;
signal \N__22687\ : std_logic;
signal \N__22684\ : std_logic;
signal \N__22681\ : std_logic;
signal \N__22680\ : std_logic;
signal \N__22677\ : std_logic;
signal \N__22674\ : std_logic;
signal \N__22671\ : std_logic;
signal \N__22670\ : std_logic;
signal \N__22667\ : std_logic;
signal \N__22664\ : std_logic;
signal \N__22661\ : std_logic;
signal \N__22656\ : std_logic;
signal \N__22653\ : std_logic;
signal \N__22650\ : std_logic;
signal \N__22649\ : std_logic;
signal \N__22646\ : std_logic;
signal \N__22641\ : std_logic;
signal \N__22634\ : std_logic;
signal \N__22631\ : std_logic;
signal \N__22626\ : std_logic;
signal \N__22623\ : std_logic;
signal \N__22620\ : std_logic;
signal \N__22613\ : std_logic;
signal \N__22610\ : std_logic;
signal \N__22607\ : std_logic;
signal \N__22604\ : std_logic;
signal \N__22601\ : std_logic;
signal \N__22598\ : std_logic;
signal \N__22595\ : std_logic;
signal \N__22592\ : std_logic;
signal \N__22589\ : std_logic;
signal \N__22586\ : std_logic;
signal \N__22583\ : std_logic;
signal \N__22580\ : std_logic;
signal \N__22577\ : std_logic;
signal \N__22574\ : std_logic;
signal \N__22571\ : std_logic;
signal \N__22568\ : std_logic;
signal \N__22565\ : std_logic;
signal \N__22562\ : std_logic;
signal \N__22559\ : std_logic;
signal \N__22556\ : std_logic;
signal \N__22553\ : std_logic;
signal \N__22550\ : std_logic;
signal \N__22547\ : std_logic;
signal \N__22544\ : std_logic;
signal \N__22541\ : std_logic;
signal \N__22538\ : std_logic;
signal \N__22535\ : std_logic;
signal \N__22532\ : std_logic;
signal \N__22529\ : std_logic;
signal \N__22526\ : std_logic;
signal \N__22523\ : std_logic;
signal \N__22520\ : std_logic;
signal \N__22519\ : std_logic;
signal \N__22518\ : std_logic;
signal \N__22517\ : std_logic;
signal \N__22514\ : std_logic;
signal \N__22513\ : std_logic;
signal \N__22510\ : std_logic;
signal \N__22507\ : std_logic;
signal \N__22506\ : std_logic;
signal \N__22503\ : std_logic;
signal \N__22500\ : std_logic;
signal \N__22497\ : std_logic;
signal \N__22496\ : std_logic;
signal \N__22493\ : std_logic;
signal \N__22490\ : std_logic;
signal \N__22487\ : std_logic;
signal \N__22484\ : std_logic;
signal \N__22483\ : std_logic;
signal \N__22478\ : std_logic;
signal \N__22475\ : std_logic;
signal \N__22472\ : std_logic;
signal \N__22469\ : std_logic;
signal \N__22466\ : std_logic;
signal \N__22463\ : std_logic;
signal \N__22460\ : std_logic;
signal \N__22457\ : std_logic;
signal \N__22456\ : std_logic;
signal \N__22453\ : std_logic;
signal \N__22450\ : std_logic;
signal \N__22445\ : std_logic;
signal \N__22440\ : std_logic;
signal \N__22437\ : std_logic;
signal \N__22434\ : std_logic;
signal \N__22431\ : std_logic;
signal \N__22428\ : std_logic;
signal \N__22423\ : std_logic;
signal \N__22418\ : std_logic;
signal \N__22409\ : std_logic;
signal \N__22406\ : std_logic;
signal \N__22403\ : std_logic;
signal \N__22400\ : std_logic;
signal \N__22397\ : std_logic;
signal \N__22394\ : std_logic;
signal \N__22393\ : std_logic;
signal \N__22392\ : std_logic;
signal \N__22391\ : std_logic;
signal \N__22390\ : std_logic;
signal \N__22389\ : std_logic;
signal \N__22388\ : std_logic;
signal \N__22385\ : std_logic;
signal \N__22382\ : std_logic;
signal \N__22381\ : std_logic;
signal \N__22378\ : std_logic;
signal \N__22377\ : std_logic;
signal \N__22376\ : std_logic;
signal \N__22375\ : std_logic;
signal \N__22374\ : std_logic;
signal \N__22373\ : std_logic;
signal \N__22372\ : std_logic;
signal \N__22369\ : std_logic;
signal \N__22366\ : std_logic;
signal \N__22363\ : std_logic;
signal \N__22360\ : std_logic;
signal \N__22357\ : std_logic;
signal \N__22354\ : std_logic;
signal \N__22351\ : std_logic;
signal \N__22350\ : std_logic;
signal \N__22347\ : std_logic;
signal \N__22346\ : std_logic;
signal \N__22343\ : std_logic;
signal \N__22340\ : std_logic;
signal \N__22339\ : std_logic;
signal \N__22338\ : std_logic;
signal \N__22337\ : std_logic;
signal \N__22334\ : std_logic;
signal \N__22331\ : std_logic;
signal \N__22328\ : std_logic;
signal \N__22325\ : std_logic;
signal \N__22322\ : std_logic;
signal \N__22313\ : std_logic;
signal \N__22310\ : std_logic;
signal \N__22307\ : std_logic;
signal \N__22306\ : std_logic;
signal \N__22305\ : std_logic;
signal \N__22302\ : std_logic;
signal \N__22299\ : std_logic;
signal \N__22296\ : std_logic;
signal \N__22293\ : std_logic;
signal \N__22290\ : std_logic;
signal \N__22287\ : std_logic;
signal \N__22284\ : std_logic;
signal \N__22281\ : std_logic;
signal \N__22276\ : std_logic;
signal \N__22273\ : std_logic;
signal \N__22270\ : std_logic;
signal \N__22269\ : std_logic;
signal \N__22260\ : std_logic;
signal \N__22257\ : std_logic;
signal \N__22254\ : std_logic;
signal \N__22249\ : std_logic;
signal \N__22242\ : std_logic;
signal \N__22229\ : std_logic;
signal \N__22226\ : std_logic;
signal \N__22223\ : std_logic;
signal \N__22220\ : std_logic;
signal \N__22211\ : std_logic;
signal \N__22208\ : std_logic;
signal \N__22205\ : std_logic;
signal \N__22200\ : std_logic;
signal \N__22193\ : std_logic;
signal \N__22190\ : std_logic;
signal \N__22187\ : std_logic;
signal \N__22184\ : std_logic;
signal \N__22181\ : std_logic;
signal \N__22178\ : std_logic;
signal \N__22175\ : std_logic;
signal \N__22172\ : std_logic;
signal \N__22169\ : std_logic;
signal \N__22166\ : std_logic;
signal \N__22165\ : std_logic;
signal \N__22162\ : std_logic;
signal \N__22159\ : std_logic;
signal \N__22156\ : std_logic;
signal \N__22153\ : std_logic;
signal \N__22150\ : std_logic;
signal \N__22147\ : std_logic;
signal \N__22144\ : std_logic;
signal \N__22141\ : std_logic;
signal \N__22138\ : std_logic;
signal \N__22135\ : std_logic;
signal \N__22132\ : std_logic;
signal \N__22129\ : std_logic;
signal \N__22124\ : std_logic;
signal \N__22121\ : std_logic;
signal \N__22118\ : std_logic;
signal \N__22115\ : std_logic;
signal \N__22112\ : std_logic;
signal \N__22109\ : std_logic;
signal \N__22106\ : std_logic;
signal \N__22103\ : std_logic;
signal \N__22100\ : std_logic;
signal \N__22097\ : std_logic;
signal \N__22094\ : std_logic;
signal \N__22091\ : std_logic;
signal \N__22088\ : std_logic;
signal \N__22085\ : std_logic;
signal \N__22082\ : std_logic;
signal \N__22079\ : std_logic;
signal \N__22076\ : std_logic;
signal \N__22073\ : std_logic;
signal \N__22070\ : std_logic;
signal \N__22067\ : std_logic;
signal \N__22064\ : std_logic;
signal \N__22061\ : std_logic;
signal \N__22058\ : std_logic;
signal \N__22055\ : std_logic;
signal \N__22052\ : std_logic;
signal \N__22049\ : std_logic;
signal \N__22046\ : std_logic;
signal \N__22043\ : std_logic;
signal \N__22040\ : std_logic;
signal \N__22037\ : std_logic;
signal \N__22034\ : std_logic;
signal \N__22031\ : std_logic;
signal \N__22028\ : std_logic;
signal \N__22025\ : std_logic;
signal \N__22022\ : std_logic;
signal \N__22019\ : std_logic;
signal \N__22016\ : std_logic;
signal \N__22013\ : std_logic;
signal \N__22010\ : std_logic;
signal \N__22007\ : std_logic;
signal \N__22004\ : std_logic;
signal \N__22001\ : std_logic;
signal \N__21998\ : std_logic;
signal \N__21995\ : std_logic;
signal \N__21994\ : std_logic;
signal \N__21991\ : std_logic;
signal \N__21988\ : std_logic;
signal \N__21985\ : std_logic;
signal \N__21984\ : std_logic;
signal \N__21981\ : std_logic;
signal \N__21978\ : std_logic;
signal \N__21975\ : std_logic;
signal \N__21972\ : std_logic;
signal \N__21969\ : std_logic;
signal \N__21966\ : std_logic;
signal \N__21963\ : std_logic;
signal \N__21960\ : std_logic;
signal \N__21955\ : std_logic;
signal \N__21950\ : std_logic;
signal \N__21947\ : std_logic;
signal \N__21944\ : std_logic;
signal \N__21941\ : std_logic;
signal \N__21938\ : std_logic;
signal \N__21935\ : std_logic;
signal \N__21932\ : std_logic;
signal \N__21929\ : std_logic;
signal \N__21926\ : std_logic;
signal \N__21923\ : std_logic;
signal \N__21920\ : std_logic;
signal \N__21917\ : std_logic;
signal \N__21914\ : std_logic;
signal \N__21911\ : std_logic;
signal \N__21908\ : std_logic;
signal \N__21905\ : std_logic;
signal \N__21902\ : std_logic;
signal \N__21899\ : std_logic;
signal \N__21896\ : std_logic;
signal \N__21893\ : std_logic;
signal \N__21890\ : std_logic;
signal \N__21887\ : std_logic;
signal \N__21884\ : std_logic;
signal \N__21881\ : std_logic;
signal \N__21878\ : std_logic;
signal \N__21875\ : std_logic;
signal \N__21872\ : std_logic;
signal \N__21869\ : std_logic;
signal \N__21866\ : std_logic;
signal \N__21863\ : std_logic;
signal \N__21860\ : std_logic;
signal \N__21857\ : std_logic;
signal \N__21854\ : std_logic;
signal \N__21851\ : std_logic;
signal \N__21848\ : std_logic;
signal \N__21845\ : std_logic;
signal \N__21842\ : std_logic;
signal \N__21839\ : std_logic;
signal \N__21836\ : std_logic;
signal \N__21833\ : std_logic;
signal \N__21830\ : std_logic;
signal \N__21827\ : std_logic;
signal \N__21824\ : std_logic;
signal \N__21821\ : std_logic;
signal \N__21818\ : std_logic;
signal \N__21815\ : std_logic;
signal \N__21812\ : std_logic;
signal \N__21809\ : std_logic;
signal \N__21806\ : std_logic;
signal \N__21803\ : std_logic;
signal \N__21800\ : std_logic;
signal \N__21797\ : std_logic;
signal \N__21794\ : std_logic;
signal \N__21791\ : std_logic;
signal \N__21788\ : std_logic;
signal \N__21785\ : std_logic;
signal \N__21782\ : std_logic;
signal \N__21779\ : std_logic;
signal \N__21776\ : std_logic;
signal \N__21773\ : std_logic;
signal \N__21770\ : std_logic;
signal \N__21767\ : std_logic;
signal \N__21764\ : std_logic;
signal \N__21761\ : std_logic;
signal \N__21760\ : std_logic;
signal \N__21757\ : std_logic;
signal \N__21754\ : std_logic;
signal \N__21751\ : std_logic;
signal \N__21748\ : std_logic;
signal \N__21747\ : std_logic;
signal \N__21744\ : std_logic;
signal \N__21741\ : std_logic;
signal \N__21738\ : std_logic;
signal \N__21733\ : std_logic;
signal \N__21730\ : std_logic;
signal \N__21727\ : std_logic;
signal \N__21724\ : std_logic;
signal \N__21721\ : std_logic;
signal \N__21718\ : std_logic;
signal \N__21713\ : std_logic;
signal \N__21710\ : std_logic;
signal \N__21707\ : std_logic;
signal \N__21704\ : std_logic;
signal \N__21701\ : std_logic;
signal \N__21698\ : std_logic;
signal \N__21695\ : std_logic;
signal \N__21692\ : std_logic;
signal \N__21689\ : std_logic;
signal \N__21686\ : std_logic;
signal \N__21683\ : std_logic;
signal \N__21680\ : std_logic;
signal \N__21677\ : std_logic;
signal \N__21674\ : std_logic;
signal \N__21671\ : std_logic;
signal \N__21668\ : std_logic;
signal \N__21665\ : std_logic;
signal \N__21662\ : std_logic;
signal \N__21659\ : std_logic;
signal \N__21656\ : std_logic;
signal \N__21653\ : std_logic;
signal \N__21650\ : std_logic;
signal \N__21647\ : std_logic;
signal \N__21644\ : std_logic;
signal \N__21641\ : std_logic;
signal \N__21638\ : std_logic;
signal \N__21635\ : std_logic;
signal \N__21632\ : std_logic;
signal \N__21629\ : std_logic;
signal \N__21628\ : std_logic;
signal \N__21625\ : std_logic;
signal \N__21622\ : std_logic;
signal \N__21617\ : std_logic;
signal \N__21614\ : std_logic;
signal \N__21611\ : std_logic;
signal \N__21608\ : std_logic;
signal \N__21605\ : std_logic;
signal \N__21602\ : std_logic;
signal \N__21599\ : std_logic;
signal \N__21596\ : std_logic;
signal \N__21593\ : std_logic;
signal \N__21590\ : std_logic;
signal \N__21587\ : std_logic;
signal \N__21584\ : std_logic;
signal \N__21581\ : std_logic;
signal \N__21578\ : std_logic;
signal \N__21575\ : std_logic;
signal \N__21572\ : std_logic;
signal \N__21569\ : std_logic;
signal \N__21566\ : std_logic;
signal \N__21563\ : std_logic;
signal \N__21560\ : std_logic;
signal \N__21557\ : std_logic;
signal \N__21554\ : std_logic;
signal \N__21551\ : std_logic;
signal \N__21548\ : std_logic;
signal \N__21545\ : std_logic;
signal \N__21542\ : std_logic;
signal \N__21539\ : std_logic;
signal \N__21536\ : std_logic;
signal \N__21533\ : std_logic;
signal \N__21530\ : std_logic;
signal \N__21527\ : std_logic;
signal \N__21524\ : std_logic;
signal \N__21521\ : std_logic;
signal \N__21518\ : std_logic;
signal \N__21515\ : std_logic;
signal \N__21512\ : std_logic;
signal \N__21509\ : std_logic;
signal \N__21506\ : std_logic;
signal \N__21503\ : std_logic;
signal \N__21500\ : std_logic;
signal \N__21497\ : std_logic;
signal \N__21494\ : std_logic;
signal \N__21491\ : std_logic;
signal \N__21488\ : std_logic;
signal \N__21485\ : std_logic;
signal \N__21482\ : std_logic;
signal \N__21479\ : std_logic;
signal \N__21476\ : std_logic;
signal \N__21475\ : std_logic;
signal \N__21474\ : std_logic;
signal \N__21471\ : std_logic;
signal \N__21468\ : std_logic;
signal \N__21465\ : std_logic;
signal \N__21464\ : std_logic;
signal \N__21461\ : std_logic;
signal \N__21458\ : std_logic;
signal \N__21455\ : std_logic;
signal \N__21452\ : std_logic;
signal \N__21449\ : std_logic;
signal \N__21446\ : std_logic;
signal \N__21443\ : std_logic;
signal \N__21440\ : std_logic;
signal \N__21431\ : std_logic;
signal \N__21430\ : std_logic;
signal \N__21429\ : std_logic;
signal \N__21428\ : std_logic;
signal \N__21427\ : std_logic;
signal \N__21426\ : std_logic;
signal \N__21423\ : std_logic;
signal \N__21420\ : std_logic;
signal \N__21417\ : std_logic;
signal \N__21414\ : std_logic;
signal \N__21411\ : std_logic;
signal \N__21408\ : std_logic;
signal \N__21407\ : std_logic;
signal \N__21406\ : std_logic;
signal \N__21405\ : std_logic;
signal \N__21402\ : std_logic;
signal \N__21399\ : std_logic;
signal \N__21392\ : std_logic;
signal \N__21389\ : std_logic;
signal \N__21386\ : std_logic;
signal \N__21383\ : std_logic;
signal \N__21382\ : std_logic;
signal \N__21381\ : std_logic;
signal \N__21378\ : std_logic;
signal \N__21373\ : std_logic;
signal \N__21366\ : std_logic;
signal \N__21363\ : std_logic;
signal \N__21362\ : std_logic;
signal \N__21359\ : std_logic;
signal \N__21356\ : std_logic;
signal \N__21355\ : std_logic;
signal \N__21354\ : std_logic;
signal \N__21351\ : std_logic;
signal \N__21344\ : std_logic;
signal \N__21341\ : std_logic;
signal \N__21338\ : std_logic;
signal \N__21335\ : std_logic;
signal \N__21332\ : std_logic;
signal \N__21331\ : std_logic;
signal \N__21328\ : std_logic;
signal \N__21327\ : std_logic;
signal \N__21322\ : std_logic;
signal \N__21319\ : std_logic;
signal \N__21312\ : std_logic;
signal \N__21309\ : std_logic;
signal \N__21306\ : std_logic;
signal \N__21303\ : std_logic;
signal \N__21300\ : std_logic;
signal \N__21297\ : std_logic;
signal \N__21294\ : std_logic;
signal \N__21287\ : std_logic;
signal \N__21278\ : std_logic;
signal \N__21275\ : std_logic;
signal \N__21272\ : std_logic;
signal \N__21269\ : std_logic;
signal \N__21266\ : std_logic;
signal \N__21263\ : std_logic;
signal \N__21260\ : std_logic;
signal \N__21257\ : std_logic;
signal \N__21254\ : std_logic;
signal \N__21251\ : std_logic;
signal \N__21248\ : std_logic;
signal \N__21245\ : std_logic;
signal \N__21242\ : std_logic;
signal \N__21239\ : std_logic;
signal \N__21236\ : std_logic;
signal \N__21233\ : std_logic;
signal \N__21230\ : std_logic;
signal \N__21227\ : std_logic;
signal \N__21224\ : std_logic;
signal \N__21221\ : std_logic;
signal \N__21218\ : std_logic;
signal \N__21215\ : std_logic;
signal \N__21212\ : std_logic;
signal \N__21209\ : std_logic;
signal \N__21206\ : std_logic;
signal \N__21203\ : std_logic;
signal \N__21200\ : std_logic;
signal \N__21197\ : std_logic;
signal \N__21194\ : std_logic;
signal \N__21191\ : std_logic;
signal \N__21188\ : std_logic;
signal \N__21185\ : std_logic;
signal \N__21182\ : std_logic;
signal \N__21179\ : std_logic;
signal \N__21176\ : std_logic;
signal \N__21173\ : std_logic;
signal \N__21170\ : std_logic;
signal \N__21167\ : std_logic;
signal \N__21164\ : std_logic;
signal \N__21161\ : std_logic;
signal \N__21158\ : std_logic;
signal \N__21155\ : std_logic;
signal \N__21152\ : std_logic;
signal \N__21149\ : std_logic;
signal \N__21146\ : std_logic;
signal \N__21143\ : std_logic;
signal \N__21140\ : std_logic;
signal \N__21137\ : std_logic;
signal \N__21134\ : std_logic;
signal \N__21131\ : std_logic;
signal \N__21128\ : std_logic;
signal \N__21125\ : std_logic;
signal \N__21122\ : std_logic;
signal \N__21119\ : std_logic;
signal \N__21116\ : std_logic;
signal \N__21113\ : std_logic;
signal \N__21110\ : std_logic;
signal \N__21107\ : std_logic;
signal \N__21104\ : std_logic;
signal \N__21101\ : std_logic;
signal \N__21098\ : std_logic;
signal \N__21095\ : std_logic;
signal \N__21092\ : std_logic;
signal \N__21089\ : std_logic;
signal \N__21086\ : std_logic;
signal \N__21083\ : std_logic;
signal \N__21080\ : std_logic;
signal \N__21077\ : std_logic;
signal \N__21074\ : std_logic;
signal \N__21071\ : std_logic;
signal \N__21068\ : std_logic;
signal \N__21065\ : std_logic;
signal \N__21062\ : std_logic;
signal \N__21059\ : std_logic;
signal \N__21056\ : std_logic;
signal \N__21053\ : std_logic;
signal \N__21050\ : std_logic;
signal \N__21047\ : std_logic;
signal \N__21044\ : std_logic;
signal \N__21041\ : std_logic;
signal \N__21038\ : std_logic;
signal \N__21035\ : std_logic;
signal \N__21032\ : std_logic;
signal \N__21029\ : std_logic;
signal \N__21026\ : std_logic;
signal \N__21023\ : std_logic;
signal \N__21020\ : std_logic;
signal \N__21017\ : std_logic;
signal \N__21014\ : std_logic;
signal \N__21011\ : std_logic;
signal \N__21008\ : std_logic;
signal \N__21005\ : std_logic;
signal \N__21002\ : std_logic;
signal \N__20999\ : std_logic;
signal \N__20996\ : std_logic;
signal \N__20993\ : std_logic;
signal \N__20990\ : std_logic;
signal \N__20987\ : std_logic;
signal \N__20984\ : std_logic;
signal \N__20981\ : std_logic;
signal \N__20978\ : std_logic;
signal \N__20975\ : std_logic;
signal \N__20972\ : std_logic;
signal \N__20969\ : std_logic;
signal \N__20966\ : std_logic;
signal \N__20965\ : std_logic;
signal \N__20964\ : std_logic;
signal \N__20961\ : std_logic;
signal \N__20958\ : std_logic;
signal \N__20955\ : std_logic;
signal \N__20952\ : std_logic;
signal \N__20949\ : std_logic;
signal \N__20946\ : std_logic;
signal \N__20943\ : std_logic;
signal \N__20940\ : std_logic;
signal \N__20937\ : std_logic;
signal \N__20934\ : std_logic;
signal \N__20931\ : std_logic;
signal \N__20928\ : std_logic;
signal \N__20923\ : std_logic;
signal \N__20920\ : std_logic;
signal \N__20917\ : std_logic;
signal \N__20914\ : std_logic;
signal \N__20911\ : std_logic;
signal \N__20906\ : std_logic;
signal \N__20903\ : std_logic;
signal \N__20900\ : std_logic;
signal \N__20897\ : std_logic;
signal \N__20894\ : std_logic;
signal \N__20891\ : std_logic;
signal \N__20890\ : std_logic;
signal \N__20887\ : std_logic;
signal \N__20884\ : std_logic;
signal \N__20879\ : std_logic;
signal \N__20876\ : std_logic;
signal \N__20875\ : std_logic;
signal \N__20872\ : std_logic;
signal \N__20869\ : std_logic;
signal \N__20866\ : std_logic;
signal \N__20863\ : std_logic;
signal \N__20860\ : std_logic;
signal \N__20857\ : std_logic;
signal \N__20852\ : std_logic;
signal \N__20849\ : std_logic;
signal \N__20846\ : std_logic;
signal \N__20843\ : std_logic;
signal \N__20840\ : std_logic;
signal \N__20837\ : std_logic;
signal \N__20834\ : std_logic;
signal \N__20831\ : std_logic;
signal \N__20828\ : std_logic;
signal \N__20825\ : std_logic;
signal \N__20822\ : std_logic;
signal \N__20819\ : std_logic;
signal \N__20816\ : std_logic;
signal \N__20813\ : std_logic;
signal \N__20810\ : std_logic;
signal \N__20807\ : std_logic;
signal \N__20806\ : std_logic;
signal \N__20805\ : std_logic;
signal \N__20804\ : std_logic;
signal \N__20801\ : std_logic;
signal \N__20798\ : std_logic;
signal \N__20795\ : std_logic;
signal \N__20792\ : std_logic;
signal \N__20783\ : std_logic;
signal \N__20780\ : std_logic;
signal \N__20777\ : std_logic;
signal \N__20774\ : std_logic;
signal \N__20773\ : std_logic;
signal \N__20772\ : std_logic;
signal \N__20771\ : std_logic;
signal \N__20768\ : std_logic;
signal \N__20765\ : std_logic;
signal \N__20764\ : std_logic;
signal \N__20761\ : std_logic;
signal \N__20758\ : std_logic;
signal \N__20757\ : std_logic;
signal \N__20752\ : std_logic;
signal \N__20749\ : std_logic;
signal \N__20748\ : std_logic;
signal \N__20745\ : std_logic;
signal \N__20742\ : std_logic;
signal \N__20739\ : std_logic;
signal \N__20738\ : std_logic;
signal \N__20735\ : std_logic;
signal \N__20732\ : std_logic;
signal \N__20729\ : std_logic;
signal \N__20724\ : std_logic;
signal \N__20721\ : std_logic;
signal \N__20718\ : std_logic;
signal \N__20713\ : std_logic;
signal \N__20710\ : std_logic;
signal \N__20707\ : std_logic;
signal \N__20704\ : std_logic;
signal \N__20701\ : std_logic;
signal \N__20690\ : std_logic;
signal \N__20687\ : std_logic;
signal \N__20684\ : std_logic;
signal \N__20683\ : std_logic;
signal \N__20682\ : std_logic;
signal \N__20679\ : std_logic;
signal \N__20678\ : std_logic;
signal \N__20677\ : std_logic;
signal \N__20676\ : std_logic;
signal \N__20673\ : std_logic;
signal \N__20672\ : std_logic;
signal \N__20671\ : std_logic;
signal \N__20668\ : std_logic;
signal \N__20665\ : std_logic;
signal \N__20662\ : std_logic;
signal \N__20661\ : std_logic;
signal \N__20656\ : std_logic;
signal \N__20655\ : std_logic;
signal \N__20652\ : std_logic;
signal \N__20649\ : std_logic;
signal \N__20648\ : std_logic;
signal \N__20647\ : std_logic;
signal \N__20644\ : std_logic;
signal \N__20641\ : std_logic;
signal \N__20636\ : std_logic;
signal \N__20633\ : std_logic;
signal \N__20630\ : std_logic;
signal \N__20627\ : std_logic;
signal \N__20626\ : std_logic;
signal \N__20625\ : std_logic;
signal \N__20620\ : std_logic;
signal \N__20615\ : std_logic;
signal \N__20612\ : std_logic;
signal \N__20605\ : std_logic;
signal \N__20600\ : std_logic;
signal \N__20597\ : std_logic;
signal \N__20594\ : std_logic;
signal \N__20579\ : std_logic;
signal \N__20578\ : std_logic;
signal \N__20577\ : std_logic;
signal \N__20574\ : std_logic;
signal \N__20573\ : std_logic;
signal \N__20570\ : std_logic;
signal \N__20567\ : std_logic;
signal \N__20564\ : std_logic;
signal \N__20561\ : std_logic;
signal \N__20552\ : std_logic;
signal \N__20549\ : std_logic;
signal \N__20548\ : std_logic;
signal \N__20545\ : std_logic;
signal \N__20542\ : std_logic;
signal \N__20537\ : std_logic;
signal \N__20534\ : std_logic;
signal \N__20531\ : std_logic;
signal \N__20528\ : std_logic;
signal \N__20527\ : std_logic;
signal \N__20524\ : std_logic;
signal \N__20521\ : std_logic;
signal \N__20518\ : std_logic;
signal \N__20515\ : std_logic;
signal \N__20512\ : std_logic;
signal \N__20509\ : std_logic;
signal \N__20506\ : std_logic;
signal \N__20503\ : std_logic;
signal \N__20500\ : std_logic;
signal \N__20497\ : std_logic;
signal \N__20494\ : std_logic;
signal \N__20491\ : std_logic;
signal \N__20488\ : std_logic;
signal \N__20485\ : std_logic;
signal \N__20482\ : std_logic;
signal \N__20479\ : std_logic;
signal \N__20476\ : std_logic;
signal \N__20473\ : std_logic;
signal \N__20470\ : std_logic;
signal \N__20467\ : std_logic;
signal \N__20464\ : std_logic;
signal \N__20461\ : std_logic;
signal \N__20458\ : std_logic;
signal \N__20455\ : std_logic;
signal \N__20452\ : std_logic;
signal \N__20449\ : std_logic;
signal \N__20446\ : std_logic;
signal \N__20443\ : std_logic;
signal \N__20440\ : std_logic;
signal \N__20437\ : std_logic;
signal \N__20434\ : std_logic;
signal \N__20431\ : std_logic;
signal \N__20428\ : std_logic;
signal \N__20425\ : std_logic;
signal \N__20422\ : std_logic;
signal \N__20419\ : std_logic;
signal \N__20416\ : std_logic;
signal \N__20413\ : std_logic;
signal \N__20410\ : std_logic;
signal \N__20407\ : std_logic;
signal \N__20404\ : std_logic;
signal \N__20401\ : std_logic;
signal \N__20398\ : std_logic;
signal \N__20395\ : std_logic;
signal \N__20392\ : std_logic;
signal \N__20389\ : std_logic;
signal \N__20386\ : std_logic;
signal \N__20383\ : std_logic;
signal \N__20380\ : std_logic;
signal \N__20377\ : std_logic;
signal \N__20374\ : std_logic;
signal \N__20371\ : std_logic;
signal \N__20368\ : std_logic;
signal \N__20365\ : std_logic;
signal \N__20362\ : std_logic;
signal \N__20359\ : std_logic;
signal \N__20356\ : std_logic;
signal \N__20353\ : std_logic;
signal \N__20350\ : std_logic;
signal \N__20347\ : std_logic;
signal \N__20344\ : std_logic;
signal \N__20341\ : std_logic;
signal \N__20338\ : std_logic;
signal \N__20335\ : std_logic;
signal \N__20332\ : std_logic;
signal \N__20329\ : std_logic;
signal \N__20326\ : std_logic;
signal \N__20323\ : std_logic;
signal \N__20320\ : std_logic;
signal \N__20317\ : std_logic;
signal \N__20314\ : std_logic;
signal \N__20309\ : std_logic;
signal \N__20306\ : std_logic;
signal \N__20303\ : std_logic;
signal \N__20300\ : std_logic;
signal \N__20297\ : std_logic;
signal \N__20294\ : std_logic;
signal \N__20291\ : std_logic;
signal \N__20288\ : std_logic;
signal \N__20285\ : std_logic;
signal \N__20282\ : std_logic;
signal \N__20279\ : std_logic;
signal \N__20276\ : std_logic;
signal \N__20273\ : std_logic;
signal \N__20270\ : std_logic;
signal \N__20267\ : std_logic;
signal \N__20264\ : std_logic;
signal \N__20263\ : std_logic;
signal \N__20262\ : std_logic;
signal \N__20261\ : std_logic;
signal \N__20260\ : std_logic;
signal \N__20259\ : std_logic;
signal \N__20258\ : std_logic;
signal \N__20257\ : std_logic;
signal \N__20256\ : std_logic;
signal \N__20255\ : std_logic;
signal \N__20254\ : std_logic;
signal \N__20253\ : std_logic;
signal \N__20252\ : std_logic;
signal \N__20251\ : std_logic;
signal \N__20248\ : std_logic;
signal \N__20243\ : std_logic;
signal \N__20240\ : std_logic;
signal \N__20237\ : std_logic;
signal \N__20236\ : std_logic;
signal \N__20233\ : std_logic;
signal \N__20230\ : std_logic;
signal \N__20227\ : std_logic;
signal \N__20226\ : std_logic;
signal \N__20223\ : std_logic;
signal \N__20220\ : std_logic;
signal \N__20217\ : std_logic;
signal \N__20214\ : std_logic;
signal \N__20209\ : std_logic;
signal \N__20206\ : std_logic;
signal \N__20201\ : std_logic;
signal \N__20196\ : std_logic;
signal \N__20195\ : std_logic;
signal \N__20194\ : std_logic;
signal \N__20193\ : std_logic;
signal \N__20190\ : std_logic;
signal \N__20185\ : std_logic;
signal \N__20182\ : std_logic;
signal \N__20181\ : std_logic;
signal \N__20180\ : std_logic;
signal \N__20179\ : std_logic;
signal \N__20172\ : std_logic;
signal \N__20167\ : std_logic;
signal \N__20164\ : std_logic;
signal \N__20163\ : std_logic;
signal \N__20162\ : std_logic;
signal \N__20161\ : std_logic;
signal \N__20156\ : std_logic;
signal \N__20153\ : std_logic;
signal \N__20150\ : std_logic;
signal \N__20147\ : std_logic;
signal \N__20144\ : std_logic;
signal \N__20141\ : std_logic;
signal \N__20138\ : std_logic;
signal \N__20135\ : std_logic;
signal \N__20130\ : std_logic;
signal \N__20129\ : std_logic;
signal \N__20128\ : std_logic;
signal \N__20127\ : std_logic;
signal \N__20122\ : std_logic;
signal \N__20119\ : std_logic;
signal \N__20112\ : std_logic;
signal \N__20109\ : std_logic;
signal \N__20104\ : std_logic;
signal \N__20091\ : std_logic;
signal \N__20084\ : std_logic;
signal \N__20069\ : std_logic;
signal \N__20068\ : std_logic;
signal \N__20067\ : std_logic;
signal \N__20066\ : std_logic;
signal \N__20065\ : std_logic;
signal \N__20062\ : std_logic;
signal \N__20061\ : std_logic;
signal \N__20060\ : std_logic;
signal \N__20059\ : std_logic;
signal \N__20058\ : std_logic;
signal \N__20057\ : std_logic;
signal \N__20056\ : std_logic;
signal \N__20055\ : std_logic;
signal \N__20054\ : std_logic;
signal \N__20051\ : std_logic;
signal \N__20050\ : std_logic;
signal \N__20049\ : std_logic;
signal \N__20046\ : std_logic;
signal \N__20045\ : std_logic;
signal \N__20044\ : std_logic;
signal \N__20043\ : std_logic;
signal \N__20042\ : std_logic;
signal \N__20041\ : std_logic;
signal \N__20038\ : std_logic;
signal \N__20037\ : std_logic;
signal \N__20036\ : std_logic;
signal \N__20035\ : std_logic;
signal \N__20034\ : std_logic;
signal \N__20033\ : std_logic;
signal \N__20032\ : std_logic;
signal \N__20029\ : std_logic;
signal \N__20026\ : std_logic;
signal \N__20023\ : std_logic;
signal \N__20020\ : std_logic;
signal \N__20019\ : std_logic;
signal \N__20018\ : std_logic;
signal \N__20017\ : std_logic;
signal \N__20014\ : std_logic;
signal \N__20013\ : std_logic;
signal \N__20012\ : std_logic;
signal \N__20011\ : std_logic;
signal \N__20008\ : std_logic;
signal \N__20007\ : std_logic;
signal \N__20006\ : std_logic;
signal \N__20003\ : std_logic;
signal \N__20002\ : std_logic;
signal \N__20001\ : std_logic;
signal \N__19998\ : std_logic;
signal \N__19997\ : std_logic;
signal \N__19996\ : std_logic;
signal \N__19995\ : std_logic;
signal \N__19994\ : std_logic;
signal \N__19991\ : std_logic;
signal \N__19988\ : std_logic;
signal \N__19985\ : std_logic;
signal \N__19982\ : std_logic;
signal \N__19981\ : std_logic;
signal \N__19978\ : std_logic;
signal \N__19975\ : std_logic;
signal \N__19972\ : std_logic;
signal \N__19971\ : std_logic;
signal \N__19968\ : std_logic;
signal \N__19965\ : std_logic;
signal \N__19964\ : std_logic;
signal \N__19963\ : std_logic;
signal \N__19960\ : std_logic;
signal \N__19957\ : std_logic;
signal \N__19952\ : std_logic;
signal \N__19951\ : std_logic;
signal \N__19948\ : std_logic;
signal \N__19945\ : std_logic;
signal \N__19942\ : std_logic;
signal \N__19939\ : std_logic;
signal \N__19936\ : std_logic;
signal \N__19935\ : std_logic;
signal \N__19932\ : std_logic;
signal \N__19925\ : std_logic;
signal \N__19922\ : std_logic;
signal \N__19919\ : std_logic;
signal \N__19916\ : std_logic;
signal \N__19913\ : std_logic;
signal \N__19912\ : std_logic;
signal \N__19911\ : std_logic;
signal \N__19910\ : std_logic;
signal \N__19907\ : std_logic;
signal \N__19904\ : std_logic;
signal \N__19901\ : std_logic;
signal \N__19898\ : std_logic;
signal \N__19895\ : std_logic;
signal \N__19892\ : std_logic;
signal \N__19889\ : std_logic;
signal \N__19886\ : std_logic;
signal \N__19883\ : std_logic;
signal \N__19880\ : std_logic;
signal \N__19877\ : std_logic;
signal \N__19876\ : std_logic;
signal \N__19875\ : std_logic;
signal \N__19874\ : std_logic;
signal \N__19873\ : std_logic;
signal \N__19870\ : std_logic;
signal \N__19867\ : std_logic;
signal \N__19866\ : std_logic;
signal \N__19863\ : std_logic;
signal \N__19860\ : std_logic;
signal \N__19857\ : std_logic;
signal \N__19852\ : std_logic;
signal \N__19849\ : std_logic;
signal \N__19842\ : std_logic;
signal \N__19839\ : std_logic;
signal \N__19838\ : std_logic;
signal \N__19837\ : std_logic;
signal \N__19836\ : std_logic;
signal \N__19831\ : std_logic;
signal \N__19828\ : std_logic;
signal \N__19825\ : std_logic;
signal \N__19818\ : std_logic;
signal \N__19815\ : std_logic;
signal \N__19812\ : std_logic;
signal \N__19807\ : std_logic;
signal \N__19804\ : std_logic;
signal \N__19801\ : std_logic;
signal \N__19798\ : std_logic;
signal \N__19791\ : std_logic;
signal \N__19786\ : std_logic;
signal \N__19783\ : std_logic;
signal \N__19780\ : std_logic;
signal \N__19777\ : std_logic;
signal \N__19772\ : std_logic;
signal \N__19769\ : std_logic;
signal \N__19766\ : std_logic;
signal \N__19763\ : std_logic;
signal \N__19758\ : std_logic;
signal \N__19751\ : std_logic;
signal \N__19746\ : std_logic;
signal \N__19743\ : std_logic;
signal \N__19740\ : std_logic;
signal \N__19739\ : std_logic;
signal \N__19734\ : std_logic;
signal \N__19731\ : std_logic;
signal \N__19728\ : std_logic;
signal \N__19727\ : std_logic;
signal \N__19724\ : std_logic;
signal \N__19723\ : std_logic;
signal \N__19722\ : std_logic;
signal \N__19721\ : std_logic;
signal \N__19718\ : std_logic;
signal \N__19709\ : std_logic;
signal \N__19704\ : std_logic;
signal \N__19701\ : std_logic;
signal \N__19698\ : std_logic;
signal \N__19695\ : std_logic;
signal \N__19694\ : std_logic;
signal \N__19693\ : std_logic;
signal \N__19692\ : std_logic;
signal \N__19685\ : std_logic;
signal \N__19682\ : std_logic;
signal \N__19679\ : std_logic;
signal \N__19674\ : std_logic;
signal \N__19671\ : std_logic;
signal \N__19660\ : std_logic;
signal \N__19653\ : std_logic;
signal \N__19638\ : std_logic;
signal \N__19633\ : std_logic;
signal \N__19630\ : std_logic;
signal \N__19627\ : std_logic;
signal \N__19624\ : std_logic;
signal \N__19621\ : std_logic;
signal \N__19616\ : std_logic;
signal \N__19613\ : std_logic;
signal \N__19612\ : std_logic;
signal \N__19609\ : std_logic;
signal \N__19608\ : std_logic;
signal \N__19607\ : std_logic;
signal \N__19604\ : std_logic;
signal \N__19599\ : std_logic;
signal \N__19596\ : std_logic;
signal \N__19593\ : std_logic;
signal \N__19586\ : std_logic;
signal \N__19583\ : std_logic;
signal \N__19568\ : std_logic;
signal \N__19561\ : std_logic;
signal \N__19552\ : std_logic;
signal \N__19547\ : std_logic;
signal \N__19540\ : std_logic;
signal \N__19517\ : std_logic;
signal \N__19516\ : std_logic;
signal \N__19513\ : std_logic;
signal \N__19510\ : std_logic;
signal \N__19507\ : std_logic;
signal \N__19504\ : std_logic;
signal \N__19499\ : std_logic;
signal \N__19496\ : std_logic;
signal \N__19495\ : std_logic;
signal \N__19492\ : std_logic;
signal \N__19489\ : std_logic;
signal \N__19486\ : std_logic;
signal \N__19481\ : std_logic;
signal \N__19480\ : std_logic;
signal \N__19477\ : std_logic;
signal \N__19474\ : std_logic;
signal \N__19471\ : std_logic;
signal \N__19468\ : std_logic;
signal \N__19465\ : std_logic;
signal \N__19462\ : std_logic;
signal \N__19459\ : std_logic;
signal \N__19456\ : std_logic;
signal \N__19453\ : std_logic;
signal \N__19450\ : std_logic;
signal \N__19447\ : std_logic;
signal \N__19444\ : std_logic;
signal \N__19441\ : std_logic;
signal \N__19438\ : std_logic;
signal \N__19435\ : std_logic;
signal \N__19432\ : std_logic;
signal \N__19429\ : std_logic;
signal \N__19426\ : std_logic;
signal \N__19423\ : std_logic;
signal \N__19420\ : std_logic;
signal \N__19417\ : std_logic;
signal \N__19414\ : std_logic;
signal \N__19411\ : std_logic;
signal \N__19408\ : std_logic;
signal \N__19405\ : std_logic;
signal \N__19402\ : std_logic;
signal \N__19399\ : std_logic;
signal \N__19396\ : std_logic;
signal \N__19393\ : std_logic;
signal \N__19390\ : std_logic;
signal \N__19387\ : std_logic;
signal \N__19384\ : std_logic;
signal \N__19381\ : std_logic;
signal \N__19378\ : std_logic;
signal \N__19375\ : std_logic;
signal \N__19372\ : std_logic;
signal \N__19369\ : std_logic;
signal \N__19366\ : std_logic;
signal \N__19363\ : std_logic;
signal \N__19360\ : std_logic;
signal \N__19357\ : std_logic;
signal \N__19354\ : std_logic;
signal \N__19351\ : std_logic;
signal \N__19348\ : std_logic;
signal \N__19345\ : std_logic;
signal \N__19342\ : std_logic;
signal \N__19339\ : std_logic;
signal \N__19336\ : std_logic;
signal \N__19333\ : std_logic;
signal \N__19330\ : std_logic;
signal \N__19327\ : std_logic;
signal \N__19324\ : std_logic;
signal \N__19321\ : std_logic;
signal \N__19318\ : std_logic;
signal \N__19315\ : std_logic;
signal \N__19312\ : std_logic;
signal \N__19309\ : std_logic;
signal \N__19306\ : std_logic;
signal \N__19303\ : std_logic;
signal \N__19300\ : std_logic;
signal \N__19297\ : std_logic;
signal \N__19294\ : std_logic;
signal \N__19291\ : std_logic;
signal \N__19288\ : std_logic;
signal \N__19285\ : std_logic;
signal \N__19282\ : std_logic;
signal \N__19279\ : std_logic;
signal \N__19276\ : std_logic;
signal \N__19271\ : std_logic;
signal \N__19268\ : std_logic;
signal \N__19265\ : std_logic;
signal \N__19264\ : std_logic;
signal \N__19263\ : std_logic;
signal \N__19260\ : std_logic;
signal \N__19257\ : std_logic;
signal \N__19254\ : std_logic;
signal \N__19251\ : std_logic;
signal \N__19248\ : std_logic;
signal \N__19245\ : std_logic;
signal \N__19242\ : std_logic;
signal \N__19239\ : std_logic;
signal \N__19236\ : std_logic;
signal \N__19233\ : std_logic;
signal \N__19230\ : std_logic;
signal \N__19227\ : std_logic;
signal \N__19224\ : std_logic;
signal \N__19221\ : std_logic;
signal \N__19218\ : std_logic;
signal \N__19213\ : std_logic;
signal \N__19210\ : std_logic;
signal \N__19205\ : std_logic;
signal \N__19202\ : std_logic;
signal \N__19199\ : std_logic;
signal \N__19196\ : std_logic;
signal \N__19193\ : std_logic;
signal \N__19190\ : std_logic;
signal \N__19187\ : std_logic;
signal \N__19184\ : std_logic;
signal \N__19181\ : std_logic;
signal \N__19178\ : std_logic;
signal \N__19175\ : std_logic;
signal \N__19172\ : std_logic;
signal \N__19169\ : std_logic;
signal \N__19166\ : std_logic;
signal \N__19163\ : std_logic;
signal \N__19160\ : std_logic;
signal \N__19157\ : std_logic;
signal \N__19154\ : std_logic;
signal \N__19151\ : std_logic;
signal \N__19148\ : std_logic;
signal \N__19147\ : std_logic;
signal \N__19146\ : std_logic;
signal \N__19143\ : std_logic;
signal \N__19140\ : std_logic;
signal \N__19137\ : std_logic;
signal \N__19136\ : std_logic;
signal \N__19135\ : std_logic;
signal \N__19130\ : std_logic;
signal \N__19127\ : std_logic;
signal \N__19124\ : std_logic;
signal \N__19121\ : std_logic;
signal \N__19120\ : std_logic;
signal \N__19119\ : std_logic;
signal \N__19112\ : std_logic;
signal \N__19111\ : std_logic;
signal \N__19108\ : std_logic;
signal \N__19105\ : std_logic;
signal \N__19102\ : std_logic;
signal \N__19099\ : std_logic;
signal \N__19096\ : std_logic;
signal \N__19093\ : std_logic;
signal \N__19090\ : std_logic;
signal \N__19087\ : std_logic;
signal \N__19082\ : std_logic;
signal \N__19081\ : std_logic;
signal \N__19078\ : std_logic;
signal \N__19073\ : std_logic;
signal \N__19070\ : std_logic;
signal \N__19067\ : std_logic;
signal \N__19064\ : std_logic;
signal \N__19061\ : std_logic;
signal \N__19056\ : std_logic;
signal \N__19051\ : std_logic;
signal \N__19048\ : std_logic;
signal \N__19043\ : std_logic;
signal \N__19040\ : std_logic;
signal \N__19037\ : std_logic;
signal \N__19036\ : std_logic;
signal \N__19035\ : std_logic;
signal \N__19034\ : std_logic;
signal \N__19031\ : std_logic;
signal \N__19028\ : std_logic;
signal \N__19025\ : std_logic;
signal \N__19022\ : std_logic;
signal \N__19021\ : std_logic;
signal \N__19016\ : std_logic;
signal \N__19013\ : std_logic;
signal \N__19010\ : std_logic;
signal \N__19007\ : std_logic;
signal \N__19006\ : std_logic;
signal \N__19003\ : std_logic;
signal \N__19002\ : std_logic;
signal \N__19001\ : std_logic;
signal \N__18998\ : std_logic;
signal \N__18995\ : std_logic;
signal \N__18992\ : std_logic;
signal \N__18989\ : std_logic;
signal \N__18986\ : std_logic;
signal \N__18983\ : std_logic;
signal \N__18980\ : std_logic;
signal \N__18977\ : std_logic;
signal \N__18974\ : std_logic;
signal \N__18971\ : std_logic;
signal \N__18968\ : std_logic;
signal \N__18963\ : std_logic;
signal \N__18960\ : std_logic;
signal \N__18959\ : std_logic;
signal \N__18956\ : std_logic;
signal \N__18951\ : std_logic;
signal \N__18944\ : std_logic;
signal \N__18941\ : std_logic;
signal \N__18932\ : std_logic;
signal \N__18929\ : std_logic;
signal \N__18926\ : std_logic;
signal \N__18925\ : std_logic;
signal \N__18920\ : std_logic;
signal \N__18919\ : std_logic;
signal \N__18918\ : std_logic;
signal \N__18915\ : std_logic;
signal \N__18912\ : std_logic;
signal \N__18909\ : std_logic;
signal \N__18908\ : std_logic;
signal \N__18901\ : std_logic;
signal \N__18898\ : std_logic;
signal \N__18897\ : std_logic;
signal \N__18896\ : std_logic;
signal \N__18895\ : std_logic;
signal \N__18894\ : std_logic;
signal \N__18893\ : std_logic;
signal \N__18892\ : std_logic;
signal \N__18887\ : std_logic;
signal \N__18880\ : std_logic;
signal \N__18873\ : std_logic;
signal \N__18872\ : std_logic;
signal \N__18871\ : std_logic;
signal \N__18870\ : std_logic;
signal \N__18863\ : std_logic;
signal \N__18862\ : std_logic;
signal \N__18855\ : std_logic;
signal \N__18854\ : std_logic;
signal \N__18851\ : std_logic;
signal \N__18848\ : std_logic;
signal \N__18845\ : std_logic;
signal \N__18844\ : std_logic;
signal \N__18843\ : std_logic;
signal \N__18840\ : std_logic;
signal \N__18835\ : std_logic;
signal \N__18832\ : std_logic;
signal \N__18827\ : std_logic;
signal \N__18818\ : std_logic;
signal \N__18815\ : std_logic;
signal \N__18812\ : std_logic;
signal \N__18809\ : std_logic;
signal \N__18806\ : std_logic;
signal \N__18805\ : std_logic;
signal \N__18802\ : std_logic;
signal \N__18799\ : std_logic;
signal \N__18798\ : std_logic;
signal \N__18793\ : std_logic;
signal \N__18790\ : std_logic;
signal \N__18785\ : std_logic;
signal \N__18784\ : std_logic;
signal \N__18781\ : std_logic;
signal \N__18778\ : std_logic;
signal \N__18777\ : std_logic;
signal \N__18772\ : std_logic;
signal \N__18769\ : std_logic;
signal \N__18768\ : std_logic;
signal \N__18767\ : std_logic;
signal \N__18766\ : std_logic;
signal \N__18763\ : std_logic;
signal \N__18760\ : std_logic;
signal \N__18757\ : std_logic;
signal \N__18756\ : std_logic;
signal \N__18755\ : std_logic;
signal \N__18754\ : std_logic;
signal \N__18753\ : std_logic;
signal \N__18750\ : std_logic;
signal \N__18747\ : std_logic;
signal \N__18744\ : std_logic;
signal \N__18741\ : std_logic;
signal \N__18738\ : std_logic;
signal \N__18737\ : std_logic;
signal \N__18734\ : std_logic;
signal \N__18733\ : std_logic;
signal \N__18730\ : std_logic;
signal \N__18727\ : std_logic;
signal \N__18724\ : std_logic;
signal \N__18721\ : std_logic;
signal \N__18718\ : std_logic;
signal \N__18713\ : std_logic;
signal \N__18710\ : std_logic;
signal \N__18697\ : std_logic;
signal \N__18694\ : std_logic;
signal \N__18691\ : std_logic;
signal \N__18686\ : std_logic;
signal \N__18683\ : std_logic;
signal \N__18682\ : std_logic;
signal \N__18681\ : std_logic;
signal \N__18680\ : std_logic;
signal \N__18675\ : std_logic;
signal \N__18670\ : std_logic;
signal \N__18669\ : std_logic;
signal \N__18666\ : std_logic;
signal \N__18665\ : std_logic;
signal \N__18664\ : std_logic;
signal \N__18663\ : std_logic;
signal \N__18662\ : std_logic;
signal \N__18661\ : std_logic;
signal \N__18660\ : std_logic;
signal \N__18659\ : std_logic;
signal \N__18654\ : std_logic;
signal \N__18651\ : std_logic;
signal \N__18648\ : std_logic;
signal \N__18645\ : std_logic;
signal \N__18642\ : std_logic;
signal \N__18635\ : std_logic;
signal \N__18632\ : std_logic;
signal \N__18627\ : std_logic;
signal \N__18624\ : std_logic;
signal \N__18621\ : std_logic;
signal \N__18602\ : std_logic;
signal \N__18599\ : std_logic;
signal \N__18596\ : std_logic;
signal \N__18593\ : std_logic;
signal \N__18592\ : std_logic;
signal \N__18591\ : std_logic;
signal \N__18588\ : std_logic;
signal \N__18585\ : std_logic;
signal \N__18582\ : std_logic;
signal \N__18581\ : std_logic;
signal \N__18580\ : std_logic;
signal \N__18579\ : std_logic;
signal \N__18572\ : std_logic;
signal \N__18569\ : std_logic;
signal \N__18566\ : std_logic;
signal \N__18563\ : std_logic;
signal \N__18558\ : std_logic;
signal \N__18557\ : std_logic;
signal \N__18556\ : std_logic;
signal \N__18553\ : std_logic;
signal \N__18550\ : std_logic;
signal \N__18547\ : std_logic;
signal \N__18544\ : std_logic;
signal \N__18541\ : std_logic;
signal \N__18538\ : std_logic;
signal \N__18535\ : std_logic;
signal \N__18532\ : std_logic;
signal \N__18529\ : std_logic;
signal \N__18526\ : std_logic;
signal \N__18525\ : std_logic;
signal \N__18520\ : std_logic;
signal \N__18517\ : std_logic;
signal \N__18512\ : std_logic;
signal \N__18509\ : std_logic;
signal \N__18500\ : std_logic;
signal \N__18497\ : std_logic;
signal \N__18494\ : std_logic;
signal \N__18491\ : std_logic;
signal \N__18488\ : std_logic;
signal \N__18485\ : std_logic;
signal \N__18482\ : std_logic;
signal \N__18479\ : std_logic;
signal \N__18476\ : std_logic;
signal \N__18473\ : std_logic;
signal \N__18470\ : std_logic;
signal \N__18467\ : std_logic;
signal \N__18464\ : std_logic;
signal \N__18461\ : std_logic;
signal \N__18458\ : std_logic;
signal \N__18455\ : std_logic;
signal \N__18452\ : std_logic;
signal \N__18449\ : std_logic;
signal \N__18446\ : std_logic;
signal \N__18443\ : std_logic;
signal \N__18440\ : std_logic;
signal \N__18437\ : std_logic;
signal \N__18434\ : std_logic;
signal \N__18431\ : std_logic;
signal \N__18428\ : std_logic;
signal \N__18427\ : std_logic;
signal \N__18424\ : std_logic;
signal \N__18421\ : std_logic;
signal \N__18416\ : std_logic;
signal \N__18415\ : std_logic;
signal \N__18412\ : std_logic;
signal \N__18409\ : std_logic;
signal \N__18404\ : std_logic;
signal \N__18401\ : std_logic;
signal \N__18400\ : std_logic;
signal \N__18397\ : std_logic;
signal \N__18394\ : std_logic;
signal \N__18389\ : std_logic;
signal \N__18386\ : std_logic;
signal \N__18385\ : std_logic;
signal \N__18382\ : std_logic;
signal \N__18379\ : std_logic;
signal \N__18374\ : std_logic;
signal \N__18371\ : std_logic;
signal \N__18370\ : std_logic;
signal \N__18367\ : std_logic;
signal \N__18364\ : std_logic;
signal \N__18359\ : std_logic;
signal \N__18356\ : std_logic;
signal \N__18355\ : std_logic;
signal \N__18352\ : std_logic;
signal \N__18349\ : std_logic;
signal \N__18344\ : std_logic;
signal \N__18341\ : std_logic;
signal \N__18338\ : std_logic;
signal \N__18337\ : std_logic;
signal \N__18334\ : std_logic;
signal \N__18331\ : std_logic;
signal \N__18326\ : std_logic;
signal \N__18325\ : std_logic;
signal \N__18322\ : std_logic;
signal \N__18319\ : std_logic;
signal \N__18316\ : std_logic;
signal \N__18313\ : std_logic;
signal \N__18310\ : std_logic;
signal \N__18307\ : std_logic;
signal \N__18302\ : std_logic;
signal \N__18299\ : std_logic;
signal \N__18296\ : std_logic;
signal \N__18293\ : std_logic;
signal \N__18290\ : std_logic;
signal \N__18287\ : std_logic;
signal \N__18284\ : std_logic;
signal \N__18281\ : std_logic;
signal \N__18280\ : std_logic;
signal \N__18277\ : std_logic;
signal \N__18274\ : std_logic;
signal \N__18271\ : std_logic;
signal \N__18268\ : std_logic;
signal \N__18265\ : std_logic;
signal \N__18262\ : std_logic;
signal \N__18259\ : std_logic;
signal \N__18256\ : std_logic;
signal \N__18253\ : std_logic;
signal \N__18250\ : std_logic;
signal \N__18247\ : std_logic;
signal \N__18244\ : std_logic;
signal \N__18241\ : std_logic;
signal \N__18238\ : std_logic;
signal \N__18235\ : std_logic;
signal \N__18232\ : std_logic;
signal \N__18229\ : std_logic;
signal \N__18226\ : std_logic;
signal \N__18223\ : std_logic;
signal \N__18220\ : std_logic;
signal \N__18217\ : std_logic;
signal \N__18214\ : std_logic;
signal \N__18211\ : std_logic;
signal \N__18208\ : std_logic;
signal \N__18205\ : std_logic;
signal \N__18202\ : std_logic;
signal \N__18199\ : std_logic;
signal \N__18196\ : std_logic;
signal \N__18193\ : std_logic;
signal \N__18190\ : std_logic;
signal \N__18187\ : std_logic;
signal \N__18184\ : std_logic;
signal \N__18181\ : std_logic;
signal \N__18178\ : std_logic;
signal \N__18175\ : std_logic;
signal \N__18172\ : std_logic;
signal \N__18169\ : std_logic;
signal \N__18166\ : std_logic;
signal \N__18163\ : std_logic;
signal \N__18160\ : std_logic;
signal \N__18157\ : std_logic;
signal \N__18154\ : std_logic;
signal \N__18151\ : std_logic;
signal \N__18148\ : std_logic;
signal \N__18145\ : std_logic;
signal \N__18142\ : std_logic;
signal \N__18139\ : std_logic;
signal \N__18136\ : std_logic;
signal \N__18133\ : std_logic;
signal \N__18130\ : std_logic;
signal \N__18127\ : std_logic;
signal \N__18124\ : std_logic;
signal \N__18121\ : std_logic;
signal \N__18118\ : std_logic;
signal \N__18115\ : std_logic;
signal \N__18112\ : std_logic;
signal \N__18109\ : std_logic;
signal \N__18106\ : std_logic;
signal \N__18103\ : std_logic;
signal \N__18100\ : std_logic;
signal \N__18099\ : std_logic;
signal \N__18096\ : std_logic;
signal \N__18093\ : std_logic;
signal \N__18090\ : std_logic;
signal \N__18087\ : std_logic;
signal \N__18084\ : std_logic;
signal \N__18081\ : std_logic;
signal \N__18080\ : std_logic;
signal \N__18077\ : std_logic;
signal \N__18074\ : std_logic;
signal \N__18071\ : std_logic;
signal \N__18068\ : std_logic;
signal \N__18063\ : std_logic;
signal \N__18056\ : std_logic;
signal \N__18053\ : std_logic;
signal \N__18050\ : std_logic;
signal \N__18047\ : std_logic;
signal \N__18044\ : std_logic;
signal \N__18043\ : std_logic;
signal \N__18040\ : std_logic;
signal \N__18037\ : std_logic;
signal \N__18034\ : std_logic;
signal \N__18031\ : std_logic;
signal \N__18028\ : std_logic;
signal \N__18025\ : std_logic;
signal \N__18022\ : std_logic;
signal \N__18019\ : std_logic;
signal \N__18016\ : std_logic;
signal \N__18013\ : std_logic;
signal \N__18010\ : std_logic;
signal \N__18007\ : std_logic;
signal \N__18004\ : std_logic;
signal \N__18001\ : std_logic;
signal \N__17998\ : std_logic;
signal \N__17995\ : std_logic;
signal \N__17992\ : std_logic;
signal \N__17989\ : std_logic;
signal \N__17986\ : std_logic;
signal \N__17983\ : std_logic;
signal \N__17980\ : std_logic;
signal \N__17977\ : std_logic;
signal \N__17974\ : std_logic;
signal \N__17971\ : std_logic;
signal \N__17968\ : std_logic;
signal \N__17965\ : std_logic;
signal \N__17962\ : std_logic;
signal \N__17959\ : std_logic;
signal \N__17956\ : std_logic;
signal \N__17953\ : std_logic;
signal \N__17950\ : std_logic;
signal \N__17947\ : std_logic;
signal \N__17944\ : std_logic;
signal \N__17941\ : std_logic;
signal \N__17938\ : std_logic;
signal \N__17935\ : std_logic;
signal \N__17932\ : std_logic;
signal \N__17929\ : std_logic;
signal \N__17926\ : std_logic;
signal \N__17923\ : std_logic;
signal \N__17920\ : std_logic;
signal \N__17917\ : std_logic;
signal \N__17914\ : std_logic;
signal \N__17911\ : std_logic;
signal \N__17908\ : std_logic;
signal \N__17905\ : std_logic;
signal \N__17902\ : std_logic;
signal \N__17899\ : std_logic;
signal \N__17896\ : std_logic;
signal \N__17893\ : std_logic;
signal \N__17890\ : std_logic;
signal \N__17887\ : std_logic;
signal \N__17884\ : std_logic;
signal \N__17881\ : std_logic;
signal \N__17878\ : std_logic;
signal \N__17875\ : std_logic;
signal \N__17872\ : std_logic;
signal \N__17869\ : std_logic;
signal \N__17866\ : std_logic;
signal \N__17863\ : std_logic;
signal \N__17862\ : std_logic;
signal \N__17859\ : std_logic;
signal \N__17856\ : std_logic;
signal \N__17853\ : std_logic;
signal \N__17850\ : std_logic;
signal \N__17847\ : std_logic;
signal \N__17846\ : std_logic;
signal \N__17843\ : std_logic;
signal \N__17840\ : std_logic;
signal \N__17837\ : std_logic;
signal \N__17834\ : std_logic;
signal \N__17827\ : std_logic;
signal \N__17822\ : std_logic;
signal \N__17819\ : std_logic;
signal \N__17816\ : std_logic;
signal \N__17813\ : std_logic;
signal \N__17810\ : std_logic;
signal \N__17807\ : std_logic;
signal \N__17806\ : std_logic;
signal \N__17803\ : std_logic;
signal \N__17800\ : std_logic;
signal \N__17797\ : std_logic;
signal \N__17794\ : std_logic;
signal \N__17791\ : std_logic;
signal \N__17788\ : std_logic;
signal \N__17785\ : std_logic;
signal \N__17782\ : std_logic;
signal \N__17779\ : std_logic;
signal \N__17776\ : std_logic;
signal \N__17773\ : std_logic;
signal \N__17770\ : std_logic;
signal \N__17767\ : std_logic;
signal \N__17764\ : std_logic;
signal \N__17761\ : std_logic;
signal \N__17758\ : std_logic;
signal \N__17755\ : std_logic;
signal \N__17752\ : std_logic;
signal \N__17749\ : std_logic;
signal \N__17746\ : std_logic;
signal \N__17743\ : std_logic;
signal \N__17740\ : std_logic;
signal \N__17737\ : std_logic;
signal \N__17734\ : std_logic;
signal \N__17731\ : std_logic;
signal \N__17728\ : std_logic;
signal \N__17725\ : std_logic;
signal \N__17722\ : std_logic;
signal \N__17719\ : std_logic;
signal \N__17716\ : std_logic;
signal \N__17713\ : std_logic;
signal \N__17710\ : std_logic;
signal \N__17707\ : std_logic;
signal \N__17704\ : std_logic;
signal \N__17701\ : std_logic;
signal \N__17698\ : std_logic;
signal \N__17695\ : std_logic;
signal \N__17692\ : std_logic;
signal \N__17689\ : std_logic;
signal \N__17686\ : std_logic;
signal \N__17683\ : std_logic;
signal \N__17680\ : std_logic;
signal \N__17677\ : std_logic;
signal \N__17674\ : std_logic;
signal \N__17671\ : std_logic;
signal \N__17668\ : std_logic;
signal \N__17665\ : std_logic;
signal \N__17662\ : std_logic;
signal \N__17659\ : std_logic;
signal \N__17656\ : std_logic;
signal \N__17653\ : std_logic;
signal \N__17650\ : std_logic;
signal \N__17647\ : std_logic;
signal \N__17644\ : std_logic;
signal \N__17641\ : std_logic;
signal \N__17638\ : std_logic;
signal \N__17635\ : std_logic;
signal \N__17632\ : std_logic;
signal \N__17629\ : std_logic;
signal \N__17626\ : std_logic;
signal \N__17625\ : std_logic;
signal \N__17622\ : std_logic;
signal \N__17619\ : std_logic;
signal \N__17616\ : std_logic;
signal \N__17613\ : std_logic;
signal \N__17610\ : std_logic;
signal \N__17607\ : std_logic;
signal \N__17604\ : std_logic;
signal \N__17601\ : std_logic;
signal \N__17598\ : std_logic;
signal \N__17597\ : std_logic;
signal \N__17594\ : std_logic;
signal \N__17591\ : std_logic;
signal \N__17588\ : std_logic;
signal \N__17585\ : std_logic;
signal \N__17582\ : std_logic;
signal \N__17579\ : std_logic;
signal \N__17570\ : std_logic;
signal \N__17567\ : std_logic;
signal \N__17566\ : std_logic;
signal \N__17565\ : std_logic;
signal \N__17562\ : std_logic;
signal \N__17559\ : std_logic;
signal \N__17556\ : std_logic;
signal \N__17555\ : std_logic;
signal \N__17554\ : std_logic;
signal \N__17549\ : std_logic;
signal \N__17546\ : std_logic;
signal \N__17543\ : std_logic;
signal \N__17542\ : std_logic;
signal \N__17541\ : std_logic;
signal \N__17538\ : std_logic;
signal \N__17531\ : std_logic;
signal \N__17528\ : std_logic;
signal \N__17525\ : std_logic;
signal \N__17522\ : std_logic;
signal \N__17517\ : std_logic;
signal \N__17514\ : std_logic;
signal \N__17513\ : std_logic;
signal \N__17510\ : std_logic;
signal \N__17505\ : std_logic;
signal \N__17502\ : std_logic;
signal \N__17495\ : std_logic;
signal \N__17492\ : std_logic;
signal \N__17489\ : std_logic;
signal \N__17486\ : std_logic;
signal \N__17483\ : std_logic;
signal \N__17480\ : std_logic;
signal \N__17477\ : std_logic;
signal \N__17474\ : std_logic;
signal \N__17473\ : std_logic;
signal \N__17470\ : std_logic;
signal \N__17467\ : std_logic;
signal \N__17462\ : std_logic;
signal \N__17461\ : std_logic;
signal \N__17456\ : std_logic;
signal \N__17453\ : std_logic;
signal \N__17450\ : std_logic;
signal \N__17447\ : std_logic;
signal \N__17444\ : std_logic;
signal \N__17441\ : std_logic;
signal \N__17438\ : std_logic;
signal \N__17437\ : std_logic;
signal \N__17434\ : std_logic;
signal \N__17431\ : std_logic;
signal \N__17428\ : std_logic;
signal \N__17425\ : std_logic;
signal \N__17422\ : std_logic;
signal \N__17419\ : std_logic;
signal \N__17416\ : std_logic;
signal \N__17413\ : std_logic;
signal \N__17410\ : std_logic;
signal \N__17407\ : std_logic;
signal \N__17404\ : std_logic;
signal \N__17401\ : std_logic;
signal \N__17398\ : std_logic;
signal \N__17395\ : std_logic;
signal \N__17392\ : std_logic;
signal \N__17389\ : std_logic;
signal \N__17386\ : std_logic;
signal \N__17383\ : std_logic;
signal \N__17380\ : std_logic;
signal \N__17377\ : std_logic;
signal \N__17374\ : std_logic;
signal \N__17371\ : std_logic;
signal \N__17368\ : std_logic;
signal \N__17365\ : std_logic;
signal \N__17362\ : std_logic;
signal \N__17359\ : std_logic;
signal \N__17356\ : std_logic;
signal \N__17353\ : std_logic;
signal \N__17350\ : std_logic;
signal \N__17347\ : std_logic;
signal \N__17344\ : std_logic;
signal \N__17341\ : std_logic;
signal \N__17338\ : std_logic;
signal \N__17335\ : std_logic;
signal \N__17332\ : std_logic;
signal \N__17329\ : std_logic;
signal \N__17326\ : std_logic;
signal \N__17323\ : std_logic;
signal \N__17320\ : std_logic;
signal \N__17317\ : std_logic;
signal \N__17314\ : std_logic;
signal \N__17311\ : std_logic;
signal \N__17308\ : std_logic;
signal \N__17305\ : std_logic;
signal \N__17302\ : std_logic;
signal \N__17299\ : std_logic;
signal \N__17296\ : std_logic;
signal \N__17293\ : std_logic;
signal \N__17290\ : std_logic;
signal \N__17287\ : std_logic;
signal \N__17284\ : std_logic;
signal \N__17281\ : std_logic;
signal \N__17278\ : std_logic;
signal \N__17275\ : std_logic;
signal \N__17272\ : std_logic;
signal \N__17269\ : std_logic;
signal \N__17266\ : std_logic;
signal \N__17263\ : std_logic;
signal \N__17260\ : std_logic;
signal \N__17257\ : std_logic;
signal \N__17254\ : std_logic;
signal \N__17251\ : std_logic;
signal \N__17248\ : std_logic;
signal \N__17245\ : std_logic;
signal \N__17244\ : std_logic;
signal \N__17241\ : std_logic;
signal \N__17238\ : std_logic;
signal \N__17235\ : std_logic;
signal \N__17232\ : std_logic;
signal \N__17229\ : std_logic;
signal \N__17226\ : std_logic;
signal \N__17223\ : std_logic;
signal \N__17220\ : std_logic;
signal \N__17219\ : std_logic;
signal \N__17216\ : std_logic;
signal \N__17213\ : std_logic;
signal \N__17210\ : std_logic;
signal \N__17207\ : std_logic;
signal \N__17204\ : std_logic;
signal \N__17201\ : std_logic;
signal \N__17198\ : std_logic;
signal \N__17189\ : std_logic;
signal \N__17186\ : std_logic;
signal \N__17183\ : std_logic;
signal \N__17180\ : std_logic;
signal \N__17177\ : std_logic;
signal \N__17176\ : std_logic;
signal \N__17173\ : std_logic;
signal \N__17170\ : std_logic;
signal \N__17167\ : std_logic;
signal \N__17164\ : std_logic;
signal \N__17161\ : std_logic;
signal \N__17158\ : std_logic;
signal \N__17155\ : std_logic;
signal \N__17152\ : std_logic;
signal \N__17149\ : std_logic;
signal \N__17146\ : std_logic;
signal \N__17143\ : std_logic;
signal \N__17140\ : std_logic;
signal \N__17137\ : std_logic;
signal \N__17134\ : std_logic;
signal \N__17131\ : std_logic;
signal \N__17128\ : std_logic;
signal \N__17125\ : std_logic;
signal \N__17122\ : std_logic;
signal \N__17119\ : std_logic;
signal \N__17116\ : std_logic;
signal \N__17113\ : std_logic;
signal \N__17110\ : std_logic;
signal \N__17107\ : std_logic;
signal \N__17104\ : std_logic;
signal \N__17101\ : std_logic;
signal \N__17098\ : std_logic;
signal \N__17095\ : std_logic;
signal \N__17092\ : std_logic;
signal \N__17089\ : std_logic;
signal \N__17086\ : std_logic;
signal \N__17083\ : std_logic;
signal \N__17080\ : std_logic;
signal \N__17077\ : std_logic;
signal \N__17074\ : std_logic;
signal \N__17071\ : std_logic;
signal \N__17068\ : std_logic;
signal \N__17065\ : std_logic;
signal \N__17062\ : std_logic;
signal \N__17059\ : std_logic;
signal \N__17056\ : std_logic;
signal \N__17053\ : std_logic;
signal \N__17050\ : std_logic;
signal \N__17047\ : std_logic;
signal \N__17044\ : std_logic;
signal \N__17041\ : std_logic;
signal \N__17038\ : std_logic;
signal \N__17035\ : std_logic;
signal \N__17032\ : std_logic;
signal \N__17029\ : std_logic;
signal \N__17026\ : std_logic;
signal \N__17023\ : std_logic;
signal \N__17020\ : std_logic;
signal \N__17017\ : std_logic;
signal \N__17014\ : std_logic;
signal \N__17011\ : std_logic;
signal \N__17008\ : std_logic;
signal \N__17005\ : std_logic;
signal \N__17002\ : std_logic;
signal \N__16999\ : std_logic;
signal \N__16996\ : std_logic;
signal \N__16993\ : std_logic;
signal \N__16992\ : std_logic;
signal \N__16989\ : std_logic;
signal \N__16986\ : std_logic;
signal \N__16983\ : std_logic;
signal \N__16980\ : std_logic;
signal \N__16977\ : std_logic;
signal \N__16976\ : std_logic;
signal \N__16973\ : std_logic;
signal \N__16970\ : std_logic;
signal \N__16967\ : std_logic;
signal \N__16964\ : std_logic;
signal \N__16961\ : std_logic;
signal \N__16958\ : std_logic;
signal \N__16955\ : std_logic;
signal \N__16952\ : std_logic;
signal \N__16949\ : std_logic;
signal \N__16946\ : std_logic;
signal \N__16943\ : std_logic;
signal \N__16934\ : std_logic;
signal \N__16931\ : std_logic;
signal \N__16928\ : std_logic;
signal \N__16925\ : std_logic;
signal \N__16922\ : std_logic;
signal \N__16919\ : std_logic;
signal \N__16918\ : std_logic;
signal \N__16915\ : std_logic;
signal \N__16912\ : std_logic;
signal \N__16909\ : std_logic;
signal \N__16906\ : std_logic;
signal \N__16903\ : std_logic;
signal \N__16900\ : std_logic;
signal \N__16897\ : std_logic;
signal \N__16894\ : std_logic;
signal \N__16891\ : std_logic;
signal \N__16888\ : std_logic;
signal \N__16885\ : std_logic;
signal \N__16882\ : std_logic;
signal \N__16879\ : std_logic;
signal \N__16876\ : std_logic;
signal \N__16873\ : std_logic;
signal \N__16870\ : std_logic;
signal \N__16867\ : std_logic;
signal \N__16864\ : std_logic;
signal \N__16861\ : std_logic;
signal \N__16858\ : std_logic;
signal \N__16855\ : std_logic;
signal \N__16852\ : std_logic;
signal \N__16849\ : std_logic;
signal \N__16846\ : std_logic;
signal \N__16843\ : std_logic;
signal \N__16840\ : std_logic;
signal \N__16837\ : std_logic;
signal \N__16834\ : std_logic;
signal \N__16831\ : std_logic;
signal \N__16828\ : std_logic;
signal \N__16825\ : std_logic;
signal \N__16822\ : std_logic;
signal \N__16819\ : std_logic;
signal \N__16816\ : std_logic;
signal \N__16813\ : std_logic;
signal \N__16810\ : std_logic;
signal \N__16807\ : std_logic;
signal \N__16804\ : std_logic;
signal \N__16801\ : std_logic;
signal \N__16798\ : std_logic;
signal \N__16795\ : std_logic;
signal \N__16792\ : std_logic;
signal \N__16789\ : std_logic;
signal \N__16786\ : std_logic;
signal \N__16783\ : std_logic;
signal \N__16780\ : std_logic;
signal \N__16777\ : std_logic;
signal \N__16774\ : std_logic;
signal \N__16771\ : std_logic;
signal \N__16768\ : std_logic;
signal \N__16765\ : std_logic;
signal \N__16762\ : std_logic;
signal \N__16759\ : std_logic;
signal \N__16756\ : std_logic;
signal \N__16753\ : std_logic;
signal \N__16750\ : std_logic;
signal \N__16747\ : std_logic;
signal \N__16744\ : std_logic;
signal \N__16741\ : std_logic;
signal \N__16738\ : std_logic;
signal \N__16735\ : std_logic;
signal \N__16732\ : std_logic;
signal \N__16729\ : std_logic;
signal \N__16726\ : std_logic;
signal \N__16725\ : std_logic;
signal \N__16722\ : std_logic;
signal \N__16719\ : std_logic;
signal \N__16716\ : std_logic;
signal \N__16713\ : std_logic;
signal \N__16710\ : std_logic;
signal \N__16707\ : std_logic;
signal \N__16704\ : std_logic;
signal \N__16701\ : std_logic;
signal \N__16700\ : std_logic;
signal \N__16697\ : std_logic;
signal \N__16694\ : std_logic;
signal \N__16691\ : std_logic;
signal \N__16688\ : std_logic;
signal \N__16683\ : std_logic;
signal \N__16680\ : std_logic;
signal \N__16673\ : std_logic;
signal \N__16670\ : std_logic;
signal \N__16667\ : std_logic;
signal \N__16664\ : std_logic;
signal \N__16661\ : std_logic;
signal \N__16658\ : std_logic;
signal \N__16657\ : std_logic;
signal \N__16654\ : std_logic;
signal \N__16651\ : std_logic;
signal \N__16648\ : std_logic;
signal \N__16645\ : std_logic;
signal \N__16642\ : std_logic;
signal \N__16639\ : std_logic;
signal \N__16636\ : std_logic;
signal \N__16633\ : std_logic;
signal \N__16630\ : std_logic;
signal \N__16627\ : std_logic;
signal \N__16624\ : std_logic;
signal \N__16621\ : std_logic;
signal \N__16618\ : std_logic;
signal \N__16615\ : std_logic;
signal \N__16612\ : std_logic;
signal \N__16609\ : std_logic;
signal \N__16606\ : std_logic;
signal \N__16603\ : std_logic;
signal \N__16600\ : std_logic;
signal \N__16597\ : std_logic;
signal \N__16594\ : std_logic;
signal \N__16591\ : std_logic;
signal \N__16588\ : std_logic;
signal \N__16585\ : std_logic;
signal \N__16582\ : std_logic;
signal \N__16579\ : std_logic;
signal \N__16576\ : std_logic;
signal \N__16573\ : std_logic;
signal \N__16570\ : std_logic;
signal \N__16567\ : std_logic;
signal \N__16564\ : std_logic;
signal \N__16561\ : std_logic;
signal \N__16558\ : std_logic;
signal \N__16555\ : std_logic;
signal \N__16552\ : std_logic;
signal \N__16549\ : std_logic;
signal \N__16546\ : std_logic;
signal \N__16543\ : std_logic;
signal \N__16540\ : std_logic;
signal \N__16537\ : std_logic;
signal \N__16534\ : std_logic;
signal \N__16531\ : std_logic;
signal \N__16528\ : std_logic;
signal \N__16525\ : std_logic;
signal \N__16522\ : std_logic;
signal \N__16519\ : std_logic;
signal \N__16516\ : std_logic;
signal \N__16513\ : std_logic;
signal \N__16510\ : std_logic;
signal \N__16507\ : std_logic;
signal \N__16504\ : std_logic;
signal \N__16501\ : std_logic;
signal \N__16498\ : std_logic;
signal \N__16495\ : std_logic;
signal \N__16492\ : std_logic;
signal \N__16489\ : std_logic;
signal \N__16486\ : std_logic;
signal \N__16483\ : std_logic;
signal \N__16480\ : std_logic;
signal \N__16477\ : std_logic;
signal \N__16474\ : std_logic;
signal \N__16471\ : std_logic;
signal \N__16468\ : std_logic;
signal \N__16465\ : std_logic;
signal \N__16464\ : std_logic;
signal \N__16461\ : std_logic;
signal \N__16458\ : std_logic;
signal \N__16457\ : std_logic;
signal \N__16454\ : std_logic;
signal \N__16451\ : std_logic;
signal \N__16448\ : std_logic;
signal \N__16445\ : std_logic;
signal \N__16442\ : std_logic;
signal \N__16439\ : std_logic;
signal \N__16436\ : std_logic;
signal \N__16433\ : std_logic;
signal \N__16430\ : std_logic;
signal \N__16425\ : std_logic;
signal \N__16418\ : std_logic;
signal \N__16415\ : std_logic;
signal \N__16412\ : std_logic;
signal \N__16409\ : std_logic;
signal \N__16406\ : std_logic;
signal \N__16405\ : std_logic;
signal \N__16404\ : std_logic;
signal \N__16401\ : std_logic;
signal \N__16398\ : std_logic;
signal \N__16397\ : std_logic;
signal \N__16394\ : std_logic;
signal \N__16391\ : std_logic;
signal \N__16388\ : std_logic;
signal \N__16385\ : std_logic;
signal \N__16382\ : std_logic;
signal \N__16373\ : std_logic;
signal \N__16370\ : std_logic;
signal \N__16367\ : std_logic;
signal \N__16364\ : std_logic;
signal \N__16361\ : std_logic;
signal \N__16358\ : std_logic;
signal \N__16355\ : std_logic;
signal \N__16354\ : std_logic;
signal \N__16351\ : std_logic;
signal \N__16348\ : std_logic;
signal \N__16345\ : std_logic;
signal \N__16342\ : std_logic;
signal \N__16339\ : std_logic;
signal \N__16336\ : std_logic;
signal \N__16333\ : std_logic;
signal \N__16330\ : std_logic;
signal \N__16327\ : std_logic;
signal \N__16324\ : std_logic;
signal \N__16321\ : std_logic;
signal \N__16318\ : std_logic;
signal \N__16315\ : std_logic;
signal \N__16312\ : std_logic;
signal \N__16309\ : std_logic;
signal \N__16306\ : std_logic;
signal \N__16303\ : std_logic;
signal \N__16300\ : std_logic;
signal \N__16297\ : std_logic;
signal \N__16294\ : std_logic;
signal \N__16291\ : std_logic;
signal \N__16288\ : std_logic;
signal \N__16285\ : std_logic;
signal \N__16282\ : std_logic;
signal \N__16279\ : std_logic;
signal \N__16276\ : std_logic;
signal \N__16273\ : std_logic;
signal \N__16270\ : std_logic;
signal \N__16267\ : std_logic;
signal \N__16264\ : std_logic;
signal \N__16261\ : std_logic;
signal \N__16258\ : std_logic;
signal \N__16255\ : std_logic;
signal \N__16252\ : std_logic;
signal \N__16249\ : std_logic;
signal \N__16246\ : std_logic;
signal \N__16243\ : std_logic;
signal \N__16240\ : std_logic;
signal \N__16237\ : std_logic;
signal \N__16234\ : std_logic;
signal \N__16231\ : std_logic;
signal \N__16228\ : std_logic;
signal \N__16225\ : std_logic;
signal \N__16222\ : std_logic;
signal \N__16219\ : std_logic;
signal \N__16216\ : std_logic;
signal \N__16213\ : std_logic;
signal \N__16210\ : std_logic;
signal \N__16207\ : std_logic;
signal \N__16204\ : std_logic;
signal \N__16201\ : std_logic;
signal \N__16198\ : std_logic;
signal \N__16195\ : std_logic;
signal \N__16192\ : std_logic;
signal \N__16189\ : std_logic;
signal \N__16186\ : std_logic;
signal \N__16183\ : std_logic;
signal \N__16180\ : std_logic;
signal \N__16177\ : std_logic;
signal \N__16174\ : std_logic;
signal \N__16173\ : std_logic;
signal \N__16170\ : std_logic;
signal \N__16167\ : std_logic;
signal \N__16164\ : std_logic;
signal \N__16161\ : std_logic;
signal \N__16158\ : std_logic;
signal \N__16155\ : std_logic;
signal \N__16152\ : std_logic;
signal \N__16149\ : std_logic;
signal \N__16146\ : std_logic;
signal \N__16145\ : std_logic;
signal \N__16142\ : std_logic;
signal \N__16139\ : std_logic;
signal \N__16136\ : std_logic;
signal \N__16133\ : std_logic;
signal \N__16128\ : std_logic;
signal \N__16121\ : std_logic;
signal \N__16120\ : std_logic;
signal \N__16117\ : std_logic;
signal \N__16114\ : std_logic;
signal \N__16111\ : std_logic;
signal \N__16108\ : std_logic;
signal \N__16105\ : std_logic;
signal \N__16102\ : std_logic;
signal \N__16099\ : std_logic;
signal \N__16096\ : std_logic;
signal \N__16093\ : std_logic;
signal \N__16090\ : std_logic;
signal \N__16085\ : std_logic;
signal \N__16084\ : std_logic;
signal \N__16081\ : std_logic;
signal \N__16078\ : std_logic;
signal \N__16075\ : std_logic;
signal \N__16074\ : std_logic;
signal \N__16071\ : std_logic;
signal \N__16068\ : std_logic;
signal \N__16065\ : std_logic;
signal \N__16062\ : std_logic;
signal \N__16057\ : std_logic;
signal \N__16054\ : std_logic;
signal \N__16051\ : std_logic;
signal \N__16048\ : std_logic;
signal \N__16045\ : std_logic;
signal \N__16042\ : std_logic;
signal \N__16039\ : std_logic;
signal \N__16034\ : std_logic;
signal \N__16031\ : std_logic;
signal \N__16028\ : std_logic;
signal \N__16025\ : std_logic;
signal \N__16022\ : std_logic;
signal \N__16021\ : std_logic;
signal \N__16018\ : std_logic;
signal \N__16015\ : std_logic;
signal \N__16012\ : std_logic;
signal \N__16009\ : std_logic;
signal \N__16006\ : std_logic;
signal \N__16003\ : std_logic;
signal \N__16000\ : std_logic;
signal \N__15997\ : std_logic;
signal \N__15994\ : std_logic;
signal \N__15991\ : std_logic;
signal \N__15988\ : std_logic;
signal \N__15985\ : std_logic;
signal \N__15982\ : std_logic;
signal \N__15979\ : std_logic;
signal \N__15976\ : std_logic;
signal \N__15973\ : std_logic;
signal \N__15970\ : std_logic;
signal \N__15967\ : std_logic;
signal \N__15964\ : std_logic;
signal \N__15961\ : std_logic;
signal \N__15958\ : std_logic;
signal \N__15955\ : std_logic;
signal \N__15952\ : std_logic;
signal \N__15949\ : std_logic;
signal \N__15946\ : std_logic;
signal \N__15943\ : std_logic;
signal \N__15940\ : std_logic;
signal \N__15937\ : std_logic;
signal \N__15934\ : std_logic;
signal \N__15931\ : std_logic;
signal \N__15928\ : std_logic;
signal \N__15925\ : std_logic;
signal \N__15922\ : std_logic;
signal \N__15919\ : std_logic;
signal \N__15916\ : std_logic;
signal \N__15913\ : std_logic;
signal \N__15910\ : std_logic;
signal \N__15907\ : std_logic;
signal \N__15904\ : std_logic;
signal \N__15901\ : std_logic;
signal \N__15898\ : std_logic;
signal \N__15895\ : std_logic;
signal \N__15892\ : std_logic;
signal \N__15889\ : std_logic;
signal \N__15886\ : std_logic;
signal \N__15883\ : std_logic;
signal \N__15880\ : std_logic;
signal \N__15877\ : std_logic;
signal \N__15874\ : std_logic;
signal \N__15871\ : std_logic;
signal \N__15868\ : std_logic;
signal \N__15865\ : std_logic;
signal \N__15862\ : std_logic;
signal \N__15859\ : std_logic;
signal \N__15856\ : std_logic;
signal \N__15853\ : std_logic;
signal \N__15850\ : std_logic;
signal \N__15847\ : std_logic;
signal \N__15844\ : std_logic;
signal \N__15841\ : std_logic;
signal \N__15838\ : std_logic;
signal \N__15835\ : std_logic;
signal \N__15832\ : std_logic;
signal \N__15829\ : std_logic;
signal \N__15828\ : std_logic;
signal \N__15825\ : std_logic;
signal \N__15822\ : std_logic;
signal \N__15819\ : std_logic;
signal \N__15816\ : std_logic;
signal \N__15813\ : std_logic;
signal \N__15812\ : std_logic;
signal \N__15809\ : std_logic;
signal \N__15806\ : std_logic;
signal \N__15803\ : std_logic;
signal \N__15800\ : std_logic;
signal \N__15795\ : std_logic;
signal \N__15792\ : std_logic;
signal \N__15785\ : std_logic;
signal \N__15782\ : std_logic;
signal \N__15779\ : std_logic;
signal \N__15776\ : std_logic;
signal \N__15773\ : std_logic;
signal \N__15770\ : std_logic;
signal \N__15767\ : std_logic;
signal \N__15764\ : std_logic;
signal \N__15761\ : std_logic;
signal \N__15758\ : std_logic;
signal \N__15755\ : std_logic;
signal \N__15752\ : std_logic;
signal \N__15749\ : std_logic;
signal \N__15746\ : std_logic;
signal \N__15743\ : std_logic;
signal \N__15740\ : std_logic;
signal \N__15737\ : std_logic;
signal \N__15734\ : std_logic;
signal \N__15733\ : std_logic;
signal \N__15730\ : std_logic;
signal \N__15727\ : std_logic;
signal \N__15724\ : std_logic;
signal \N__15721\ : std_logic;
signal \N__15718\ : std_logic;
signal \N__15715\ : std_logic;
signal \N__15712\ : std_logic;
signal \N__15709\ : std_logic;
signal \N__15706\ : std_logic;
signal \N__15703\ : std_logic;
signal \N__15700\ : std_logic;
signal \N__15697\ : std_logic;
signal \N__15694\ : std_logic;
signal \N__15691\ : std_logic;
signal \N__15688\ : std_logic;
signal \N__15685\ : std_logic;
signal \N__15682\ : std_logic;
signal \N__15679\ : std_logic;
signal \N__15676\ : std_logic;
signal \N__15673\ : std_logic;
signal \N__15670\ : std_logic;
signal \N__15667\ : std_logic;
signal \N__15664\ : std_logic;
signal \N__15661\ : std_logic;
signal \N__15658\ : std_logic;
signal \N__15655\ : std_logic;
signal \N__15652\ : std_logic;
signal \N__15649\ : std_logic;
signal \N__15646\ : std_logic;
signal \N__15643\ : std_logic;
signal \N__15640\ : std_logic;
signal \N__15637\ : std_logic;
signal \N__15634\ : std_logic;
signal \N__15631\ : std_logic;
signal \N__15628\ : std_logic;
signal \N__15625\ : std_logic;
signal \N__15622\ : std_logic;
signal \N__15619\ : std_logic;
signal \N__15616\ : std_logic;
signal \N__15613\ : std_logic;
signal \N__15610\ : std_logic;
signal \N__15607\ : std_logic;
signal \N__15604\ : std_logic;
signal \N__15601\ : std_logic;
signal \N__15598\ : std_logic;
signal \N__15595\ : std_logic;
signal \N__15592\ : std_logic;
signal \N__15589\ : std_logic;
signal \N__15586\ : std_logic;
signal \N__15583\ : std_logic;
signal \N__15580\ : std_logic;
signal \N__15577\ : std_logic;
signal \N__15574\ : std_logic;
signal \N__15571\ : std_logic;
signal \N__15568\ : std_logic;
signal \N__15565\ : std_logic;
signal \N__15562\ : std_logic;
signal \N__15559\ : std_logic;
signal \N__15556\ : std_logic;
signal \N__15553\ : std_logic;
signal \N__15550\ : std_logic;
signal \N__15547\ : std_logic;
signal \N__15544\ : std_logic;
signal \N__15541\ : std_logic;
signal \N__15540\ : std_logic;
signal \N__15537\ : std_logic;
signal \N__15534\ : std_logic;
signal \N__15531\ : std_logic;
signal \N__15528\ : std_logic;
signal \N__15525\ : std_logic;
signal \N__15522\ : std_logic;
signal \N__15519\ : std_logic;
signal \N__15516\ : std_logic;
signal \N__15515\ : std_logic;
signal \N__15512\ : std_logic;
signal \N__15509\ : std_logic;
signal \N__15506\ : std_logic;
signal \N__15503\ : std_logic;
signal \N__15496\ : std_logic;
signal \N__15491\ : std_logic;
signal \N__15488\ : std_logic;
signal \N__15485\ : std_logic;
signal \N__15482\ : std_logic;
signal \N__15481\ : std_logic;
signal \N__15478\ : std_logic;
signal \N__15475\ : std_logic;
signal \N__15472\ : std_logic;
signal \N__15469\ : std_logic;
signal \N__15466\ : std_logic;
signal \N__15463\ : std_logic;
signal \N__15460\ : std_logic;
signal \N__15457\ : std_logic;
signal \N__15454\ : std_logic;
signal \N__15451\ : std_logic;
signal \N__15448\ : std_logic;
signal \N__15445\ : std_logic;
signal \N__15442\ : std_logic;
signal \N__15439\ : std_logic;
signal \N__15436\ : std_logic;
signal \N__15433\ : std_logic;
signal \N__15430\ : std_logic;
signal \N__15427\ : std_logic;
signal \N__15424\ : std_logic;
signal \N__15421\ : std_logic;
signal \N__15418\ : std_logic;
signal \N__15415\ : std_logic;
signal \N__15412\ : std_logic;
signal \N__15409\ : std_logic;
signal \N__15406\ : std_logic;
signal \N__15403\ : std_logic;
signal \N__15400\ : std_logic;
signal \N__15397\ : std_logic;
signal \N__15394\ : std_logic;
signal \N__15391\ : std_logic;
signal \N__15388\ : std_logic;
signal \N__15385\ : std_logic;
signal \N__15382\ : std_logic;
signal \N__15379\ : std_logic;
signal \N__15376\ : std_logic;
signal \N__15373\ : std_logic;
signal \N__15370\ : std_logic;
signal \N__15367\ : std_logic;
signal \N__15364\ : std_logic;
signal \N__15361\ : std_logic;
signal \N__15358\ : std_logic;
signal \N__15355\ : std_logic;
signal \N__15352\ : std_logic;
signal \N__15349\ : std_logic;
signal \N__15346\ : std_logic;
signal \N__15343\ : std_logic;
signal \N__15340\ : std_logic;
signal \N__15337\ : std_logic;
signal \N__15334\ : std_logic;
signal \N__15331\ : std_logic;
signal \N__15328\ : std_logic;
signal \N__15325\ : std_logic;
signal \N__15322\ : std_logic;
signal \N__15319\ : std_logic;
signal \N__15316\ : std_logic;
signal \N__15313\ : std_logic;
signal \N__15310\ : std_logic;
signal \N__15307\ : std_logic;
signal \N__15304\ : std_logic;
signal \N__15301\ : std_logic;
signal \N__15298\ : std_logic;
signal \N__15295\ : std_logic;
signal \N__15292\ : std_logic;
signal \N__15289\ : std_logic;
signal \N__15288\ : std_logic;
signal \N__15285\ : std_logic;
signal \N__15282\ : std_logic;
signal \N__15279\ : std_logic;
signal \N__15276\ : std_logic;
signal \N__15273\ : std_logic;
signal \N__15272\ : std_logic;
signal \N__15269\ : std_logic;
signal \N__15266\ : std_logic;
signal \N__15263\ : std_logic;
signal \N__15260\ : std_logic;
signal \N__15255\ : std_logic;
signal \N__15252\ : std_logic;
signal \N__15245\ : std_logic;
signal \N__15242\ : std_logic;
signal \N__15239\ : std_logic;
signal \N__15236\ : std_logic;
signal \N__15233\ : std_logic;
signal \N__15230\ : std_logic;
signal \N__15227\ : std_logic;
signal \N__15224\ : std_logic;
signal \N__15221\ : std_logic;
signal \N__15218\ : std_logic;
signal \N__15215\ : std_logic;
signal \N__15212\ : std_logic;
signal \N__15209\ : std_logic;
signal \N__15206\ : std_logic;
signal \N__15203\ : std_logic;
signal \N__15200\ : std_logic;
signal \N__15199\ : std_logic;
signal \N__15196\ : std_logic;
signal \N__15193\ : std_logic;
signal \N__15188\ : std_logic;
signal \N__15185\ : std_logic;
signal \N__15182\ : std_logic;
signal \N__15179\ : std_logic;
signal \N__15176\ : std_logic;
signal \N__15175\ : std_logic;
signal \N__15174\ : std_logic;
signal \N__15173\ : std_logic;
signal \N__15170\ : std_logic;
signal \N__15167\ : std_logic;
signal \N__15164\ : std_logic;
signal \N__15161\ : std_logic;
signal \N__15156\ : std_logic;
signal \N__15153\ : std_logic;
signal \N__15146\ : std_logic;
signal \N__15145\ : std_logic;
signal \N__15144\ : std_logic;
signal \N__15143\ : std_logic;
signal \N__15142\ : std_logic;
signal \N__15141\ : std_logic;
signal \N__15140\ : std_logic;
signal \N__15137\ : std_logic;
signal \N__15134\ : std_logic;
signal \N__15131\ : std_logic;
signal \N__15128\ : std_logic;
signal \N__15127\ : std_logic;
signal \N__15126\ : std_logic;
signal \N__15123\ : std_logic;
signal \N__15120\ : std_logic;
signal \N__15119\ : std_logic;
signal \N__15116\ : std_logic;
signal \N__15115\ : std_logic;
signal \N__15114\ : std_logic;
signal \N__15111\ : std_logic;
signal \N__15106\ : std_logic;
signal \N__15103\ : std_logic;
signal \N__15098\ : std_logic;
signal \N__15097\ : std_logic;
signal \N__15096\ : std_logic;
signal \N__15093\ : std_logic;
signal \N__15090\ : std_logic;
signal \N__15087\ : std_logic;
signal \N__15084\ : std_logic;
signal \N__15081\ : std_logic;
signal \N__15078\ : std_logic;
signal \N__15069\ : std_logic;
signal \N__15066\ : std_logic;
signal \N__15063\ : std_logic;
signal \N__15044\ : std_logic;
signal \N__15041\ : std_logic;
signal \N__15038\ : std_logic;
signal \N__15035\ : std_logic;
signal \N__15032\ : std_logic;
signal \N__15031\ : std_logic;
signal \N__15028\ : std_logic;
signal \N__15025\ : std_logic;
signal \N__15024\ : std_logic;
signal \N__15019\ : std_logic;
signal \N__15016\ : std_logic;
signal \N__15015\ : std_logic;
signal \N__15010\ : std_logic;
signal \N__15007\ : std_logic;
signal \N__15002\ : std_logic;
signal \N__14999\ : std_logic;
signal \N__14996\ : std_logic;
signal \N__14993\ : std_logic;
signal \N__14992\ : std_logic;
signal \N__14989\ : std_logic;
signal \N__14988\ : std_logic;
signal \N__14987\ : std_logic;
signal \N__14984\ : std_logic;
signal \N__14981\ : std_logic;
signal \N__14978\ : std_logic;
signal \N__14975\ : std_logic;
signal \N__14972\ : std_logic;
signal \N__14965\ : std_logic;
signal \N__14962\ : std_logic;
signal \N__14959\ : std_logic;
signal \N__14956\ : std_logic;
signal \N__14953\ : std_logic;
signal \N__14950\ : std_logic;
signal \N__14947\ : std_logic;
signal \N__14944\ : std_logic;
signal \N__14939\ : std_logic;
signal \N__14936\ : std_logic;
signal \N__14933\ : std_logic;
signal \N__14930\ : std_logic;
signal \N__14927\ : std_logic;
signal \N__14924\ : std_logic;
signal \N__14923\ : std_logic;
signal \N__14922\ : std_logic;
signal \N__14921\ : std_logic;
signal \N__14920\ : std_logic;
signal \N__14919\ : std_logic;
signal \N__14918\ : std_logic;
signal \N__14917\ : std_logic;
signal \N__14916\ : std_logic;
signal \N__14913\ : std_logic;
signal \N__14910\ : std_logic;
signal \N__14903\ : std_logic;
signal \N__14896\ : std_logic;
signal \N__14893\ : std_logic;
signal \N__14882\ : std_logic;
signal \N__14881\ : std_logic;
signal \N__14880\ : std_logic;
signal \N__14879\ : std_logic;
signal \N__14876\ : std_logic;
signal \N__14869\ : std_logic;
signal \N__14868\ : std_logic;
signal \N__14867\ : std_logic;
signal \N__14866\ : std_logic;
signal \N__14865\ : std_logic;
signal \N__14864\ : std_logic;
signal \N__14861\ : std_logic;
signal \N__14858\ : std_logic;
signal \N__14855\ : std_logic;
signal \N__14852\ : std_logic;
signal \N__14847\ : std_logic;
signal \N__14844\ : std_logic;
signal \N__14839\ : std_logic;
signal \N__14828\ : std_logic;
signal \N__14827\ : std_logic;
signal \N__14826\ : std_logic;
signal \N__14825\ : std_logic;
signal \N__14824\ : std_logic;
signal \N__14823\ : std_logic;
signal \N__14822\ : std_logic;
signal \N__14821\ : std_logic;
signal \N__14818\ : std_logic;
signal \N__14817\ : std_logic;
signal \N__14814\ : std_logic;
signal \N__14811\ : std_logic;
signal \N__14808\ : std_logic;
signal \N__14805\ : std_logic;
signal \N__14802\ : std_logic;
signal \N__14799\ : std_logic;
signal \N__14796\ : std_logic;
signal \N__14793\ : std_logic;
signal \N__14790\ : std_logic;
signal \N__14787\ : std_logic;
signal \N__14784\ : std_logic;
signal \N__14781\ : std_logic;
signal \N__14776\ : std_logic;
signal \N__14771\ : std_logic;
signal \N__14768\ : std_logic;
signal \N__14753\ : std_logic;
signal \N__14750\ : std_logic;
signal \N__14749\ : std_logic;
signal \N__14748\ : std_logic;
signal \N__14745\ : std_logic;
signal \N__14742\ : std_logic;
signal \N__14741\ : std_logic;
signal \N__14738\ : std_logic;
signal \N__14735\ : std_logic;
signal \N__14732\ : std_logic;
signal \N__14729\ : std_logic;
signal \N__14726\ : std_logic;
signal \N__14723\ : std_logic;
signal \N__14720\ : std_logic;
signal \N__14717\ : std_logic;
signal \N__14714\ : std_logic;
signal \N__14711\ : std_logic;
signal \N__14706\ : std_logic;
signal \N__14703\ : std_logic;
signal \N__14698\ : std_logic;
signal \N__14693\ : std_logic;
signal \N__14690\ : std_logic;
signal \N__14687\ : std_logic;
signal \N__14684\ : std_logic;
signal \N__14681\ : std_logic;
signal \N__14678\ : std_logic;
signal \N__14675\ : std_logic;
signal \N__14672\ : std_logic;
signal \N__14671\ : std_logic;
signal \N__14668\ : std_logic;
signal \N__14665\ : std_logic;
signal \N__14662\ : std_logic;
signal \N__14659\ : std_logic;
signal \N__14654\ : std_logic;
signal \N__14651\ : std_logic;
signal \N__14648\ : std_logic;
signal \N__14645\ : std_logic;
signal \N__14642\ : std_logic;
signal \N__14639\ : std_logic;
signal \N__14636\ : std_logic;
signal \N__14633\ : std_logic;
signal \N__14630\ : std_logic;
signal \N__14627\ : std_logic;
signal \N__14624\ : std_logic;
signal \N__14621\ : std_logic;
signal \N__14618\ : std_logic;
signal \N__14615\ : std_logic;
signal \N__14612\ : std_logic;
signal \N__14609\ : std_logic;
signal \N__14606\ : std_logic;
signal \N__14603\ : std_logic;
signal \N__14600\ : std_logic;
signal \N__14597\ : std_logic;
signal \N__14594\ : std_logic;
signal \N__14591\ : std_logic;
signal \N__14588\ : std_logic;
signal \N__14585\ : std_logic;
signal \N__14582\ : std_logic;
signal \N__14579\ : std_logic;
signal \N__14578\ : std_logic;
signal \N__14575\ : std_logic;
signal \N__14574\ : std_logic;
signal \N__14573\ : std_logic;
signal \N__14570\ : std_logic;
signal \N__14567\ : std_logic;
signal \N__14564\ : std_logic;
signal \N__14561\ : std_logic;
signal \N__14558\ : std_logic;
signal \N__14549\ : std_logic;
signal \N__14546\ : std_logic;
signal \N__14543\ : std_logic;
signal \N__14540\ : std_logic;
signal \N__14539\ : std_logic;
signal \N__14536\ : std_logic;
signal \N__14535\ : std_logic;
signal \N__14534\ : std_logic;
signal \N__14531\ : std_logic;
signal \N__14528\ : std_logic;
signal \N__14523\ : std_logic;
signal \N__14520\ : std_logic;
signal \N__14513\ : std_logic;
signal \N__14510\ : std_logic;
signal \N__14507\ : std_logic;
signal \N__14504\ : std_logic;
signal \N__14503\ : std_logic;
signal \N__14502\ : std_logic;
signal \N__14499\ : std_logic;
signal \N__14496\ : std_logic;
signal \N__14493\ : std_logic;
signal \N__14492\ : std_logic;
signal \N__14489\ : std_logic;
signal \N__14486\ : std_logic;
signal \N__14483\ : std_logic;
signal \N__14480\ : std_logic;
signal \N__14471\ : std_logic;
signal \N__14468\ : std_logic;
signal \N__14465\ : std_logic;
signal \N__14462\ : std_logic;
signal \N__14461\ : std_logic;
signal \N__14460\ : std_logic;
signal \N__14457\ : std_logic;
signal \N__14454\ : std_logic;
signal \N__14451\ : std_logic;
signal \N__14450\ : std_logic;
signal \N__14443\ : std_logic;
signal \N__14440\ : std_logic;
signal \N__14435\ : std_logic;
signal \N__14432\ : std_logic;
signal \N__14429\ : std_logic;
signal \N__14426\ : std_logic;
signal \N__14423\ : std_logic;
signal \N__14420\ : std_logic;
signal \N__14417\ : std_logic;
signal \N__14414\ : std_logic;
signal \N__14413\ : std_logic;
signal \N__14410\ : std_logic;
signal \N__14407\ : std_logic;
signal \N__14402\ : std_logic;
signal \N__14399\ : std_logic;
signal \N__14396\ : std_logic;
signal \N__14393\ : std_logic;
signal \N__14390\ : std_logic;
signal \N__14389\ : std_logic;
signal \N__14386\ : std_logic;
signal \N__14383\ : std_logic;
signal \N__14380\ : std_logic;
signal \N__14377\ : std_logic;
signal \N__14374\ : std_logic;
signal \N__14371\ : std_logic;
signal \N__14368\ : std_logic;
signal \N__14365\ : std_logic;
signal \N__14360\ : std_logic;
signal \N__14357\ : std_logic;
signal \N__14354\ : std_logic;
signal \N__14351\ : std_logic;
signal \N__14348\ : std_logic;
signal \N__14345\ : std_logic;
signal \N__14344\ : std_logic;
signal \N__14341\ : std_logic;
signal \N__14336\ : std_logic;
signal \N__14335\ : std_logic;
signal \N__14332\ : std_logic;
signal \N__14329\ : std_logic;
signal \N__14324\ : std_logic;
signal \N__14321\ : std_logic;
signal \N__14318\ : std_logic;
signal \N__14315\ : std_logic;
signal \N__14312\ : std_logic;
signal \N__14309\ : std_logic;
signal \N__14306\ : std_logic;
signal \N__14305\ : std_logic;
signal \N__14302\ : std_logic;
signal \N__14299\ : std_logic;
signal \N__14294\ : std_logic;
signal \N__14291\ : std_logic;
signal \N__14288\ : std_logic;
signal \N__14287\ : std_logic;
signal \N__14284\ : std_logic;
signal \N__14281\ : std_logic;
signal \N__14278\ : std_logic;
signal \N__14277\ : std_logic;
signal \N__14274\ : std_logic;
signal \N__14273\ : std_logic;
signal \N__14270\ : std_logic;
signal \N__14269\ : std_logic;
signal \N__14266\ : std_logic;
signal \N__14263\ : std_logic;
signal \N__14260\ : std_logic;
signal \N__14257\ : std_logic;
signal \N__14254\ : std_logic;
signal \N__14247\ : std_logic;
signal \N__14240\ : std_logic;
signal \N__14237\ : std_logic;
signal \N__14234\ : std_logic;
signal \N__14231\ : std_logic;
signal \N__14228\ : std_logic;
signal \N__14225\ : std_logic;
signal \N__14222\ : std_logic;
signal \N__14219\ : std_logic;
signal \N__14216\ : std_logic;
signal \N__14213\ : std_logic;
signal \N__14212\ : std_logic;
signal \N__14211\ : std_logic;
signal \N__14210\ : std_logic;
signal \N__14207\ : std_logic;
signal \N__14204\ : std_logic;
signal \N__14201\ : std_logic;
signal \N__14198\ : std_logic;
signal \N__14195\ : std_logic;
signal \N__14190\ : std_logic;
signal \N__14187\ : std_logic;
signal \N__14180\ : std_logic;
signal \N__14177\ : std_logic;
signal \N__14176\ : std_logic;
signal \N__14173\ : std_logic;
signal \N__14170\ : std_logic;
signal \N__14165\ : std_logic;
signal \N__14164\ : std_logic;
signal \N__14161\ : std_logic;
signal \N__14158\ : std_logic;
signal \N__14155\ : std_logic;
signal \N__14152\ : std_logic;
signal \N__14149\ : std_logic;
signal \N__14144\ : std_logic;
signal \N__14141\ : std_logic;
signal \N__14138\ : std_logic;
signal \N__14135\ : std_logic;
signal \N__14132\ : std_logic;
signal \N__14129\ : std_logic;
signal \N__14126\ : std_logic;
signal \N__14125\ : std_logic;
signal \N__14122\ : std_logic;
signal \N__14119\ : std_logic;
signal \N__14114\ : std_logic;
signal \N__14113\ : std_logic;
signal \N__14110\ : std_logic;
signal \N__14107\ : std_logic;
signal \N__14104\ : std_logic;
signal \N__14101\ : std_logic;
signal \N__14098\ : std_logic;
signal \N__14095\ : std_logic;
signal \N__14092\ : std_logic;
signal \N__14089\ : std_logic;
signal \N__14086\ : std_logic;
signal \N__14083\ : std_logic;
signal \N__14080\ : std_logic;
signal \N__14077\ : std_logic;
signal \N__14074\ : std_logic;
signal \N__14071\ : std_logic;
signal \N__14068\ : std_logic;
signal \N__14065\ : std_logic;
signal \N__14062\ : std_logic;
signal \N__14059\ : std_logic;
signal \N__14056\ : std_logic;
signal \N__14053\ : std_logic;
signal \N__14050\ : std_logic;
signal \N__14047\ : std_logic;
signal \N__14044\ : std_logic;
signal \N__14041\ : std_logic;
signal \N__14038\ : std_logic;
signal \N__14035\ : std_logic;
signal \N__14032\ : std_logic;
signal \N__14029\ : std_logic;
signal \N__14026\ : std_logic;
signal \N__14023\ : std_logic;
signal \N__14020\ : std_logic;
signal \N__14017\ : std_logic;
signal \N__14014\ : std_logic;
signal \N__14011\ : std_logic;
signal \N__14008\ : std_logic;
signal \N__14005\ : std_logic;
signal \N__14002\ : std_logic;
signal \N__13999\ : std_logic;
signal \N__13996\ : std_logic;
signal \N__13993\ : std_logic;
signal \N__13990\ : std_logic;
signal \N__13987\ : std_logic;
signal \N__13984\ : std_logic;
signal \N__13981\ : std_logic;
signal \N__13978\ : std_logic;
signal \N__13975\ : std_logic;
signal \N__13972\ : std_logic;
signal \N__13969\ : std_logic;
signal \N__13966\ : std_logic;
signal \N__13963\ : std_logic;
signal \N__13960\ : std_logic;
signal \N__13957\ : std_logic;
signal \N__13954\ : std_logic;
signal \N__13951\ : std_logic;
signal \N__13948\ : std_logic;
signal \N__13945\ : std_logic;
signal \N__13942\ : std_logic;
signal \N__13939\ : std_logic;
signal \N__13936\ : std_logic;
signal \N__13933\ : std_logic;
signal \N__13930\ : std_logic;
signal \N__13927\ : std_logic;
signal \N__13924\ : std_logic;
signal \N__13921\ : std_logic;
signal \N__13918\ : std_logic;
signal \N__13915\ : std_logic;
signal \N__13912\ : std_logic;
signal \N__13909\ : std_logic;
signal \N__13906\ : std_logic;
signal \N__13903\ : std_logic;
signal \N__13900\ : std_logic;
signal \N__13895\ : std_logic;
signal \N__13894\ : std_logic;
signal \N__13891\ : std_logic;
signal \N__13888\ : std_logic;
signal \N__13883\ : std_logic;
signal \N__13880\ : std_logic;
signal \N__13877\ : std_logic;
signal \N__13874\ : std_logic;
signal \N__13871\ : std_logic;
signal \N__13870\ : std_logic;
signal \N__13867\ : std_logic;
signal \N__13864\ : std_logic;
signal \N__13861\ : std_logic;
signal \N__13858\ : std_logic;
signal \N__13855\ : std_logic;
signal \N__13852\ : std_logic;
signal \N__13849\ : std_logic;
signal \N__13846\ : std_logic;
signal \N__13843\ : std_logic;
signal \N__13840\ : std_logic;
signal \N__13837\ : std_logic;
signal \N__13834\ : std_logic;
signal \N__13831\ : std_logic;
signal \N__13828\ : std_logic;
signal \N__13825\ : std_logic;
signal \N__13822\ : std_logic;
signal \N__13819\ : std_logic;
signal \N__13816\ : std_logic;
signal \N__13813\ : std_logic;
signal \N__13810\ : std_logic;
signal \N__13807\ : std_logic;
signal \N__13804\ : std_logic;
signal \N__13801\ : std_logic;
signal \N__13798\ : std_logic;
signal \N__13795\ : std_logic;
signal \N__13792\ : std_logic;
signal \N__13789\ : std_logic;
signal \N__13786\ : std_logic;
signal \N__13783\ : std_logic;
signal \N__13780\ : std_logic;
signal \N__13777\ : std_logic;
signal \N__13774\ : std_logic;
signal \N__13771\ : std_logic;
signal \N__13768\ : std_logic;
signal \N__13765\ : std_logic;
signal \N__13762\ : std_logic;
signal \N__13759\ : std_logic;
signal \N__13756\ : std_logic;
signal \N__13753\ : std_logic;
signal \N__13750\ : std_logic;
signal \N__13747\ : std_logic;
signal \N__13744\ : std_logic;
signal \N__13741\ : std_logic;
signal \N__13738\ : std_logic;
signal \N__13735\ : std_logic;
signal \N__13732\ : std_logic;
signal \N__13729\ : std_logic;
signal \N__13726\ : std_logic;
signal \N__13723\ : std_logic;
signal \N__13720\ : std_logic;
signal \N__13717\ : std_logic;
signal \N__13714\ : std_logic;
signal \N__13711\ : std_logic;
signal \N__13708\ : std_logic;
signal \N__13705\ : std_logic;
signal \N__13702\ : std_logic;
signal \N__13699\ : std_logic;
signal \N__13696\ : std_logic;
signal \N__13693\ : std_logic;
signal \N__13690\ : std_logic;
signal \N__13687\ : std_logic;
signal \N__13684\ : std_logic;
signal \N__13681\ : std_logic;
signal \N__13678\ : std_logic;
signal \N__13675\ : std_logic;
signal \N__13672\ : std_logic;
signal \N__13669\ : std_logic;
signal \N__13666\ : std_logic;
signal \N__13661\ : std_logic;
signal \N__13658\ : std_logic;
signal \N__13655\ : std_logic;
signal \N__13652\ : std_logic;
signal \N__13649\ : std_logic;
signal \N__13646\ : std_logic;
signal \N__13643\ : std_logic;
signal \N__13640\ : std_logic;
signal \N__13637\ : std_logic;
signal \N__13634\ : std_logic;
signal \N__13631\ : std_logic;
signal \N__13628\ : std_logic;
signal \N__13625\ : std_logic;
signal \N__13622\ : std_logic;
signal \N__13619\ : std_logic;
signal \N__13616\ : std_logic;
signal \N__13615\ : std_logic;
signal \N__13612\ : std_logic;
signal \N__13609\ : std_logic;
signal \N__13604\ : std_logic;
signal \N__13601\ : std_logic;
signal \N__13600\ : std_logic;
signal \N__13597\ : std_logic;
signal \N__13594\ : std_logic;
signal \N__13591\ : std_logic;
signal \N__13586\ : std_logic;
signal \N__13583\ : std_logic;
signal \N__13580\ : std_logic;
signal \N__13577\ : std_logic;
signal \N__13574\ : std_logic;
signal \N__13571\ : std_logic;
signal \N__13568\ : std_logic;
signal \N__13565\ : std_logic;
signal \N__13562\ : std_logic;
signal \N__13559\ : std_logic;
signal \N__13556\ : std_logic;
signal \N__13553\ : std_logic;
signal \N__13550\ : std_logic;
signal \N__13547\ : std_logic;
signal \N__13544\ : std_logic;
signal \N__13541\ : std_logic;
signal \N__13538\ : std_logic;
signal \N__13535\ : std_logic;
signal \N__13534\ : std_logic;
signal \N__13533\ : std_logic;
signal \N__13532\ : std_logic;
signal \N__13529\ : std_logic;
signal \N__13526\ : std_logic;
signal \N__13523\ : std_logic;
signal \N__13520\ : std_logic;
signal \N__13511\ : std_logic;
signal \N__13508\ : std_logic;
signal \N__13505\ : std_logic;
signal \N__13502\ : std_logic;
signal \N__13499\ : std_logic;
signal \N__13496\ : std_logic;
signal \N__13493\ : std_logic;
signal \N__13490\ : std_logic;
signal \N__13487\ : std_logic;
signal \N__13486\ : std_logic;
signal \N__13483\ : std_logic;
signal \N__13482\ : std_logic;
signal \N__13479\ : std_logic;
signal \N__13478\ : std_logic;
signal \N__13475\ : std_logic;
signal \N__13472\ : std_logic;
signal \N__13469\ : std_logic;
signal \N__13466\ : std_logic;
signal \N__13457\ : std_logic;
signal \N__13454\ : std_logic;
signal \N__13451\ : std_logic;
signal \N__13448\ : std_logic;
signal \N__13445\ : std_logic;
signal \N__13442\ : std_logic;
signal \N__13439\ : std_logic;
signal \N__13436\ : std_logic;
signal \N__13433\ : std_logic;
signal \N__13430\ : std_logic;
signal \N__13427\ : std_logic;
signal \N__13424\ : std_logic;
signal \N__13421\ : std_logic;
signal \N__13418\ : std_logic;
signal \N__13415\ : std_logic;
signal \N__13414\ : std_logic;
signal \N__13413\ : std_logic;
signal \N__13410\ : std_logic;
signal \N__13407\ : std_logic;
signal \N__13404\ : std_logic;
signal \N__13403\ : std_logic;
signal \N__13396\ : std_logic;
signal \N__13393\ : std_logic;
signal \N__13390\ : std_logic;
signal \N__13387\ : std_logic;
signal \N__13384\ : std_logic;
signal \N__13381\ : std_logic;
signal \N__13378\ : std_logic;
signal \N__13375\ : std_logic;
signal \N__13370\ : std_logic;
signal \N__13367\ : std_logic;
signal \N__13364\ : std_logic;
signal \N__13361\ : std_logic;
signal \N__13358\ : std_logic;
signal \N__13355\ : std_logic;
signal \N__13352\ : std_logic;
signal \N__13349\ : std_logic;
signal \N__13346\ : std_logic;
signal \N__13343\ : std_logic;
signal \N__13340\ : std_logic;
signal \N__13337\ : std_logic;
signal \N__13334\ : std_logic;
signal \N__13331\ : std_logic;
signal \N__13328\ : std_logic;
signal \N__13325\ : std_logic;
signal \N__13322\ : std_logic;
signal \N__13319\ : std_logic;
signal \N__13316\ : std_logic;
signal \N__13313\ : std_logic;
signal \N__13310\ : std_logic;
signal \N__13309\ : std_logic;
signal \N__13306\ : std_logic;
signal \N__13305\ : std_logic;
signal \N__13304\ : std_logic;
signal \N__13301\ : std_logic;
signal \N__13298\ : std_logic;
signal \N__13293\ : std_logic;
signal \N__13286\ : std_logic;
signal \N__13283\ : std_logic;
signal \N__13280\ : std_logic;
signal \N__13279\ : std_logic;
signal \N__13276\ : std_logic;
signal \N__13273\ : std_logic;
signal \N__13268\ : std_logic;
signal \N__13265\ : std_logic;
signal \N__13264\ : std_logic;
signal \N__13263\ : std_logic;
signal \N__13262\ : std_logic;
signal \N__13259\ : std_logic;
signal \N__13256\ : std_logic;
signal \N__13253\ : std_logic;
signal \N__13250\ : std_logic;
signal \N__13247\ : std_logic;
signal \N__13238\ : std_logic;
signal \N__13235\ : std_logic;
signal \N__13232\ : std_logic;
signal \N__13229\ : std_logic;
signal \N__13226\ : std_logic;
signal \N__13223\ : std_logic;
signal \N__13220\ : std_logic;
signal \N__13219\ : std_logic;
signal \N__13218\ : std_logic;
signal \N__13217\ : std_logic;
signal \N__13214\ : std_logic;
signal \N__13211\ : std_logic;
signal \N__13206\ : std_logic;
signal \N__13199\ : std_logic;
signal \N__13198\ : std_logic;
signal \N__13195\ : std_logic;
signal \N__13194\ : std_logic;
signal \N__13193\ : std_logic;
signal \N__13190\ : std_logic;
signal \N__13187\ : std_logic;
signal \N__13184\ : std_logic;
signal \N__13181\ : std_logic;
signal \N__13178\ : std_logic;
signal \N__13169\ : std_logic;
signal \N__13166\ : std_logic;
signal \N__13165\ : std_logic;
signal \N__13164\ : std_logic;
signal \N__13163\ : std_logic;
signal \N__13160\ : std_logic;
signal \N__13157\ : std_logic;
signal \N__13152\ : std_logic;
signal \N__13145\ : std_logic;
signal \N__13142\ : std_logic;
signal \N__13139\ : std_logic;
signal \N__13136\ : std_logic;
signal \N__13135\ : std_logic;
signal \N__13134\ : std_logic;
signal \N__13133\ : std_logic;
signal \N__13130\ : std_logic;
signal \N__13127\ : std_logic;
signal \N__13122\ : std_logic;
signal \N__13115\ : std_logic;
signal \N__13114\ : std_logic;
signal \N__13111\ : std_logic;
signal \N__13110\ : std_logic;
signal \N__13109\ : std_logic;
signal \N__13106\ : std_logic;
signal \N__13103\ : std_logic;
signal \N__13100\ : std_logic;
signal \N__13097\ : std_logic;
signal \N__13088\ : std_logic;
signal \N__13085\ : std_logic;
signal \N__13082\ : std_logic;
signal \N__13079\ : std_logic;
signal \N__13076\ : std_logic;
signal \N__13073\ : std_logic;
signal \N__13072\ : std_logic;
signal \N__13071\ : std_logic;
signal \N__13068\ : std_logic;
signal \N__13065\ : std_logic;
signal \N__13062\ : std_logic;
signal \N__13061\ : std_logic;
signal \N__13054\ : std_logic;
signal \N__13051\ : std_logic;
signal \N__13048\ : std_logic;
signal \N__13045\ : std_logic;
signal \N__13040\ : std_logic;
signal \N__13037\ : std_logic;
signal \N__13034\ : std_logic;
signal \N__13031\ : std_logic;
signal \N__13028\ : std_logic;
signal \N__13025\ : std_logic;
signal \N__13024\ : std_logic;
signal \N__13021\ : std_logic;
signal \N__13018\ : std_logic;
signal \N__13017\ : std_logic;
signal \N__13016\ : std_logic;
signal \N__13011\ : std_logic;
signal \N__13008\ : std_logic;
signal \N__13005\ : std_logic;
signal \N__12998\ : std_logic;
signal \N__12995\ : std_logic;
signal \N__12992\ : std_logic;
signal \N__12989\ : std_logic;
signal \N__12988\ : std_logic;
signal \N__12987\ : std_logic;
signal \N__12984\ : std_logic;
signal \N__12981\ : std_logic;
signal \N__12978\ : std_logic;
signal \N__12971\ : std_logic;
signal \N__12970\ : std_logic;
signal \N__12969\ : std_logic;
signal \N__12966\ : std_logic;
signal \N__12963\ : std_logic;
signal \N__12960\ : std_logic;
signal \N__12953\ : std_logic;
signal \N__12952\ : std_logic;
signal \N__12951\ : std_logic;
signal \N__12948\ : std_logic;
signal \N__12945\ : std_logic;
signal \N__12942\ : std_logic;
signal \N__12935\ : std_logic;
signal \N__12932\ : std_logic;
signal \N__12929\ : std_logic;
signal \N__12926\ : std_logic;
signal \N__12923\ : std_logic;
signal \N__12920\ : std_logic;
signal \N__12917\ : std_logic;
signal \N__12914\ : std_logic;
signal \N__12913\ : std_logic;
signal \N__12910\ : std_logic;
signal \N__12907\ : std_logic;
signal \N__12902\ : std_logic;
signal \N__12901\ : std_logic;
signal \N__12900\ : std_logic;
signal \N__12897\ : std_logic;
signal \N__12894\ : std_logic;
signal \N__12891\ : std_logic;
signal \N__12890\ : std_logic;
signal \N__12887\ : std_logic;
signal \N__12882\ : std_logic;
signal \N__12879\ : std_logic;
signal \N__12876\ : std_logic;
signal \N__12871\ : std_logic;
signal \N__12866\ : std_logic;
signal \N__12863\ : std_logic;
signal \N__12860\ : std_logic;
signal \N__12857\ : std_logic;
signal \N__12854\ : std_logic;
signal \N__12853\ : std_logic;
signal \N__12852\ : std_logic;
signal \N__12849\ : std_logic;
signal \N__12846\ : std_logic;
signal \N__12843\ : std_logic;
signal \N__12836\ : std_logic;
signal \N__12835\ : std_logic;
signal \N__12832\ : std_logic;
signal \N__12829\ : std_logic;
signal \N__12826\ : std_logic;
signal \N__12821\ : std_logic;
signal \N__12818\ : std_logic;
signal \N__12815\ : std_logic;
signal \N__12812\ : std_logic;
signal \N__12811\ : std_logic;
signal \N__12810\ : std_logic;
signal \N__12807\ : std_logic;
signal \N__12804\ : std_logic;
signal \N__12801\ : std_logic;
signal \N__12794\ : std_logic;
signal \N__12793\ : std_logic;
signal \N__12792\ : std_logic;
signal \N__12789\ : std_logic;
signal \N__12786\ : std_logic;
signal \N__12783\ : std_logic;
signal \N__12776\ : std_logic;
signal \N__12773\ : std_logic;
signal \N__12770\ : std_logic;
signal \N__12767\ : std_logic;
signal \N__12764\ : std_logic;
signal \N__12761\ : std_logic;
signal \N__12758\ : std_logic;
signal \N__12755\ : std_logic;
signal \N__12752\ : std_logic;
signal \N__12749\ : std_logic;
signal \N__12746\ : std_logic;
signal \N__12743\ : std_logic;
signal \N__12740\ : std_logic;
signal \N__12737\ : std_logic;
signal \N__12734\ : std_logic;
signal \N__12731\ : std_logic;
signal \N__12728\ : std_logic;
signal \N__12727\ : std_logic;
signal \N__12726\ : std_logic;
signal \N__12723\ : std_logic;
signal \N__12720\ : std_logic;
signal \N__12717\ : std_logic;
signal \N__12714\ : std_logic;
signal \N__12711\ : std_logic;
signal \N__12708\ : std_logic;
signal \N__12705\ : std_logic;
signal \N__12702\ : std_logic;
signal \N__12699\ : std_logic;
signal \N__12696\ : std_logic;
signal \N__12693\ : std_logic;
signal \N__12690\ : std_logic;
signal \N__12687\ : std_logic;
signal \N__12684\ : std_logic;
signal \N__12677\ : std_logic;
signal \N__12674\ : std_logic;
signal \N__12671\ : std_logic;
signal \N__12668\ : std_logic;
signal \N__12665\ : std_logic;
signal \N__12662\ : std_logic;
signal \N__12659\ : std_logic;
signal \N__12656\ : std_logic;
signal \N__12653\ : std_logic;
signal \N__12650\ : std_logic;
signal \N__12647\ : std_logic;
signal \N__12644\ : std_logic;
signal \N__12641\ : std_logic;
signal \N__12640\ : std_logic;
signal \N__12639\ : std_logic;
signal \N__12636\ : std_logic;
signal \N__12633\ : std_logic;
signal \N__12630\ : std_logic;
signal \N__12627\ : std_logic;
signal \N__12626\ : std_logic;
signal \N__12623\ : std_logic;
signal \N__12620\ : std_logic;
signal \N__12617\ : std_logic;
signal \N__12614\ : std_logic;
signal \N__12611\ : std_logic;
signal \N__12608\ : std_logic;
signal \N__12603\ : std_logic;
signal \N__12600\ : std_logic;
signal \N__12597\ : std_logic;
signal \N__12594\ : std_logic;
signal \N__12591\ : std_logic;
signal \N__12588\ : std_logic;
signal \N__12585\ : std_logic;
signal \N__12578\ : std_logic;
signal \N__12577\ : std_logic;
signal \N__12574\ : std_logic;
signal \N__12571\ : std_logic;
signal \N__12566\ : std_logic;
signal \N__12565\ : std_logic;
signal \N__12562\ : std_logic;
signal \N__12559\ : std_logic;
signal \N__12554\ : std_logic;
signal \N__12553\ : std_logic;
signal \N__12550\ : std_logic;
signal \N__12547\ : std_logic;
signal \N__12542\ : std_logic;
signal \N__12539\ : std_logic;
signal \N__12536\ : std_logic;
signal \N__12535\ : std_logic;
signal \N__12534\ : std_logic;
signal \N__12531\ : std_logic;
signal \N__12526\ : std_logic;
signal \N__12521\ : std_logic;
signal \N__12520\ : std_logic;
signal \N__12519\ : std_logic;
signal \N__12516\ : std_logic;
signal \N__12511\ : std_logic;
signal \N__12506\ : std_logic;
signal \N__12503\ : std_logic;
signal \N__12502\ : std_logic;
signal \N__12499\ : std_logic;
signal \N__12496\ : std_logic;
signal \N__12493\ : std_logic;
signal \N__12490\ : std_logic;
signal \N__12485\ : std_logic;
signal \N__12484\ : std_logic;
signal \N__12483\ : std_logic;
signal \N__12480\ : std_logic;
signal \N__12477\ : std_logic;
signal \N__12474\ : std_logic;
signal \N__12473\ : std_logic;
signal \N__12468\ : std_logic;
signal \N__12463\ : std_logic;
signal \N__12458\ : std_logic;
signal \N__12457\ : std_logic;
signal \N__12456\ : std_logic;
signal \N__12455\ : std_logic;
signal \N__12452\ : std_logic;
signal \N__12449\ : std_logic;
signal \N__12444\ : std_logic;
signal \N__12439\ : std_logic;
signal \N__12434\ : std_logic;
signal \N__12431\ : std_logic;
signal \N__12428\ : std_logic;
signal \N__12427\ : std_logic;
signal \N__12424\ : std_logic;
signal \N__12421\ : std_logic;
signal \N__12416\ : std_logic;
signal \N__12415\ : std_logic;
signal \N__12412\ : std_logic;
signal \N__12409\ : std_logic;
signal \N__12408\ : std_logic;
signal \N__12407\ : std_logic;
signal \N__12406\ : std_logic;
signal \N__12403\ : std_logic;
signal \N__12400\ : std_logic;
signal \N__12397\ : std_logic;
signal \N__12394\ : std_logic;
signal \N__12391\ : std_logic;
signal \N__12384\ : std_logic;
signal \N__12377\ : std_logic;
signal \N__12374\ : std_logic;
signal \N__12371\ : std_logic;
signal \N__12370\ : std_logic;
signal \N__12367\ : std_logic;
signal \N__12364\ : std_logic;
signal \N__12359\ : std_logic;
signal \N__12356\ : std_logic;
signal \N__12355\ : std_logic;
signal \N__12352\ : std_logic;
signal \N__12349\ : std_logic;
signal \N__12346\ : std_logic;
signal \N__12343\ : std_logic;
signal \N__12340\ : std_logic;
signal \N__12337\ : std_logic;
signal \N__12334\ : std_logic;
signal \N__12331\ : std_logic;
signal \N__12328\ : std_logic;
signal \N__12325\ : std_logic;
signal \N__12322\ : std_logic;
signal \N__12319\ : std_logic;
signal \N__12316\ : std_logic;
signal \N__12313\ : std_logic;
signal \N__12310\ : std_logic;
signal \N__12307\ : std_logic;
signal \N__12304\ : std_logic;
signal \N__12301\ : std_logic;
signal \N__12298\ : std_logic;
signal \N__12295\ : std_logic;
signal \N__12292\ : std_logic;
signal \N__12289\ : std_logic;
signal \N__12286\ : std_logic;
signal \N__12283\ : std_logic;
signal \N__12280\ : std_logic;
signal \N__12277\ : std_logic;
signal \N__12274\ : std_logic;
signal \N__12271\ : std_logic;
signal \N__12268\ : std_logic;
signal \N__12265\ : std_logic;
signal \N__12262\ : std_logic;
signal \N__12259\ : std_logic;
signal \N__12256\ : std_logic;
signal \N__12253\ : std_logic;
signal \N__12250\ : std_logic;
signal \N__12247\ : std_logic;
signal \N__12244\ : std_logic;
signal \N__12241\ : std_logic;
signal \N__12238\ : std_logic;
signal \N__12235\ : std_logic;
signal \N__12232\ : std_logic;
signal \N__12229\ : std_logic;
signal \N__12226\ : std_logic;
signal \N__12223\ : std_logic;
signal \N__12220\ : std_logic;
signal \N__12217\ : std_logic;
signal \N__12214\ : std_logic;
signal \N__12211\ : std_logic;
signal \N__12208\ : std_logic;
signal \N__12205\ : std_logic;
signal \N__12202\ : std_logic;
signal \N__12199\ : std_logic;
signal \N__12196\ : std_logic;
signal \N__12193\ : std_logic;
signal \N__12190\ : std_logic;
signal \N__12187\ : std_logic;
signal \N__12184\ : std_logic;
signal \N__12181\ : std_logic;
signal \N__12178\ : std_logic;
signal \N__12175\ : std_logic;
signal \N__12172\ : std_logic;
signal \N__12169\ : std_logic;
signal \N__12166\ : std_logic;
signal \N__12163\ : std_logic;
signal \N__12160\ : std_logic;
signal \N__12157\ : std_logic;
signal \N__12154\ : std_logic;
signal \N__12151\ : std_logic;
signal \N__12148\ : std_logic;
signal \N__12145\ : std_logic;
signal \N__12140\ : std_logic;
signal \N__12137\ : std_logic;
signal \N__12134\ : std_logic;
signal \N__12131\ : std_logic;
signal \N__12128\ : std_logic;
signal \N__12125\ : std_logic;
signal \N__12122\ : std_logic;
signal \N__12119\ : std_logic;
signal \N__12116\ : std_logic;
signal \N__12113\ : std_logic;
signal \N__12110\ : std_logic;
signal \N__12107\ : std_logic;
signal \N__12104\ : std_logic;
signal \N__12103\ : std_logic;
signal \N__12098\ : std_logic;
signal \N__12095\ : std_logic;
signal \N__12092\ : std_logic;
signal \N__12091\ : std_logic;
signal \N__12088\ : std_logic;
signal \N__12085\ : std_logic;
signal \N__12082\ : std_logic;
signal \N__12079\ : std_logic;
signal \N__12076\ : std_logic;
signal \N__12073\ : std_logic;
signal \N__12070\ : std_logic;
signal \N__12067\ : std_logic;
signal \N__12064\ : std_logic;
signal \N__12061\ : std_logic;
signal \N__12058\ : std_logic;
signal \N__12055\ : std_logic;
signal \N__12052\ : std_logic;
signal \N__12049\ : std_logic;
signal \N__12046\ : std_logic;
signal \N__12043\ : std_logic;
signal \N__12040\ : std_logic;
signal \N__12037\ : std_logic;
signal \N__12034\ : std_logic;
signal \N__12031\ : std_logic;
signal \N__12028\ : std_logic;
signal \N__12025\ : std_logic;
signal \N__12022\ : std_logic;
signal \N__12019\ : std_logic;
signal \N__12016\ : std_logic;
signal \N__12013\ : std_logic;
signal \N__12010\ : std_logic;
signal \N__12007\ : std_logic;
signal \N__12004\ : std_logic;
signal \N__12001\ : std_logic;
signal \N__11998\ : std_logic;
signal \N__11995\ : std_logic;
signal \N__11992\ : std_logic;
signal \N__11989\ : std_logic;
signal \N__11986\ : std_logic;
signal \N__11983\ : std_logic;
signal \N__11980\ : std_logic;
signal \N__11977\ : std_logic;
signal \N__11974\ : std_logic;
signal \N__11971\ : std_logic;
signal \N__11968\ : std_logic;
signal \N__11965\ : std_logic;
signal \N__11962\ : std_logic;
signal \N__11959\ : std_logic;
signal \N__11956\ : std_logic;
signal \N__11953\ : std_logic;
signal \N__11950\ : std_logic;
signal \N__11947\ : std_logic;
signal \N__11944\ : std_logic;
signal \N__11941\ : std_logic;
signal \N__11938\ : std_logic;
signal \N__11935\ : std_logic;
signal \N__11932\ : std_logic;
signal \N__11929\ : std_logic;
signal \N__11926\ : std_logic;
signal \N__11923\ : std_logic;
signal \N__11920\ : std_logic;
signal \N__11917\ : std_logic;
signal \N__11914\ : std_logic;
signal \N__11911\ : std_logic;
signal \N__11908\ : std_logic;
signal \N__11905\ : std_logic;
signal \N__11902\ : std_logic;
signal \N__11899\ : std_logic;
signal \N__11896\ : std_logic;
signal \N__11893\ : std_logic;
signal \N__11890\ : std_logic;
signal \N__11887\ : std_logic;
signal \N__11884\ : std_logic;
signal \N__11881\ : std_logic;
signal \N__11878\ : std_logic;
signal \N__11873\ : std_logic;
signal \N__11872\ : std_logic;
signal \N__11869\ : std_logic;
signal \N__11866\ : std_logic;
signal \N__11861\ : std_logic;
signal \N__11860\ : std_logic;
signal \N__11857\ : std_logic;
signal \N__11856\ : std_logic;
signal \N__11853\ : std_logic;
signal \N__11850\ : std_logic;
signal \N__11847\ : std_logic;
signal \N__11846\ : std_logic;
signal \N__11843\ : std_logic;
signal \N__11840\ : std_logic;
signal \N__11837\ : std_logic;
signal \N__11834\ : std_logic;
signal \N__11829\ : std_logic;
signal \N__11826\ : std_logic;
signal \N__11819\ : std_logic;
signal \N__11818\ : std_logic;
signal \N__11815\ : std_logic;
signal \N__11812\ : std_logic;
signal \N__11809\ : std_logic;
signal \N__11804\ : std_logic;
signal \N__11801\ : std_logic;
signal \N__11800\ : std_logic;
signal \N__11797\ : std_logic;
signal \N__11794\ : std_logic;
signal \N__11789\ : std_logic;
signal \N__11786\ : std_logic;
signal \N__11783\ : std_logic;
signal \N__11780\ : std_logic;
signal \N__11779\ : std_logic;
signal \N__11776\ : std_logic;
signal \N__11773\ : std_logic;
signal \N__11770\ : std_logic;
signal \N__11767\ : std_logic;
signal \N__11764\ : std_logic;
signal \N__11761\ : std_logic;
signal \N__11758\ : std_logic;
signal \N__11755\ : std_logic;
signal \N__11752\ : std_logic;
signal \N__11749\ : std_logic;
signal \N__11746\ : std_logic;
signal \N__11743\ : std_logic;
signal \N__11740\ : std_logic;
signal \N__11737\ : std_logic;
signal \N__11734\ : std_logic;
signal \N__11731\ : std_logic;
signal \N__11728\ : std_logic;
signal \N__11725\ : std_logic;
signal \N__11722\ : std_logic;
signal \N__11719\ : std_logic;
signal \N__11716\ : std_logic;
signal \N__11713\ : std_logic;
signal \N__11710\ : std_logic;
signal \N__11707\ : std_logic;
signal \N__11704\ : std_logic;
signal \N__11701\ : std_logic;
signal \N__11698\ : std_logic;
signal \N__11695\ : std_logic;
signal \N__11692\ : std_logic;
signal \N__11689\ : std_logic;
signal \N__11686\ : std_logic;
signal \N__11683\ : std_logic;
signal \N__11680\ : std_logic;
signal \N__11677\ : std_logic;
signal \N__11674\ : std_logic;
signal \N__11671\ : std_logic;
signal \N__11668\ : std_logic;
signal \N__11665\ : std_logic;
signal \N__11662\ : std_logic;
signal \N__11659\ : std_logic;
signal \N__11656\ : std_logic;
signal \N__11653\ : std_logic;
signal \N__11650\ : std_logic;
signal \N__11647\ : std_logic;
signal \N__11644\ : std_logic;
signal \N__11641\ : std_logic;
signal \N__11638\ : std_logic;
signal \N__11635\ : std_logic;
signal \N__11632\ : std_logic;
signal \N__11629\ : std_logic;
signal \N__11626\ : std_logic;
signal \N__11623\ : std_logic;
signal \N__11620\ : std_logic;
signal \N__11617\ : std_logic;
signal \N__11614\ : std_logic;
signal \N__11611\ : std_logic;
signal \N__11608\ : std_logic;
signal \N__11605\ : std_logic;
signal \N__11602\ : std_logic;
signal \N__11599\ : std_logic;
signal \N__11596\ : std_logic;
signal \N__11593\ : std_logic;
signal \N__11590\ : std_logic;
signal \N__11587\ : std_logic;
signal \N__11584\ : std_logic;
signal \N__11581\ : std_logic;
signal \N__11578\ : std_logic;
signal \N__11575\ : std_logic;
signal \N__11572\ : std_logic;
signal \N__11569\ : std_logic;
signal \N__11566\ : std_logic;
signal \N__11563\ : std_logic;
signal \N__11560\ : std_logic;
signal \N__11555\ : std_logic;
signal \N__11554\ : std_logic;
signal \N__11549\ : std_logic;
signal \N__11548\ : std_logic;
signal \N__11545\ : std_logic;
signal \N__11544\ : std_logic;
signal \N__11543\ : std_logic;
signal \N__11540\ : std_logic;
signal \N__11537\ : std_logic;
signal \N__11534\ : std_logic;
signal \N__11531\ : std_logic;
signal \N__11522\ : std_logic;
signal \N__11519\ : std_logic;
signal \N__11516\ : std_logic;
signal \N__11513\ : std_logic;
signal \N__11510\ : std_logic;
signal \N__11507\ : std_logic;
signal \N__11504\ : std_logic;
signal \N__11503\ : std_logic;
signal \N__11500\ : std_logic;
signal \N__11497\ : std_logic;
signal \N__11494\ : std_logic;
signal \N__11491\ : std_logic;
signal \N__11488\ : std_logic;
signal \N__11485\ : std_logic;
signal \N__11482\ : std_logic;
signal \N__11479\ : std_logic;
signal \N__11476\ : std_logic;
signal \N__11473\ : std_logic;
signal \N__11470\ : std_logic;
signal \N__11467\ : std_logic;
signal \N__11464\ : std_logic;
signal \N__11461\ : std_logic;
signal \N__11458\ : std_logic;
signal \N__11455\ : std_logic;
signal \N__11452\ : std_logic;
signal \N__11449\ : std_logic;
signal \N__11446\ : std_logic;
signal \N__11443\ : std_logic;
signal \N__11440\ : std_logic;
signal \N__11437\ : std_logic;
signal \N__11434\ : std_logic;
signal \N__11431\ : std_logic;
signal \N__11428\ : std_logic;
signal \N__11425\ : std_logic;
signal \N__11422\ : std_logic;
signal \N__11419\ : std_logic;
signal \N__11416\ : std_logic;
signal \N__11413\ : std_logic;
signal \N__11410\ : std_logic;
signal \N__11407\ : std_logic;
signal \N__11404\ : std_logic;
signal \N__11401\ : std_logic;
signal \N__11398\ : std_logic;
signal \N__11395\ : std_logic;
signal \N__11392\ : std_logic;
signal \N__11389\ : std_logic;
signal \N__11386\ : std_logic;
signal \N__11383\ : std_logic;
signal \N__11380\ : std_logic;
signal \N__11377\ : std_logic;
signal \N__11374\ : std_logic;
signal \N__11371\ : std_logic;
signal \N__11368\ : std_logic;
signal \N__11365\ : std_logic;
signal \N__11362\ : std_logic;
signal \N__11359\ : std_logic;
signal \N__11356\ : std_logic;
signal \N__11353\ : std_logic;
signal \N__11350\ : std_logic;
signal \N__11347\ : std_logic;
signal \N__11344\ : std_logic;
signal \N__11341\ : std_logic;
signal \N__11338\ : std_logic;
signal \N__11335\ : std_logic;
signal \N__11332\ : std_logic;
signal \N__11329\ : std_logic;
signal \N__11326\ : std_logic;
signal \N__11323\ : std_logic;
signal \N__11320\ : std_logic;
signal \N__11317\ : std_logic;
signal \N__11314\ : std_logic;
signal \N__11311\ : std_logic;
signal \N__11308\ : std_logic;
signal \N__11305\ : std_logic;
signal \N__11302\ : std_logic;
signal \N__11299\ : std_logic;
signal \N__11296\ : std_logic;
signal \N__11293\ : std_logic;
signal \N__11288\ : std_logic;
signal \N__11285\ : std_logic;
signal \N__11284\ : std_logic;
signal \N__11283\ : std_logic;
signal \N__11278\ : std_logic;
signal \N__11275\ : std_logic;
signal \N__11274\ : std_logic;
signal \N__11271\ : std_logic;
signal \N__11266\ : std_logic;
signal \N__11261\ : std_logic;
signal \N__11258\ : std_logic;
signal \N__11255\ : std_logic;
signal \N__11252\ : std_logic;
signal \N__11251\ : std_logic;
signal \N__11246\ : std_logic;
signal \N__11243\ : std_logic;
signal \N__11240\ : std_logic;
signal \N__11239\ : std_logic;
signal \N__11236\ : std_logic;
signal \N__11233\ : std_logic;
signal \N__11230\ : std_logic;
signal \N__11227\ : std_logic;
signal \N__11224\ : std_logic;
signal \N__11221\ : std_logic;
signal \N__11218\ : std_logic;
signal \N__11215\ : std_logic;
signal \N__11212\ : std_logic;
signal \N__11209\ : std_logic;
signal \N__11206\ : std_logic;
signal \N__11203\ : std_logic;
signal \N__11200\ : std_logic;
signal \N__11197\ : std_logic;
signal \N__11194\ : std_logic;
signal \N__11191\ : std_logic;
signal \N__11188\ : std_logic;
signal \N__11185\ : std_logic;
signal \N__11182\ : std_logic;
signal \N__11179\ : std_logic;
signal \N__11176\ : std_logic;
signal \N__11173\ : std_logic;
signal \N__11170\ : std_logic;
signal \N__11167\ : std_logic;
signal \N__11164\ : std_logic;
signal \N__11161\ : std_logic;
signal \N__11158\ : std_logic;
signal \N__11155\ : std_logic;
signal \N__11152\ : std_logic;
signal \N__11149\ : std_logic;
signal \N__11146\ : std_logic;
signal \N__11143\ : std_logic;
signal \N__11140\ : std_logic;
signal \N__11137\ : std_logic;
signal \N__11134\ : std_logic;
signal \N__11131\ : std_logic;
signal \N__11128\ : std_logic;
signal \N__11125\ : std_logic;
signal \N__11122\ : std_logic;
signal \N__11119\ : std_logic;
signal \N__11116\ : std_logic;
signal \N__11113\ : std_logic;
signal \N__11110\ : std_logic;
signal \N__11107\ : std_logic;
signal \N__11104\ : std_logic;
signal \N__11101\ : std_logic;
signal \N__11098\ : std_logic;
signal \N__11095\ : std_logic;
signal \N__11092\ : std_logic;
signal \N__11089\ : std_logic;
signal \N__11086\ : std_logic;
signal \N__11083\ : std_logic;
signal \N__11080\ : std_logic;
signal \N__11077\ : std_logic;
signal \N__11074\ : std_logic;
signal \N__11071\ : std_logic;
signal \N__11068\ : std_logic;
signal \N__11065\ : std_logic;
signal \N__11062\ : std_logic;
signal \N__11059\ : std_logic;
signal \N__11056\ : std_logic;
signal \N__11053\ : std_logic;
signal \N__11050\ : std_logic;
signal \N__11047\ : std_logic;
signal \N__11044\ : std_logic;
signal \N__11041\ : std_logic;
signal \N__11038\ : std_logic;
signal \N__11035\ : std_logic;
signal \N__11032\ : std_logic;
signal \N__11029\ : std_logic;
signal \N__11026\ : std_logic;
signal \N__11023\ : std_logic;
signal \N__11020\ : std_logic;
signal \N__11015\ : std_logic;
signal \N__11014\ : std_logic;
signal \N__11013\ : std_logic;
signal \N__11010\ : std_logic;
signal \N__11009\ : std_logic;
signal \N__11006\ : std_logic;
signal \N__11003\ : std_logic;
signal \N__11000\ : std_logic;
signal \N__10997\ : std_logic;
signal \N__10988\ : std_logic;
signal \N__10985\ : std_logic;
signal \N__10982\ : std_logic;
signal \N__10979\ : std_logic;
signal \N__10976\ : std_logic;
signal \N__10975\ : std_logic;
signal \N__10972\ : std_logic;
signal \N__10969\ : std_logic;
signal \N__10964\ : std_logic;
signal \N__10963\ : std_logic;
signal \N__10962\ : std_logic;
signal \N__10959\ : std_logic;
signal \N__10958\ : std_logic;
signal \N__10955\ : std_logic;
signal \N__10952\ : std_logic;
signal \N__10949\ : std_logic;
signal \N__10946\ : std_logic;
signal \N__10937\ : std_logic;
signal \N__10934\ : std_logic;
signal \N__10931\ : std_logic;
signal \N__10928\ : std_logic;
signal \N__10925\ : std_logic;
signal \N__10922\ : std_logic;
signal \N__10919\ : std_logic;
signal \N__10916\ : std_logic;
signal \N__10913\ : std_logic;
signal \N__10910\ : std_logic;
signal \N__10907\ : std_logic;
signal \N__10904\ : std_logic;
signal \N__10901\ : std_logic;
signal \N__10898\ : std_logic;
signal \N__10895\ : std_logic;
signal \N__10892\ : std_logic;
signal \N__10889\ : std_logic;
signal \N__10886\ : std_logic;
signal \N__10883\ : std_logic;
signal \N__10880\ : std_logic;
signal \N__10877\ : std_logic;
signal \N__10874\ : std_logic;
signal \N__10871\ : std_logic;
signal \N__10870\ : std_logic;
signal \N__10865\ : std_logic;
signal \N__10862\ : std_logic;
signal \N__10861\ : std_logic;
signal \N__10860\ : std_logic;
signal \N__10857\ : std_logic;
signal \N__10852\ : std_logic;
signal \N__10847\ : std_logic;
signal \N__10844\ : std_logic;
signal \N__10841\ : std_logic;
signal \N__10838\ : std_logic;
signal \N__10835\ : std_logic;
signal \N__10832\ : std_logic;
signal \N__10829\ : std_logic;
signal \N__10826\ : std_logic;
signal \N__10823\ : std_logic;
signal \N__10820\ : std_logic;
signal \N__10819\ : std_logic;
signal \N__10818\ : std_logic;
signal \N__10815\ : std_logic;
signal \N__10810\ : std_logic;
signal \N__10809\ : std_logic;
signal \N__10808\ : std_logic;
signal \N__10807\ : std_logic;
signal \N__10804\ : std_logic;
signal \N__10801\ : std_logic;
signal \N__10794\ : std_logic;
signal \N__10787\ : std_logic;
signal \N__10784\ : std_logic;
signal \N__10781\ : std_logic;
signal \N__10778\ : std_logic;
signal \N__10775\ : std_logic;
signal \N__10772\ : std_logic;
signal \N__10769\ : std_logic;
signal \N__10766\ : std_logic;
signal \N__10763\ : std_logic;
signal \N__10760\ : std_logic;
signal \N__10757\ : std_logic;
signal \N__10754\ : std_logic;
signal \N__10751\ : std_logic;
signal \N__10748\ : std_logic;
signal \N__10745\ : std_logic;
signal \N__10742\ : std_logic;
signal \N__10739\ : std_logic;
signal \N__10736\ : std_logic;
signal \N__10735\ : std_logic;
signal \N__10732\ : std_logic;
signal \N__10729\ : std_logic;
signal \N__10728\ : std_logic;
signal \N__10725\ : std_logic;
signal \N__10724\ : std_logic;
signal \N__10721\ : std_logic;
signal \N__10718\ : std_logic;
signal \N__10717\ : std_logic;
signal \N__10716\ : std_logic;
signal \N__10715\ : std_logic;
signal \N__10712\ : std_logic;
signal \N__10709\ : std_logic;
signal \N__10708\ : std_logic;
signal \N__10703\ : std_logic;
signal \N__10700\ : std_logic;
signal \N__10697\ : std_logic;
signal \N__10694\ : std_logic;
signal \N__10689\ : std_logic;
signal \N__10686\ : std_logic;
signal \N__10679\ : std_logic;
signal \N__10676\ : std_logic;
signal \N__10673\ : std_logic;
signal \N__10670\ : std_logic;
signal \N__10665\ : std_logic;
signal \N__10660\ : std_logic;
signal \N__10657\ : std_logic;
signal \N__10654\ : std_logic;
signal \N__10649\ : std_logic;
signal \N__10646\ : std_logic;
signal \N__10643\ : std_logic;
signal \N__10640\ : std_logic;
signal \N__10637\ : std_logic;
signal \N__10634\ : std_logic;
signal \N__10631\ : std_logic;
signal \N__10628\ : std_logic;
signal \N__10625\ : std_logic;
signal \N__10622\ : std_logic;
signal \N__10619\ : std_logic;
signal \N__10616\ : std_logic;
signal \N__10613\ : std_logic;
signal \N__10610\ : std_logic;
signal \N__10609\ : std_logic;
signal \N__10606\ : std_logic;
signal \N__10603\ : std_logic;
signal \N__10602\ : std_logic;
signal \N__10601\ : std_logic;
signal \N__10600\ : std_logic;
signal \N__10599\ : std_logic;
signal \N__10596\ : std_logic;
signal \N__10595\ : std_logic;
signal \N__10594\ : std_logic;
signal \N__10591\ : std_logic;
signal \N__10588\ : std_logic;
signal \N__10585\ : std_logic;
signal \N__10582\ : std_logic;
signal \N__10579\ : std_logic;
signal \N__10576\ : std_logic;
signal \N__10573\ : std_logic;
signal \N__10570\ : std_logic;
signal \N__10565\ : std_logic;
signal \N__10560\ : std_logic;
signal \N__10557\ : std_logic;
signal \N__10552\ : std_logic;
signal \N__10549\ : std_logic;
signal \N__10546\ : std_logic;
signal \N__10541\ : std_logic;
signal \N__10536\ : std_logic;
signal \N__10531\ : std_logic;
signal \N__10528\ : std_logic;
signal \N__10523\ : std_logic;
signal \N__10520\ : std_logic;
signal \N__10517\ : std_logic;
signal \N__10514\ : std_logic;
signal \N__10513\ : std_logic;
signal \N__10510\ : std_logic;
signal \N__10507\ : std_logic;
signal \N__10504\ : std_logic;
signal \N__10501\ : std_logic;
signal \N__10500\ : std_logic;
signal \N__10497\ : std_logic;
signal \N__10496\ : std_logic;
signal \N__10493\ : std_logic;
signal \N__10490\ : std_logic;
signal \N__10489\ : std_logic;
signal \N__10486\ : std_logic;
signal \N__10483\ : std_logic;
signal \N__10482\ : std_logic;
signal \N__10477\ : std_logic;
signal \N__10476\ : std_logic;
signal \N__10475\ : std_logic;
signal \N__10472\ : std_logic;
signal \N__10467\ : std_logic;
signal \N__10464\ : std_logic;
signal \N__10461\ : std_logic;
signal \N__10458\ : std_logic;
signal \N__10455\ : std_logic;
signal \N__10452\ : std_logic;
signal \N__10449\ : std_logic;
signal \N__10446\ : std_logic;
signal \N__10439\ : std_logic;
signal \N__10436\ : std_logic;
signal \N__10431\ : std_logic;
signal \N__10428\ : std_logic;
signal \N__10423\ : std_logic;
signal \N__10418\ : std_logic;
signal \N__10415\ : std_logic;
signal \N__10412\ : std_logic;
signal \N__10409\ : std_logic;
signal \N__10406\ : std_logic;
signal \N__10403\ : std_logic;
signal \N__10400\ : std_logic;
signal \N__10399\ : std_logic;
signal \N__10396\ : std_logic;
signal \N__10395\ : std_logic;
signal \N__10394\ : std_logic;
signal \N__10391\ : std_logic;
signal \N__10384\ : std_logic;
signal \N__10379\ : std_logic;
signal \N__10378\ : std_logic;
signal \N__10377\ : std_logic;
signal \N__10376\ : std_logic;
signal \N__10373\ : std_logic;
signal \N__10366\ : std_logic;
signal \N__10361\ : std_logic;
signal \N__10358\ : std_logic;
signal \N__10357\ : std_logic;
signal \N__10356\ : std_logic;
signal \N__10355\ : std_logic;
signal \N__10352\ : std_logic;
signal \N__10349\ : std_logic;
signal \N__10344\ : std_logic;
signal \N__10341\ : std_logic;
signal \N__10334\ : std_logic;
signal \N__10331\ : std_logic;
signal \N__10328\ : std_logic;
signal \N__10327\ : std_logic;
signal \N__10326\ : std_logic;
signal \N__10325\ : std_logic;
signal \N__10322\ : std_logic;
signal \N__10319\ : std_logic;
signal \N__10314\ : std_logic;
signal \N__10311\ : std_logic;
signal \N__10304\ : std_logic;
signal \N__10301\ : std_logic;
signal \N__10298\ : std_logic;
signal \N__10295\ : std_logic;
signal \N__10294\ : std_logic;
signal \N__10293\ : std_logic;
signal \N__10290\ : std_logic;
signal \N__10287\ : std_logic;
signal \N__10284\ : std_logic;
signal \N__10277\ : std_logic;
signal \N__10276\ : std_logic;
signal \N__10275\ : std_logic;
signal \N__10272\ : std_logic;
signal \N__10269\ : std_logic;
signal \N__10264\ : std_logic;
signal \N__10259\ : std_logic;
signal \N__10256\ : std_logic;
signal \N__10253\ : std_logic;
signal \N__10250\ : std_logic;
signal \N__10247\ : std_logic;
signal \N__10246\ : std_logic;
signal \N__10243\ : std_logic;
signal \N__10240\ : std_logic;
signal \N__10237\ : std_logic;
signal \N__10234\ : std_logic;
signal \N__10231\ : std_logic;
signal \N__10228\ : std_logic;
signal \N__10225\ : std_logic;
signal \N__10220\ : std_logic;
signal \N__10219\ : std_logic;
signal \N__10216\ : std_logic;
signal \N__10213\ : std_logic;
signal \N__10210\ : std_logic;
signal \N__10207\ : std_logic;
signal \N__10204\ : std_logic;
signal \N__10201\ : std_logic;
signal \N__10198\ : std_logic;
signal \N__10195\ : std_logic;
signal \N__10192\ : std_logic;
signal \N__10189\ : std_logic;
signal \N__10186\ : std_logic;
signal \N__10183\ : std_logic;
signal \N__10180\ : std_logic;
signal \N__10177\ : std_logic;
signal \N__10174\ : std_logic;
signal \N__10171\ : std_logic;
signal \N__10168\ : std_logic;
signal \N__10165\ : std_logic;
signal \N__10162\ : std_logic;
signal \N__10159\ : std_logic;
signal \N__10156\ : std_logic;
signal \N__10153\ : std_logic;
signal \N__10150\ : std_logic;
signal \N__10147\ : std_logic;
signal \N__10144\ : std_logic;
signal \N__10141\ : std_logic;
signal \N__10138\ : std_logic;
signal \N__10135\ : std_logic;
signal \N__10132\ : std_logic;
signal \N__10129\ : std_logic;
signal \N__10126\ : std_logic;
signal \N__10123\ : std_logic;
signal \N__10120\ : std_logic;
signal \N__10117\ : std_logic;
signal \N__10114\ : std_logic;
signal \N__10111\ : std_logic;
signal \N__10108\ : std_logic;
signal \N__10105\ : std_logic;
signal \N__10102\ : std_logic;
signal \N__10099\ : std_logic;
signal \N__10096\ : std_logic;
signal \N__10093\ : std_logic;
signal \N__10090\ : std_logic;
signal \N__10087\ : std_logic;
signal \N__10084\ : std_logic;
signal \N__10081\ : std_logic;
signal \N__10078\ : std_logic;
signal \N__10075\ : std_logic;
signal \N__10072\ : std_logic;
signal \N__10069\ : std_logic;
signal \N__10066\ : std_logic;
signal \N__10063\ : std_logic;
signal \N__10060\ : std_logic;
signal \N__10057\ : std_logic;
signal \N__10054\ : std_logic;
signal \N__10051\ : std_logic;
signal \N__10048\ : std_logic;
signal \N__10045\ : std_logic;
signal \N__10042\ : std_logic;
signal \N__10039\ : std_logic;
signal \N__10036\ : std_logic;
signal \N__10033\ : std_logic;
signal \N__10030\ : std_logic;
signal \N__10027\ : std_logic;
signal \N__10024\ : std_logic;
signal \N__10021\ : std_logic;
signal \N__10018\ : std_logic;
signal \N__10015\ : std_logic;
signal \N__10012\ : std_logic;
signal \N__10009\ : std_logic;
signal \N__10006\ : std_logic;
signal \N__10001\ : std_logic;
signal \N__9998\ : std_logic;
signal \N__9995\ : std_logic;
signal \N__9992\ : std_logic;
signal \N__9989\ : std_logic;
signal \N__9988\ : std_logic;
signal \N__9985\ : std_logic;
signal \N__9984\ : std_logic;
signal \N__9981\ : std_logic;
signal \N__9978\ : std_logic;
signal \N__9975\ : std_logic;
signal \N__9968\ : std_logic;
signal \N__9965\ : std_logic;
signal \N__9964\ : std_logic;
signal \N__9961\ : std_logic;
signal \N__9960\ : std_logic;
signal \N__9957\ : std_logic;
signal \N__9954\ : std_logic;
signal \N__9951\ : std_logic;
signal \N__9944\ : std_logic;
signal \N__9941\ : std_logic;
signal \N__9938\ : std_logic;
signal \N__9937\ : std_logic;
signal \N__9936\ : std_logic;
signal \N__9933\ : std_logic;
signal \N__9930\ : std_logic;
signal \N__9927\ : std_logic;
signal \N__9920\ : std_logic;
signal \N__9917\ : std_logic;
signal \N__9916\ : std_logic;
signal \N__9913\ : std_logic;
signal \N__9910\ : std_logic;
signal \N__9905\ : std_logic;
signal \N__9902\ : std_logic;
signal \N__9899\ : std_logic;
signal \N__9896\ : std_logic;
signal \N__9895\ : std_logic;
signal \N__9894\ : std_logic;
signal \N__9893\ : std_logic;
signal \N__9888\ : std_logic;
signal \N__9885\ : std_logic;
signal \N__9882\ : std_logic;
signal \N__9879\ : std_logic;
signal \N__9872\ : std_logic;
signal \N__9869\ : std_logic;
signal \N__9866\ : std_logic;
signal \N__9865\ : std_logic;
signal \N__9862\ : std_logic;
signal \N__9861\ : std_logic;
signal \N__9860\ : std_logic;
signal \N__9855\ : std_logic;
signal \N__9852\ : std_logic;
signal \N__9849\ : std_logic;
signal \N__9846\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9838\ : std_logic;
signal \N__9835\ : std_logic;
signal \N__9832\ : std_logic;
signal \N__9829\ : std_logic;
signal \N__9824\ : std_logic;
signal \N__9823\ : std_logic;
signal \N__9822\ : std_logic;
signal \N__9819\ : std_logic;
signal \N__9818\ : std_logic;
signal \N__9815\ : std_logic;
signal \N__9812\ : std_logic;
signal \N__9809\ : std_logic;
signal \N__9806\ : std_logic;
signal \N__9803\ : std_logic;
signal \N__9800\ : std_logic;
signal \N__9793\ : std_logic;
signal \N__9790\ : std_logic;
signal \N__9785\ : std_logic;
signal \N__9782\ : std_logic;
signal \N__9779\ : std_logic;
signal \N__9778\ : std_logic;
signal \N__9775\ : std_logic;
signal \N__9772\ : std_logic;
signal \N__9767\ : std_logic;
signal \N__9764\ : std_logic;
signal \N__9761\ : std_logic;
signal \N__9758\ : std_logic;
signal \N__9755\ : std_logic;
signal \N__9754\ : std_logic;
signal \N__9751\ : std_logic;
signal \N__9748\ : std_logic;
signal \N__9743\ : std_logic;
signal \N__9740\ : std_logic;
signal \N__9739\ : std_logic;
signal \N__9736\ : std_logic;
signal \N__9733\ : std_logic;
signal \N__9728\ : std_logic;
signal \N__9725\ : std_logic;
signal \N__9722\ : std_logic;
signal \N__9719\ : std_logic;
signal \N__9716\ : std_logic;
signal \N__9715\ : std_logic;
signal \N__9714\ : std_logic;
signal \N__9711\ : std_logic;
signal \N__9708\ : std_logic;
signal \N__9705\ : std_logic;
signal \N__9698\ : std_logic;
signal \N__9697\ : std_logic;
signal \N__9696\ : std_logic;
signal \N__9693\ : std_logic;
signal \N__9690\ : std_logic;
signal \N__9687\ : std_logic;
signal \N__9680\ : std_logic;
signal \N__9677\ : std_logic;
signal \N__9674\ : std_logic;
signal \N__9671\ : std_logic;
signal \N__9668\ : std_logic;
signal \N__9665\ : std_logic;
signal \N__9662\ : std_logic;
signal \N__9659\ : std_logic;
signal \N__9656\ : std_logic;
signal \N__9653\ : std_logic;
signal \N__9650\ : std_logic;
signal \N__9647\ : std_logic;
signal \N__9644\ : std_logic;
signal \N__9641\ : std_logic;
signal \N__9638\ : std_logic;
signal \N__9635\ : std_logic;
signal \N__9632\ : std_logic;
signal \N__9631\ : std_logic;
signal \N__9630\ : std_logic;
signal \N__9627\ : std_logic;
signal \N__9624\ : std_logic;
signal \N__9621\ : std_logic;
signal \N__9618\ : std_logic;
signal \N__9613\ : std_logic;
signal \N__9610\ : std_logic;
signal \N__9607\ : std_logic;
signal \N__9602\ : std_logic;
signal \N__9599\ : std_logic;
signal \N__9596\ : std_logic;
signal \N__9593\ : std_logic;
signal \N__9590\ : std_logic;
signal \N__9587\ : std_logic;
signal \N__9584\ : std_logic;
signal \N__9581\ : std_logic;
signal \N__9578\ : std_logic;
signal \N__9575\ : std_logic;
signal \N__9572\ : std_logic;
signal \N__9569\ : std_logic;
signal \N__9566\ : std_logic;
signal \N__9563\ : std_logic;
signal \N__9560\ : std_logic;
signal \N__9557\ : std_logic;
signal \N__9554\ : std_logic;
signal \N__9551\ : std_logic;
signal \N__9548\ : std_logic;
signal \N__9545\ : std_logic;
signal \N__9542\ : std_logic;
signal \N__9539\ : std_logic;
signal \N__9536\ : std_logic;
signal \N__9533\ : std_logic;
signal \N__9530\ : std_logic;
signal \N__9527\ : std_logic;
signal \N__9524\ : std_logic;
signal \N__9523\ : std_logic;
signal \N__9520\ : std_logic;
signal \N__9517\ : std_logic;
signal \N__9516\ : std_logic;
signal \N__9515\ : std_logic;
signal \N__9514\ : std_logic;
signal \N__9513\ : std_logic;
signal \N__9512\ : std_logic;
signal \N__9509\ : std_logic;
signal \N__9506\ : std_logic;
signal \N__9503\ : std_logic;
signal \N__9502\ : std_logic;
signal \N__9499\ : std_logic;
signal \N__9498\ : std_logic;
signal \N__9497\ : std_logic;
signal \N__9496\ : std_logic;
signal \N__9495\ : std_logic;
signal \N__9492\ : std_logic;
signal \N__9489\ : std_logic;
signal \N__9486\ : std_logic;
signal \N__9485\ : std_logic;
signal \N__9484\ : std_logic;
signal \N__9477\ : std_logic;
signal \N__9474\ : std_logic;
signal \N__9471\ : std_logic;
signal \N__9468\ : std_logic;
signal \N__9465\ : std_logic;
signal \N__9462\ : std_logic;
signal \N__9459\ : std_logic;
signal \N__9456\ : std_logic;
signal \N__9451\ : std_logic;
signal \N__9448\ : std_logic;
signal \N__9445\ : std_logic;
signal \N__9442\ : std_logic;
signal \N__9435\ : std_logic;
signal \N__9428\ : std_logic;
signal \N__9421\ : std_logic;
signal \N__9418\ : std_logic;
signal \N__9415\ : std_logic;
signal \N__9412\ : std_logic;
signal \N__9409\ : std_logic;
signal \N__9406\ : std_logic;
signal \N__9403\ : std_logic;
signal \N__9392\ : std_logic;
signal \N__9389\ : std_logic;
signal \N__9386\ : std_logic;
signal \N__9383\ : std_logic;
signal \N__9380\ : std_logic;
signal \N__9377\ : std_logic;
signal \N__9374\ : std_logic;
signal \N__9371\ : std_logic;
signal \N__9368\ : std_logic;
signal \N__9365\ : std_logic;
signal \N__9362\ : std_logic;
signal \N__9359\ : std_logic;
signal \N__9356\ : std_logic;
signal \N__9353\ : std_logic;
signal \N__9350\ : std_logic;
signal \N__9347\ : std_logic;
signal \N__9344\ : std_logic;
signal \N__9341\ : std_logic;
signal \N__9338\ : std_logic;
signal \N__9335\ : std_logic;
signal \N__9332\ : std_logic;
signal \N__9329\ : std_logic;
signal \N__9326\ : std_logic;
signal \N__9323\ : std_logic;
signal \N__9320\ : std_logic;
signal \N__9317\ : std_logic;
signal \N__9314\ : std_logic;
signal \N__9311\ : std_logic;
signal \N__9308\ : std_logic;
signal \N__9305\ : std_logic;
signal \N__9302\ : std_logic;
signal \N__9299\ : std_logic;
signal \N__9296\ : std_logic;
signal \N__9293\ : std_logic;
signal \N__9290\ : std_logic;
signal \N__9287\ : std_logic;
signal \N__9284\ : std_logic;
signal \N__9281\ : std_logic;
signal \N__9278\ : std_logic;
signal \N__9275\ : std_logic;
signal \N__9272\ : std_logic;
signal \N__9269\ : std_logic;
signal \N__9266\ : std_logic;
signal \N__9263\ : std_logic;
signal \N__9260\ : std_logic;
signal \N__9257\ : std_logic;
signal \N__9254\ : std_logic;
signal \N__9251\ : std_logic;
signal \N__9248\ : std_logic;
signal \N__9245\ : std_logic;
signal \N__9242\ : std_logic;
signal \N__9239\ : std_logic;
signal \N__9236\ : std_logic;
signal \N__9233\ : std_logic;
signal \N__9230\ : std_logic;
signal \N__9227\ : std_logic;
signal \N__9224\ : std_logic;
signal \N__9221\ : std_logic;
signal \N__9218\ : std_logic;
signal \N__9215\ : std_logic;
signal \N__9212\ : std_logic;
signal \N__9209\ : std_logic;
signal \N__9206\ : std_logic;
signal \N__9203\ : std_logic;
signal \N__9200\ : std_logic;
signal \N__9197\ : std_logic;
signal \N__9194\ : std_logic;
signal \N__9191\ : std_logic;
signal \N__9188\ : std_logic;
signal \N__9185\ : std_logic;
signal \N__9182\ : std_logic;
signal \N__9179\ : std_logic;
signal \N__9176\ : std_logic;
signal \N__9173\ : std_logic;
signal \N__9170\ : std_logic;
signal \N__9167\ : std_logic;
signal \N__9164\ : std_logic;
signal \N__9161\ : std_logic;
signal \N__9158\ : std_logic;
signal \N__9155\ : std_logic;
signal \N__9152\ : std_logic;
signal \N__9149\ : std_logic;
signal \N__9146\ : std_logic;
signal \N__9143\ : std_logic;
signal \N__9140\ : std_logic;
signal \N__9137\ : std_logic;
signal \N__9134\ : std_logic;
signal \N__9131\ : std_logic;
signal \N__9128\ : std_logic;
signal \N__9125\ : std_logic;
signal \N__9122\ : std_logic;
signal \N__9119\ : std_logic;
signal \N__9116\ : std_logic;
signal \N__9113\ : std_logic;
signal \N__9110\ : std_logic;
signal \N__9107\ : std_logic;
signal \N__9104\ : std_logic;
signal \N__9101\ : std_logic;
signal \N__9098\ : std_logic;
signal \N__9097\ : std_logic;
signal \N__9094\ : std_logic;
signal \N__9091\ : std_logic;
signal \N__9086\ : std_logic;
signal \N__9083\ : std_logic;
signal \N__9080\ : std_logic;
signal \N__9077\ : std_logic;
signal \N__9074\ : std_logic;
signal \N__9071\ : std_logic;
signal \N__9070\ : std_logic;
signal \N__9069\ : std_logic;
signal \N__9068\ : std_logic;
signal \N__9065\ : std_logic;
signal \N__9062\ : std_logic;
signal \N__9059\ : std_logic;
signal \N__9058\ : std_logic;
signal \N__9057\ : std_logic;
signal \N__9054\ : std_logic;
signal \N__9051\ : std_logic;
signal \N__9048\ : std_logic;
signal \N__9045\ : std_logic;
signal \N__9042\ : std_logic;
signal \N__9039\ : std_logic;
signal \N__9038\ : std_logic;
signal \N__9035\ : std_logic;
signal \N__9032\ : std_logic;
signal \N__9027\ : std_logic;
signal \N__9024\ : std_logic;
signal \N__9021\ : std_logic;
signal \N__9018\ : std_logic;
signal \N__9015\ : std_logic;
signal \N__9010\ : std_logic;
signal \N__9007\ : std_logic;
signal \N__9002\ : std_logic;
signal \N__9001\ : std_logic;
signal \N__8992\ : std_logic;
signal \N__8989\ : std_logic;
signal \N__8984\ : std_logic;
signal \N__8981\ : std_logic;
signal \N__8978\ : std_logic;
signal \N__8975\ : std_logic;
signal \N__8972\ : std_logic;
signal \N__8969\ : std_logic;
signal \N__8968\ : std_logic;
signal \N__8965\ : std_logic;
signal \N__8962\ : std_logic;
signal \N__8959\ : std_logic;
signal \N__8956\ : std_logic;
signal \N__8953\ : std_logic;
signal \N__8950\ : std_logic;
signal \N__8947\ : std_logic;
signal \N__8944\ : std_logic;
signal \N__8941\ : std_logic;
signal \N__8938\ : std_logic;
signal \N__8935\ : std_logic;
signal \N__8932\ : std_logic;
signal \N__8929\ : std_logic;
signal \N__8926\ : std_logic;
signal \N__8923\ : std_logic;
signal \N__8920\ : std_logic;
signal \N__8917\ : std_logic;
signal \N__8914\ : std_logic;
signal \N__8911\ : std_logic;
signal \N__8908\ : std_logic;
signal \N__8905\ : std_logic;
signal \N__8902\ : std_logic;
signal \N__8899\ : std_logic;
signal \N__8896\ : std_logic;
signal \N__8893\ : std_logic;
signal \N__8890\ : std_logic;
signal \N__8887\ : std_logic;
signal \N__8884\ : std_logic;
signal \N__8881\ : std_logic;
signal \N__8878\ : std_logic;
signal \N__8875\ : std_logic;
signal \N__8872\ : std_logic;
signal \N__8869\ : std_logic;
signal \N__8866\ : std_logic;
signal \N__8863\ : std_logic;
signal \N__8860\ : std_logic;
signal \N__8857\ : std_logic;
signal \N__8854\ : std_logic;
signal \N__8851\ : std_logic;
signal \N__8848\ : std_logic;
signal \N__8845\ : std_logic;
signal \N__8842\ : std_logic;
signal \N__8839\ : std_logic;
signal \N__8836\ : std_logic;
signal \N__8833\ : std_logic;
signal \N__8830\ : std_logic;
signal \N__8827\ : std_logic;
signal \N__8824\ : std_logic;
signal \N__8821\ : std_logic;
signal \N__8818\ : std_logic;
signal \N__8815\ : std_logic;
signal \N__8812\ : std_logic;
signal \N__8809\ : std_logic;
signal \N__8806\ : std_logic;
signal \N__8803\ : std_logic;
signal \N__8800\ : std_logic;
signal \N__8797\ : std_logic;
signal \N__8794\ : std_logic;
signal \N__8791\ : std_logic;
signal \N__8788\ : std_logic;
signal \N__8785\ : std_logic;
signal \N__8782\ : std_logic;
signal \N__8779\ : std_logic;
signal \N__8776\ : std_logic;
signal \N__8773\ : std_logic;
signal \N__8770\ : std_logic;
signal \N__8767\ : std_logic;
signal \N__8764\ : std_logic;
signal \N__8761\ : std_logic;
signal \N__8756\ : std_logic;
signal \N__8753\ : std_logic;
signal \N__8750\ : std_logic;
signal \N__8747\ : std_logic;
signal \N__8744\ : std_logic;
signal \N__8741\ : std_logic;
signal \N__8738\ : std_logic;
signal \N__8735\ : std_logic;
signal \N__8732\ : std_logic;
signal \N__8729\ : std_logic;
signal \N__8726\ : std_logic;
signal \N__8723\ : std_logic;
signal \N__8720\ : std_logic;
signal \N__8717\ : std_logic;
signal \N__8714\ : std_logic;
signal \N__8711\ : std_logic;
signal \N__8708\ : std_logic;
signal \N__8705\ : std_logic;
signal \N__8702\ : std_logic;
signal \N__8699\ : std_logic;
signal \N__8696\ : std_logic;
signal \N__8693\ : std_logic;
signal \N__8690\ : std_logic;
signal \N__8687\ : std_logic;
signal \N__8684\ : std_logic;
signal \N__8681\ : std_logic;
signal \N__8678\ : std_logic;
signal \N__8675\ : std_logic;
signal \N__8672\ : std_logic;
signal \N__8669\ : std_logic;
signal \N__8666\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8660\ : std_logic;
signal \N__8657\ : std_logic;
signal \N__8654\ : std_logic;
signal \N__8651\ : std_logic;
signal \N__8648\ : std_logic;
signal \N__8645\ : std_logic;
signal \N__8642\ : std_logic;
signal \N__8639\ : std_logic;
signal \N__8636\ : std_logic;
signal \N__8633\ : std_logic;
signal \N__8630\ : std_logic;
signal \N__8627\ : std_logic;
signal \N__8624\ : std_logic;
signal \N__8621\ : std_logic;
signal \N__8618\ : std_logic;
signal \N__8615\ : std_logic;
signal \N__8612\ : std_logic;
signal \N__8609\ : std_logic;
signal \N__8606\ : std_logic;
signal \N__8603\ : std_logic;
signal \N__8600\ : std_logic;
signal \N__8597\ : std_logic;
signal \N__8594\ : std_logic;
signal \N__8591\ : std_logic;
signal \N__8588\ : std_logic;
signal \N__8585\ : std_logic;
signal \N__8582\ : std_logic;
signal \N__8579\ : std_logic;
signal \N__8576\ : std_logic;
signal \N__8573\ : std_logic;
signal \N__8570\ : std_logic;
signal \N__8567\ : std_logic;
signal \N__8564\ : std_logic;
signal \N__8561\ : std_logic;
signal \N__8558\ : std_logic;
signal \N__8555\ : std_logic;
signal \N__8552\ : std_logic;
signal \N__8549\ : std_logic;
signal \N__8546\ : std_logic;
signal \N__8543\ : std_logic;
signal \N__8540\ : std_logic;
signal \N__8537\ : std_logic;
signal \N__8534\ : std_logic;
signal \N__8531\ : std_logic;
signal \N__8528\ : std_logic;
signal \N__8525\ : std_logic;
signal \N__8522\ : std_logic;
signal \N__8519\ : std_logic;
signal \N__8516\ : std_logic;
signal \N__8513\ : std_logic;
signal \N__8510\ : std_logic;
signal \N__8507\ : std_logic;
signal \N__8504\ : std_logic;
signal \N__8501\ : std_logic;
signal \N__8498\ : std_logic;
signal \N__8495\ : std_logic;
signal \N__8492\ : std_logic;
signal \N__8489\ : std_logic;
signal \N__8486\ : std_logic;
signal \N__8483\ : std_logic;
signal \N__8480\ : std_logic;
signal \N__8477\ : std_logic;
signal \N__8474\ : std_logic;
signal \N__8471\ : std_logic;
signal \N__8468\ : std_logic;
signal \N__8465\ : std_logic;
signal \N__8462\ : std_logic;
signal \N__8459\ : std_logic;
signal \N__8456\ : std_logic;
signal \N__8453\ : std_logic;
signal \N__8450\ : std_logic;
signal \N__8447\ : std_logic;
signal \N__8444\ : std_logic;
signal \N__8441\ : std_logic;
signal \N__8438\ : std_logic;
signal \N__8435\ : std_logic;
signal \N__8432\ : std_logic;
signal \N__8429\ : std_logic;
signal \N__8426\ : std_logic;
signal \N__8423\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8414\ : std_logic;
signal \N__8411\ : std_logic;
signal \N__8408\ : std_logic;
signal \N__8405\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_37\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_36\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_31\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_32\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_33\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_38\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_35\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_34\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_9\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_8\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_22\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_21\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_20\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_19\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_18\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_15\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_23\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_17\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_16\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_14\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_39\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_41\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_40\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_13\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_12\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_7\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_6\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_11\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_10\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_73\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_72\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_63\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_71\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_70\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_66\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_67\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_65\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_64\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_69\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_68\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_24\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_25\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_43\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_42\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_44\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_45\ : std_logic;
signal \DEBUG_c_5_c\ : std_logic;
signal \RX_DATA_3\ : std_logic;
signal \tvp_video_buffer.BUFFER_0_5\ : std_logic;
signal \tvp_video_buffer.BUFFER_1_5\ : std_logic;
signal n27 : std_logic;
signal \line_buffer.n603\ : std_logic;
signal \line_buffer.n595\ : std_logic;
signal \line_buffer.n602\ : std_logic;
signal \line_buffer.n594\ : std_logic;
signal \TVP_VIDEO_c_2\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_74\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_75\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_78\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_79\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_77\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_76\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_62\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_61\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_80\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_82\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_81\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_83\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_85\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_84\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_26\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_27\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_28\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_30\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_29\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_47\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_46\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_49\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_48\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_53\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_52\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_51\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_50\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_60\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_59\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_58\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_54\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_55\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_57\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_56\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_86\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_96\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_99\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_98\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_97\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_95\ : std_logic;
signal \transmit_module.n3683\ : std_logic;
signal \transmit_module.video_signal_controller.n6_cascade_\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_11\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_12\ : std_logic;
signal \bfn_11_17_0_\ : std_logic;
signal \transmit_module.video_signal_controller.n3183\ : std_logic;
signal \transmit_module.video_signal_controller.n3184\ : std_logic;
signal \transmit_module.video_signal_controller.n3185\ : std_logic;
signal \transmit_module.video_signal_controller.n3186\ : std_logic;
signal \transmit_module.video_signal_controller.n3187\ : std_logic;
signal \transmit_module.video_signal_controller.n3188\ : std_logic;
signal \transmit_module.video_signal_controller.n3189\ : std_logic;
signal \transmit_module.video_signal_controller.n3190\ : std_logic;
signal \bfn_11_18_0_\ : std_logic;
signal \transmit_module.video_signal_controller.n3191\ : std_logic;
signal \transmit_module.video_signal_controller.n3192\ : std_logic;
signal \transmit_module.video_signal_controller.n3193\ : std_logic;
signal \tvp_video_buffer.BUFFER_0_2\ : std_logic;
signal \TVP_VIDEO_c_3\ : std_logic;
signal \tvp_video_buffer.BUFFER_0_3\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_15\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_14\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_94\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_93\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_92\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_87\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_89\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_88\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_91\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_90\ : std_logic;
signal \transmit_module.n2209\ : std_logic;
signal \bfn_12_14_0_\ : std_logic;
signal \transmit_module.video_signal_controller.n3194\ : std_logic;
signal \transmit_module.video_signal_controller.n3195\ : std_logic;
signal \transmit_module.video_signal_controller.n3196\ : std_logic;
signal \transmit_module.video_signal_controller.n3197\ : std_logic;
signal \transmit_module.video_signal_controller.n3198\ : std_logic;
signal \transmit_module.video_signal_controller.n3199\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_7\ : std_logic;
signal \transmit_module.video_signal_controller.n3200\ : std_logic;
signal \transmit_module.video_signal_controller.n3201\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_8\ : std_logic;
signal \bfn_12_15_0_\ : std_logic;
signal \transmit_module.video_signal_controller.n3202\ : std_logic;
signal \transmit_module.video_signal_controller.n3203\ : std_logic;
signal \transmit_module.video_signal_controller.n3204\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_11\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_10\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_5\ : std_logic;
signal \transmit_module.video_signal_controller.n3485_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_6\ : std_logic;
signal \transmit_module.video_signal_controller.n3676\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_9\ : std_logic;
signal \transmit_module.video_signal_controller.n3464_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.n3378\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_5\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_3\ : std_logic;
signal \transmit_module.video_signal_controller.n6_adj_622\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_4\ : std_logic;
signal \transmit_module.video_signal_controller.n2019\ : std_logic;
signal \transmit_module.video_signal_controller.n2050\ : std_logic;
signal \transmit_module.video_signal_controller.n2050_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.n2398\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_3\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_4\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_6\ : std_logic;
signal \transmit_module.video_signal_controller.n3482_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_5\ : std_logic;
signal \transmit_module.video_signal_controller.n55\ : std_logic;
signal \transmit_module.video_signal_controller.n3478_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_7\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_0\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_13\ : std_logic;
signal \transmit_module.n2073\ : std_logic;
signal n20 : std_logic;
signal \tvp_video_buffer.BUFFER_1_2\ : std_logic;
signal \RX_DATA_0\ : std_logic;
signal \TVP_VIDEO_c_4\ : std_logic;
signal \tvp_video_buffer.BUFFER_0_4\ : std_logic;
signal \TVP_VIDEO_c_8\ : std_logic;
signal \tvp_video_buffer.BUFFER_1_3\ : std_logic;
signal \RX_DATA_1\ : std_logic;
signal \tvp_video_buffer.BUFFER_1_4\ : std_logic;
signal \RX_DATA_2\ : std_logic;
signal \tvp_video_buffer.BUFFER_0_8\ : std_logic;
signal \tvp_video_buffer.BUFFER_1_8\ : std_logic;
signal \bfn_13_9_0_\ : std_logic;
signal \receive_module.rx_counter.n3210\ : std_logic;
signal \receive_module.rx_counter.n3211\ : std_logic;
signal \receive_module.rx_counter.n3212\ : std_logic;
signal \receive_module.rx_counter.n3213\ : std_logic;
signal \receive_module.rx_counter.n3214\ : std_logic;
signal \receive_module.rx_counter.n3215\ : std_logic;
signal \receive_module.rx_counter.n3216\ : std_logic;
signal \receive_module.rx_counter.n3217\ : std_logic;
signal \bfn_13_10_0_\ : std_logic;
signal \receive_module.rx_counter.n3218\ : std_logic;
signal \bfn_13_11_0_\ : std_logic;
signal \receive_module.rx_counter.n3175\ : std_logic;
signal \receive_module.rx_counter.n3176\ : std_logic;
signal \receive_module.rx_counter.n3177\ : std_logic;
signal \receive_module.rx_counter.n3178\ : std_logic;
signal \receive_module.rx_counter.n3179\ : std_logic;
signal \receive_module.rx_counter.n3180\ : std_logic;
signal \receive_module.rx_counter.n3181\ : std_logic;
signal \receive_module.rx_counter.n3182\ : std_logic;
signal \bfn_13_12_0_\ : std_logic;
signal \receive_module.rx_counter.n10\ : std_logic;
signal \receive_module.rx_counter.n14_cascade_\ : std_logic;
signal \line_buffer.n539\ : std_logic;
signal \line_buffer.n531\ : std_logic;
signal \transmit_module.old_VGA_HS\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_7\ : std_logic;
signal \transmit_module.video_signal_controller.n7\ : std_logic;
signal \ADV_HSYNC_c\ : std_logic;
signal \transmit_module.n141_cascade_\ : std_logic;
signal n22 : std_logic;
signal \transmit_module.VGA_VISIBLE_Y\ : std_logic;
signal \transmit_module.n140\ : std_logic;
signal \transmit_module.n140_cascade_\ : std_logic;
signal \transmit_module.n109\ : std_logic;
signal n21 : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_1\ : std_logic;
signal \transmit_module.video_signal_controller.n3520\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_0\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_Y_2\ : std_logic;
signal \transmit_module.video_signal_controller.n2958\ : std_logic;
signal \transmit_module.video_signal_controller.n2975\ : std_logic;
signal \transmit_module.n142\ : std_logic;
signal \transmit_module.n142_cascade_\ : std_logic;
signal \transmit_module.n111\ : std_logic;
signal n23 : std_logic;
signal \transmit_module.video_signal_controller.n3366\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_8\ : std_logic;
signal \transmit_module.video_signal_controller.n2017\ : std_logic;
signal \transmit_module.video_signal_controller.n3007_cascade_\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_VISIBLE_N_588\ : std_logic;
signal \transmit_module.n143\ : std_logic;
signal \transmit_module.n143_cascade_\ : std_logic;
signal n24 : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_10\ : std_logic;
signal \transmit_module.video_signal_controller.n3007\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_2\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_1\ : std_logic;
signal \transmit_module.video_signal_controller.n3679\ : std_logic;
signal \transmit_module.n108\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_9\ : std_logic;
signal \transmit_module.video_signal_controller.n6_adj_623\ : std_logic;
signal \transmit_module.n139\ : std_logic;
signal \transmit_module.n138_cascade_\ : std_logic;
signal n19 : std_logic;
signal \line_buffer.n3531\ : std_logic;
signal \line_buffer.n3530\ : std_logic;
signal \line_buffer.n3620\ : std_logic;
signal \line_buffer.n571\ : std_logic;
signal \line_buffer.n563\ : std_logic;
signal \line_buffer.n3534\ : std_logic;
signal \TX_DATA_7\ : std_logic;
signal \ADV_B_c\ : std_logic;
signal \line_buffer.n474\ : std_logic;
signal \line_buffer.n466\ : std_logic;
signal \line_buffer.n3533\ : std_logic;
signal \line_buffer.n542\ : std_logic;
signal \receive_module.rx_counter.X_1\ : std_logic;
signal \receive_module.rx_counter.X_0\ : std_logic;
signal \receive_module.rx_counter.X_2\ : std_logic;
signal \receive_module.rx_counter.n3225_cascade_\ : std_logic;
signal \receive_module.rx_counter.n3458_cascade_\ : std_logic;
signal \receive_module.rx_counter.X_4\ : std_logic;
signal \receive_module.rx_counter.X_6\ : std_logic;
signal \receive_module.rx_counter.n3\ : std_logic;
signal \receive_module.rx_counter.X_3\ : std_logic;
signal \receive_module.rx_counter.X_5\ : std_logic;
signal \receive_module.rx_counter.X_7\ : std_logic;
signal \receive_module.rx_counter.n6\ : std_logic;
signal \receive_module.rx_counter.n7_cascade_\ : std_logic;
signal \receive_module.rx_counter.n3225\ : std_logic;
signal \receive_module.rx_counter.old_HS\ : std_logic;
signal \receive_module.rx_counter.n2081\ : std_logic;
signal \line_buffer.n573\ : std_logic;
signal \receive_module.rx_counter.n3429\ : std_logic;
signal \receive_module.rx_counter.X_8\ : std_logic;
signal \receive_module.rx_counter.X_9\ : std_logic;
signal \receive_module.rx_counter.n39\ : std_logic;
signal \receive_module.rx_counter.Y_6\ : std_logic;
signal \receive_module.rx_counter.Y_5\ : std_logic;
signal \receive_module.rx_counter.n5_cascade_\ : std_logic;
signal \receive_module.rx_counter.Y_7\ : std_logic;
signal \receive_module.rx_counter.n3455_cascade_\ : std_logic;
signal \receive_module.rx_counter.n3680\ : std_logic;
signal \receive_module.rx_counter.Y_8\ : std_logic;
signal \receive_module.rx_counter.n3481\ : std_logic;
signal \receive_module.rx_counter.n4_adj_612_cascade_\ : std_logic;
signal \receive_module.rx_counter.n54\ : std_logic;
signal \receive_module.rx_counter.Y_1\ : std_logic;
signal \receive_module.rx_counter.Y_0\ : std_logic;
signal \receive_module.rx_counter.Y_2\ : std_logic;
signal \receive_module.rx_counter.n3453\ : std_logic;
signal \receive_module.rx_counter.Y_3\ : std_logic;
signal \receive_module.rx_counter.Y_4\ : std_logic;
signal \receive_module.rx_counter.n4\ : std_logic;
signal \RX_TX_SYNC\ : std_logic;
signal \line_buffer.n477\ : std_logic;
signal \line_buffer.n541\ : std_logic;
signal \line_buffer.n605\ : std_logic;
signal \line_buffer.n568\ : std_logic;
signal \line_buffer.n560\ : std_logic;
signal \sync_buffer.BUFFER_0_0\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_6\ : std_logic;
signal \bfn_14_15_0_\ : std_logic;
signal \transmit_module.n131\ : std_logic;
signal \transmit_module.n3162\ : std_logic;
signal \transmit_module.n3163\ : std_logic;
signal \transmit_module.n3164\ : std_logic;
signal \transmit_module.n128\ : std_logic;
signal \transmit_module.n3165\ : std_logic;
signal \transmit_module.TX_ADDR_5\ : std_logic;
signal \transmit_module.n127\ : std_logic;
signal \transmit_module.n3166\ : std_logic;
signal \transmit_module.n126\ : std_logic;
signal \transmit_module.n3167\ : std_logic;
signal \transmit_module.TX_ADDR_7\ : std_logic;
signal \transmit_module.n125\ : std_logic;
signal \transmit_module.n3168\ : std_logic;
signal \transmit_module.n3169\ : std_logic;
signal \transmit_module.n124\ : std_logic;
signal \bfn_14_16_0_\ : std_logic;
signal \transmit_module.n123\ : std_logic;
signal \transmit_module.n3170\ : std_logic;
signal \transmit_module.n3171\ : std_logic;
signal \transmit_module.n121\ : std_logic;
signal \transmit_module.n3172\ : std_logic;
signal \transmit_module.n120\ : std_logic;
signal \transmit_module.n3173\ : std_logic;
signal \transmit_module.n3174\ : std_logic;
signal \transmit_module.n119\ : std_logic;
signal \transmit_module.n112\ : std_logic;
signal \transmit_module.n146\ : std_logic;
signal \sync_buffer.BUFFER_1_0\ : std_logic;
signal \RX_TX_SYNC_BUFF\ : std_logic;
signal \transmit_module.n122\ : std_logic;
signal \transmit_module.n137_cascade_\ : std_logic;
signal \transmit_module.n138\ : std_logic;
signal \transmit_module.video_signal_controller.n3382\ : std_logic;
signal \transmit_module.video_signal_controller.n3017\ : std_logic;
signal \transmit_module.video_signal_controller.VGA_X_11\ : std_logic;
signal \transmit_module.video_signal_controller.n7_adj_624\ : std_logic;
signal \transmit_module.n132\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_9\ : std_logic;
signal \transmit_module.TX_ADDR_9\ : std_logic;
signal \transmit_module.n107\ : std_logic;
signal \transmit_module.n115\ : std_logic;
signal \transmit_module.n116\ : std_logic;
signal \transmit_module.n116_cascade_\ : std_logic;
signal \transmit_module.n147\ : std_logic;
signal n28 : std_logic;
signal \transmit_module.n106\ : std_logic;
signal \transmit_module.n137\ : std_logic;
signal n18 : std_logic;
signal \transmit_module.TX_ADDR_10\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_10\ : std_logic;
signal \transmit_module.TX_ADDR_8\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_8\ : std_logic;
signal \transmit_module.TX_ADDR_1\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_1\ : std_logic;
signal \transmit_module.TX_ADDR_0\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_0\ : std_logic;
signal \DEBUG_c_1_c\ : std_logic;
signal \DEBUG_c_6_c\ : std_logic;
signal \tvp_vs_buffer.BUFFER_0_0\ : std_logic;
signal \tvp_video_buffer.BUFFER_0_6\ : std_logic;
signal \TVP_HSYNC_buff\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_10\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_9\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_11\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_13\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_12\ : std_logic;
signal \bfn_15_11_0_\ : std_logic;
signal \receive_module.n3149\ : std_logic;
signal \receive_module.n3150\ : std_logic;
signal \receive_module.n3151\ : std_logic;
signal \receive_module.n3152\ : std_logic;
signal \receive_module.n3153\ : std_logic;
signal \receive_module.n3154\ : std_logic;
signal \receive_module.n3155\ : std_logic;
signal \receive_module.n3156\ : std_logic;
signal \bfn_15_12_0_\ : std_logic;
signal \receive_module.n3157\ : std_logic;
signal \receive_module.n3158\ : std_logic;
signal \receive_module.n3159\ : std_logic;
signal \receive_module.n3160\ : std_logic;
signal \receive_module.n3161\ : std_logic;
signal \line_buffer.n606\ : std_logic;
signal \line_buffer.n476\ : std_logic;
signal \receive_module.n3674\ : std_logic;
signal \RX_ADDR_11\ : std_logic;
signal \RX_ADDR_12\ : std_logic;
signal \RX_ADDR_13\ : std_logic;
signal \line_buffer.n574\ : std_logic;
signal \tvp_vs_buffer.BUFFER_1_0\ : std_logic;
signal \tvp_vs_buffer.BUFFER_2_0\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_0\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_1\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_8\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_2\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_3\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_7\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_4\ : std_logic;
signal \transmit_module.n129\ : std_logic;
signal \transmit_module.n110\ : std_logic;
signal \transmit_module.n141\ : std_logic;
signal \transmit_module.TX_ADDR_6\ : std_logic;
signal \transmit_module.VGA_VISIBLE\ : std_logic;
signal \transmit_module.n130\ : std_logic;
signal \transmit_module.n145_cascade_\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_2\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_5\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_4\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_3\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_1\ : std_logic;
signal \receive_module.n136\ : std_logic;
signal \RX_ADDR_1\ : std_logic;
signal \receive_module.n135\ : std_logic;
signal \RX_ADDR_2\ : std_logic;
signal \receive_module.n133\ : std_logic;
signal \RX_ADDR_4\ : std_logic;
signal \receive_module.n132\ : std_logic;
signal \RX_ADDR_5\ : std_logic;
signal \receive_module.n131\ : std_logic;
signal \RX_ADDR_6\ : std_logic;
signal \receive_module.n130\ : std_logic;
signal \RX_ADDR_7\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_3\ : std_logic;
signal \transmit_module.TX_ADDR_3\ : std_logic;
signal \receive_module.n128\ : std_logic;
signal \RX_ADDR_9\ : std_logic;
signal \GB_BUFFER_DEBUG_c_3_c_THRU_CO\ : std_logic;
signal n1821 : std_logic;
signal \receive_module.n129\ : std_logic;
signal \RX_ADDR_8\ : std_logic;
signal \receive_module.n137\ : std_logic;
signal \RX_ADDR_0\ : std_logic;
signal \receive_module.n134\ : std_logic;
signal \RX_ADDR_3\ : std_logic;
signal \receive_module.n127\ : std_logic;
signal \RX_ADDR_10\ : std_logic;
signal \receive_module.n3677\ : std_logic;
signal \LED_c\ : std_logic;
signal \PULSE_1HZ\ : std_logic;
signal \receive_module.rx_counter.old_VS\ : std_logic;
signal \receive_module.rx_counter.n3522_cascade_\ : std_logic;
signal \receive_module.rx_counter.n7_adj_619\ : std_logic;
signal \receive_module.rx_counter.n11\ : std_logic;
signal \receive_module.rx_counter.FRAME_COUNTER_0\ : std_logic;
signal \bfn_16_10_0_\ : std_logic;
signal \receive_module.rx_counter.FRAME_COUNTER_1\ : std_logic;
signal \receive_module.rx_counter.n3205\ : std_logic;
signal \receive_module.rx_counter.FRAME_COUNTER_2\ : std_logic;
signal \receive_module.rx_counter.n3206\ : std_logic;
signal \receive_module.rx_counter.FRAME_COUNTER_3\ : std_logic;
signal \receive_module.rx_counter.n3207\ : std_logic;
signal \receive_module.rx_counter.FRAME_COUNTER_4\ : std_logic;
signal \receive_module.rx_counter.n3208\ : std_logic;
signal \receive_module.rx_counter.n3209\ : std_logic;
signal \receive_module.rx_counter.FRAME_COUNTER_5\ : std_logic;
signal \receive_module.rx_counter.n3675\ : std_logic;
signal \receive_module.rx_counter.n2550\ : std_logic;
signal \tvp_video_buffer.BUFFER_1_6\ : std_logic;
signal \RX_DATA_6\ : std_logic;
signal \RX_DATA_4\ : std_logic;
signal \receive_module.sync_wd.n6_cascade_\ : std_logic;
signal \receive_module.sync_wd.n4_cascade_\ : std_logic;
signal \TVP_VSYNC_buff\ : std_logic;
signal \DEBUG_c_0\ : std_logic;
signal \DEBUG_c_4\ : std_logic;
signal \receive_module.sync_wd.old_visible\ : std_logic;
signal \RX_DATA_7\ : std_logic;
signal \line_buffer.n569\ : std_logic;
signal \line_buffer.n561\ : std_logic;
signal \line_buffer.n567\ : std_logic;
signal \line_buffer.n559\ : std_logic;
signal \transmit_module.TX_ADDR_4\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_4\ : std_logic;
signal \transmit_module.n2313\ : std_logic;
signal \transmit_module.ADDR_Y_COMPONENT_2\ : std_logic;
signal \transmit_module.Y_DELTA_PATTERN_0\ : std_logic;
signal \transmit_module.TX_ADDR_2\ : std_logic;
signal \transmit_module.n114\ : std_logic;
signal \transmit_module.n145\ : std_logic;
signal n26 : std_logic;
signal \line_buffer.n535\ : std_logic;
signal \line_buffer.n527\ : std_logic;
signal \transmit_module.n3678\ : std_logic;
signal \ADV_VSYNC_c\ : std_logic;
signal \transmit_module.n113\ : std_logic;
signal \transmit_module.n144\ : std_logic;
signal n25 : std_logic;
signal n1818 : std_logic;
signal \line_buffer.n470\ : std_logic;
signal \line_buffer.n462\ : std_logic;
signal \line_buffer.n3590\ : std_logic;
signal \line_buffer.n3593_cascade_\ : std_logic;
signal \line_buffer.n3629\ : std_logic;
signal \TX_DATA_3\ : std_logic;
signal \line_buffer.n471\ : std_logic;
signal \line_buffer.n463\ : std_logic;
signal \line_buffer.n3552\ : std_logic;
signal \line_buffer.n3551_cascade_\ : std_logic;
signal \line_buffer.n600\ : std_logic;
signal \line_buffer.n592\ : std_logic;
signal \TX_DATA_4\ : std_logic;
signal n1817 : std_logic;
signal \TX_DATA_1\ : std_logic;
signal n1820 : std_logic;
signal \tvp_hs_buffer.BUFFER_1_0\ : std_logic;
signal \line_buffer.n536\ : std_logic;
signal \line_buffer.n528\ : std_logic;
signal \line_buffer.n534\ : std_logic;
signal \line_buffer.n526\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_6\ : std_logic;
signal \transmit_module.X_DELTA_PATTERN_5\ : std_logic;
signal \transmit_module.n2087\ : std_logic;
signal \transmit_module.n3682\ : std_logic;
signal \line_buffer.n533\ : std_logic;
signal \line_buffer.n525\ : std_logic;
signal \line_buffer.n3653\ : std_logic;
signal \line_buffer.n468\ : std_logic;
signal \line_buffer.n460\ : std_logic;
signal \line_buffer.n3635\ : std_logic;
signal \line_buffer.n566\ : std_logic;
signal \line_buffer.n558\ : std_logic;
signal \line_buffer.n557\ : std_logic;
signal \line_buffer.n565\ : std_logic;
signal \line_buffer.n3632\ : std_logic;
signal \line_buffer.n3572\ : std_logic;
signal \line_buffer.n3602_cascade_\ : std_logic;
signal \line_buffer.n3570\ : std_logic;
signal \line_buffer.n472\ : std_logic;
signal \line_buffer.n464\ : std_logic;
signal \line_buffer.n3656\ : std_logic;
signal \line_buffer.n599\ : std_logic;
signal \line_buffer.n591\ : std_logic;
signal \line_buffer.n3626\ : std_logic;
signal \TX_DATA_2\ : std_logic;
signal n1819 : std_logic;
signal \line_buffer.n3537\ : std_logic;
signal \line_buffer.n3536\ : std_logic;
signal \line_buffer.n3614\ : std_logic;
signal \line_buffer.n469\ : std_logic;
signal \line_buffer.n461\ : std_logic;
signal \line_buffer.n3569\ : std_logic;
signal \DEBUG_c_2_c\ : std_logic;
signal \tvp_hs_buffer.BUFFER_0_0\ : std_logic;
signal \line_buffer.n598\ : std_logic;
signal \line_buffer.n590\ : std_logic;
signal \line_buffer.n3573\ : std_logic;
signal \line_buffer.n3659\ : std_logic;
signal \line_buffer.n564\ : std_logic;
signal \line_buffer.n556\ : std_logic;
signal \line_buffer.n467\ : std_logic;
signal \line_buffer.n459\ : std_logic;
signal \line_buffer.n3638\ : std_logic;
signal \line_buffer.n3641\ : std_logic;
signal \TX_DATA_0\ : std_logic;
signal \line_buffer.n532\ : std_logic;
signal \line_buffer.n524\ : std_logic;
signal \line_buffer.n3647\ : std_logic;
signal \TX_DATA_5\ : std_logic;
signal n1816 : std_logic;
signal \line_buffer.n537\ : std_logic;
signal \line_buffer.n529\ : std_logic;
signal \line_buffer.n3599\ : std_logic;
signal \line_buffer.n597\ : std_logic;
signal \line_buffer.n589\ : std_logic;
signal \line_buffer.n3650\ : std_logic;
signal \line_buffer.n570\ : std_logic;
signal \line_buffer.n562\ : std_logic;
signal \line_buffer.n3543\ : std_logic;
signal \TX_ADDR_13\ : std_logic;
signal \line_buffer.n3608_cascade_\ : std_logic;
signal \line_buffer.n3576\ : std_logic;
signal \TX_DATA_6\ : std_logic;
signal n1815 : std_logic;
signal \ADV_CLK_c\ : std_logic;
signal \transmit_module.n2388\ : std_logic;
signal \line_buffer.n596\ : std_logic;
signal \line_buffer.n588\ : std_logic;
signal \line_buffer.n3644\ : std_logic;
signal \line_buffer.n473\ : std_logic;
signal \line_buffer.n465\ : std_logic;
signal \line_buffer.n3575\ : std_logic;
signal \tvp_video_buffer.BUFFER_1_9\ : std_logic;
signal \RX_DATA_5\ : std_logic;
signal \line_buffer.n601\ : std_logic;
signal \TX_ADDR_12\ : std_logic;
signal \line_buffer.n593\ : std_logic;
signal \line_buffer.n3596\ : std_logic;
signal \DEBUG_c_7_c\ : std_logic;
signal \tvp_video_buffer.BUFFER_0_7\ : std_logic;
signal \tvp_video_buffer.BUFFER_1_7\ : std_logic;
signal \TX_ADDR_11\ : std_logic;
signal \line_buffer.n538\ : std_logic;
signal \line_buffer.n530\ : std_logic;
signal \line_buffer.n3542\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \TVP_VIDEO_c_9\ : std_logic;
signal \tvp_video_buffer.BUFFER_0_9\ : std_logic;
signal \DEBUG_c_3_c\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \TVP_CLK_wire\ : std_logic;
signal \ADV_CLK_wire\ : std_logic;
signal \TVP_HSYNC_wire\ : std_logic;
signal \TVP_VIDEO_wire\ : std_logic_vector(9 downto 0);
signal \ADV_G_wire\ : std_logic_vector(7 downto 0);
signal \ADV_R_wire\ : std_logic_vector(7 downto 0);
signal \ADV_B_wire\ : std_logic_vector(7 downto 0);
signal \ADV_SYNC_N_wire\ : std_logic;
signal \ADV_BLANK_N_wire\ : std_logic;
signal \TVP_VSYNC_wire\ : std_logic;
signal \LED_wire\ : std_logic;
signal \ADV_HSYNC_wire\ : std_logic;
signal \ADV_VSYNC_wire\ : std_logic;
signal \tx_pll.TX_PLL_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);
signal \line_buffer.mem2_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem2_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem2_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem2_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem2_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem14_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem14_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem14_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem14_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem14_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem5_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem5_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem5_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem5_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem5_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem11_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem11_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem11_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem11_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem11_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem21_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem21_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem21_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem21_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem21_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem12_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem12_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem12_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem12_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem12_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem24_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem24_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem24_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem24_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem24_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem15_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem15_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem15_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem15_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem15_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem27_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem27_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem27_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem27_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem27_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem4_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem4_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem4_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem4_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem4_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem16_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem16_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem16_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem16_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem16_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem30_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem30_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem30_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem30_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem30_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem7_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem7_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem7_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem7_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem7_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem20_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem20_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem20_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem20_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem20_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem13_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem13_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem13_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem13_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem13_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem19_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem19_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem19_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem19_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem19_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem23_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem23_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem23_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem23_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem23_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem26_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem26_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem26_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem26_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem26_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem3_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem3_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem3_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem3_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem3_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem17_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem17_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem17_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem17_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem17_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem31_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem31_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem31_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem31_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem31_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem9_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem9_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem9_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem9_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem9_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem29_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem29_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem29_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem29_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem29_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem6_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem6_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem6_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem6_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem6_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem10_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem10_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem10_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem10_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem10_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem22_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem22_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem22_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem22_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem22_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem25_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem25_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem25_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem25_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem25_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem8_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem8_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem8_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem8_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem8_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem28_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem28_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem28_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem28_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem28_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem18_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem18_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem18_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \line_buffer.mem18_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \line_buffer.mem18_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    \TVP_CLK_wire\ <= TVP_CLK;
    ADV_CLK <= \ADV_CLK_wire\;
    \TVP_HSYNC_wire\ <= TVP_HSYNC;
    \TVP_VIDEO_wire\ <= TVP_VIDEO;
    ADV_G <= \ADV_G_wire\;
    ADV_R <= \ADV_R_wire\;
    ADV_B <= \ADV_B_wire\;
    ADV_SYNC_N <= \ADV_SYNC_N_wire\;
    ADV_BLANK_N <= \ADV_BLANK_N_wire\;
    \TVP_VSYNC_wire\ <= TVP_VSYNC;
    LED <= \LED_wire\;
    ADV_HSYNC <= \ADV_HSYNC_wire\;
    ADV_VSYNC <= \ADV_VSYNC_wire\;
    \tx_pll.TX_PLL_inst_DYNAMICDELAY_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.n474\ <= \line_buffer.mem2_physical_RDATA_wire\(11);
    \line_buffer.n473\ <= \line_buffer.mem2_physical_RDATA_wire\(3);
    \line_buffer.mem2_physical_RADDR_wire\ <= \N__13726\&\N__12214\&\N__10075\&\N__11095\&\N__11380\&\N__11947\&\N__11635\&\N__19339\&\N__20383\&\N__8833\&\N__13969\;
    \line_buffer.mem2_physical_WADDR_wire\ <= \N__17671\&\N__16225\&\N__15880\&\N__16516\&\N__16777\&\N__17032\&\N__17293\&\N__17902\&\N__15340\&\N__15592\&\N__18151\;
    \line_buffer.mem2_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem2_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__18580\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19135\&'0'&'0'&'0';
    \line_buffer.n561\ <= \line_buffer.mem14_physical_RDATA_wire\(11);
    \line_buffer.n560\ <= \line_buffer.mem14_physical_RDATA_wire\(3);
    \line_buffer.mem14_physical_RADDR_wire\ <= \N__13798\&\N__12286\&\N__10147\&\N__11167\&\N__11452\&\N__12019\&\N__11707\&\N__19411\&\N__20455\&\N__8905\&\N__14041\;
    \line_buffer.mem14_physical_WADDR_wire\ <= \N__17743\&\N__16297\&\N__15952\&\N__16588\&\N__16849\&\N__17104\&\N__17365\&\N__17974\&\N__15412\&\N__15664\&\N__18223\;
    \line_buffer.mem14_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem14_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__22506\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19002\&'0'&'0'&'0';
    \line_buffer.n571\ <= \line_buffer.mem5_physical_RDATA_wire\(11);
    \line_buffer.n570\ <= \line_buffer.mem5_physical_RDATA_wire\(3);
    \line_buffer.mem5_physical_RADDR_wire\ <= \N__13747\&\N__12223\&\N__10090\&\N__11116\&\N__11371\&\N__11968\&\N__11650\&\N__19348\&\N__20398\&\N__8836\&\N__13984\;
    \line_buffer.mem5_physical_WADDR_wire\ <= \N__17674\&\N__16222\&\N__15889\&\N__16525\&\N__16786\&\N__17047\&\N__17308\&\N__17911\&\N__15349\&\N__15601\&\N__18148\;
    \line_buffer.mem5_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem5_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__18591\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19146\&'0'&'0'&'0';
    \line_buffer.n529\ <= \line_buffer.mem11_physical_RDATA_wire\(11);
    \line_buffer.n528\ <= \line_buffer.mem11_physical_RDATA_wire\(3);
    \line_buffer.mem11_physical_RADDR_wire\ <= \N__13834\&\N__12322\&\N__10183\&\N__11203\&\N__11488\&\N__12055\&\N__11743\&\N__19447\&\N__20491\&\N__8941\&\N__14077\;
    \line_buffer.mem11_physical_WADDR_wire\ <= \N__17779\&\N__16333\&\N__15988\&\N__16624\&\N__16885\&\N__17140\&\N__17401\&\N__18010\&\N__15448\&\N__15700\&\N__18259\;
    \line_buffer.mem11_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem11_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__22518\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19034\&'0'&'0'&'0';
    \line_buffer.n591\ <= \line_buffer.mem21_physical_RDATA_wire\(11);
    \line_buffer.n590\ <= \line_buffer.mem21_physical_RDATA_wire\(3);
    \line_buffer.mem21_physical_RADDR_wire\ <= \N__13702\&\N__12190\&\N__10051\&\N__11071\&\N__11356\&\N__11923\&\N__11611\&\N__19315\&\N__20359\&\N__8809\&\N__13945\;
    \line_buffer.mem21_physical_WADDR_wire\ <= \N__17647\&\N__16201\&\N__15856\&\N__16492\&\N__16753\&\N__17008\&\N__17269\&\N__17878\&\N__15316\&\N__15568\&\N__18127\;
    \line_buffer.mem21_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem21_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__9068\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__10513\&'0'&'0'&'0';
    \line_buffer.n527\ <= \line_buffer.mem12_physical_RDATA_wire\(11);
    \line_buffer.n526\ <= \line_buffer.mem12_physical_RDATA_wire\(3);
    \line_buffer.mem12_physical_RADDR_wire\ <= \N__13822\&\N__12310\&\N__10171\&\N__11191\&\N__11476\&\N__12043\&\N__11731\&\N__19435\&\N__20479\&\N__8929\&\N__14065\;
    \line_buffer.mem12_physical_WADDR_wire\ <= \N__17767\&\N__16321\&\N__15976\&\N__16612\&\N__16873\&\N__17128\&\N__17389\&\N__17998\&\N__15436\&\N__15688\&\N__18247\;
    \line_buffer.mem12_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem12_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__9074\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__10475\&'0'&'0'&'0';
    \line_buffer.n535\ <= \line_buffer.mem24_physical_RDATA_wire\(11);
    \line_buffer.n534\ <= \line_buffer.mem24_physical_RDATA_wire\(3);
    \line_buffer.mem24_physical_RADDR_wire\ <= \N__13867\&\N__12343\&\N__10210\&\N__11236\&\N__11491\&\N__12088\&\N__11770\&\N__19468\&\N__20518\&\N__8956\&\N__14104\;
    \line_buffer.mem24_physical_WADDR_wire\ <= \N__17794\&\N__16342\&\N__16009\&\N__16645\&\N__16906\&\N__17167\&\N__17428\&\N__18031\&\N__15469\&\N__15721\&\N__18268\;
    \line_buffer.mem24_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem24_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__9057\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__10489\&'0'&'0'&'0';
    \line_buffer.n563\ <= \line_buffer.mem1_physical_RDATA_wire\(11);
    \line_buffer.n562\ <= \line_buffer.mem1_physical_RDATA_wire\(3);
    \line_buffer.mem1_physical_RADDR_wire\ <= \N__13858\&\N__12346\&\N__10207\&\N__11227\&\N__11507\&\N__12079\&\N__11767\&\N__19471\&\N__20515\&\N__8965\&\N__14101\;
    \line_buffer.mem1_physical_WADDR_wire\ <= \N__17803\&\N__16355\&\N__16012\&\N__16648\&\N__16909\&\N__17164\&\N__17425\&\N__18034\&\N__15472\&\N__15724\&\N__18281\;
    \line_buffer.mem1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__18557\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19119\&'0'&'0'&'0';
    \line_buffer.n559\ <= \line_buffer.mem15_physical_RDATA_wire\(11);
    \line_buffer.n558\ <= \line_buffer.mem15_physical_RDATA_wire\(3);
    \line_buffer.mem15_physical_RADDR_wire\ <= \N__13786\&\N__12274\&\N__10135\&\N__11155\&\N__11440\&\N__12007\&\N__11695\&\N__19399\&\N__20443\&\N__8893\&\N__14029\;
    \line_buffer.mem15_physical_WADDR_wire\ <= \N__17731\&\N__16285\&\N__15940\&\N__16576\&\N__16837\&\N__17092\&\N__17353\&\N__17962\&\N__15400\&\N__15652\&\N__18211\;
    \line_buffer.mem15_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem15_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__9069\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__10476\&'0'&'0'&'0';
    \line_buffer.n567\ <= \line_buffer.mem27_physical_RDATA_wire\(11);
    \line_buffer.n566\ <= \line_buffer.mem27_physical_RDATA_wire\(3);
    \line_buffer.mem27_physical_RADDR_wire\ <= \N__13831\&\N__12307\&\N__10174\&\N__11200\&\N__11455\&\N__12052\&\N__11734\&\N__19432\&\N__20482\&\N__8920\&\N__14068\;
    \line_buffer.mem27_physical_WADDR_wire\ <= \N__17758\&\N__16306\&\N__15973\&\N__16609\&\N__16870\&\N__17131\&\N__17392\&\N__17995\&\N__15433\&\N__15685\&\N__18232\;
    \line_buffer.mem27_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem27_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__9038\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__10482\&'0'&'0'&'0';
    \line_buffer.n539\ <= \line_buffer.mem4_physical_RDATA_wire\(11);
    \line_buffer.n538\ <= \line_buffer.mem4_physical_RDATA_wire\(3);
    \line_buffer.mem4_physical_RADDR_wire\ <= \N__13759\&\N__12235\&\N__10102\&\N__11128\&\N__11383\&\N__11980\&\N__11662\&\N__19360\&\N__20410\&\N__8848\&\N__13996\;
    \line_buffer.mem4_physical_WADDR_wire\ <= \N__17686\&\N__16234\&\N__15901\&\N__16537\&\N__16798\&\N__17059\&\N__17320\&\N__17923\&\N__15361\&\N__15613\&\N__18160\;
    \line_buffer.mem4_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem4_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__18581\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19136\&'0'&'0'&'0';
    \line_buffer.n557\ <= \line_buffer.mem16_physical_RDATA_wire\(11);
    \line_buffer.n556\ <= \line_buffer.mem16_physical_RDATA_wire\(3);
    \line_buffer.mem16_physical_RADDR_wire\ <= \N__13774\&\N__12262\&\N__10123\&\N__11143\&\N__11428\&\N__11995\&\N__11683\&\N__19387\&\N__20431\&\N__8881\&\N__14017\;
    \line_buffer.mem16_physical_WADDR_wire\ <= \N__17719\&\N__16273\&\N__15928\&\N__16564\&\N__16825\&\N__17080\&\N__17341\&\N__17950\&\N__15388\&\N__15640\&\N__18199\;
    \line_buffer.mem16_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem16_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__10601\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__10717\&'0'&'0'&'0';
    \line_buffer.n599\ <= \line_buffer.mem30_physical_RDATA_wire\(11);
    \line_buffer.n598\ <= \line_buffer.mem30_physical_RDATA_wire\(3);
    \line_buffer.mem30_physical_RADDR_wire\ <= \N__13783\&\N__12259\&\N__10126\&\N__11152\&\N__11407\&\N__12004\&\N__11686\&\N__19384\&\N__20434\&\N__8872\&\N__14020\;
    \line_buffer.mem30_physical_WADDR_wire\ <= \N__17710\&\N__16258\&\N__15925\&\N__16561\&\N__16822\&\N__17083\&\N__17344\&\N__17947\&\N__15385\&\N__15637\&\N__18184\;
    \line_buffer.mem30_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem30_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__9001\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__10496\&'0'&'0'&'0';
    \line_buffer.n466\ <= \line_buffer.mem7_physical_RDATA_wire\(11);
    \line_buffer.n465\ <= \line_buffer.mem7_physical_RDATA_wire\(3);
    \line_buffer.mem7_physical_RADDR_wire\ <= \N__13723\&\N__12199\&\N__10066\&\N__11092\&\N__11347\&\N__11944\&\N__11626\&\N__19324\&\N__20374\&\N__8812\&\N__13960\;
    \line_buffer.mem7_physical_WADDR_wire\ <= \N__17650\&\N__16198\&\N__15865\&\N__16501\&\N__16762\&\N__17023\&\N__17284\&\N__17887\&\N__15325\&\N__15577\&\N__18124\;
    \line_buffer.mem7_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem7_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__18596\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19148\&'0'&'0'&'0';
    \line_buffer.n593\ <= \line_buffer.mem20_physical_RDATA_wire\(11);
    \line_buffer.n592\ <= \line_buffer.mem20_physical_RDATA_wire\(3);
    \line_buffer.mem20_physical_RADDR_wire\ <= \N__13714\&\N__12202\&\N__10063\&\N__11083\&\N__11368\&\N__11935\&\N__11623\&\N__19327\&\N__20371\&\N__8821\&\N__13957\;
    \line_buffer.mem20_physical_WADDR_wire\ <= \N__17659\&\N__16213\&\N__15868\&\N__16504\&\N__16765\&\N__17020\&\N__17281\&\N__17890\&\N__15328\&\N__15580\&\N__18139\;
    \line_buffer.mem20_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem20_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__22517\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19043\&'0'&'0'&'0';
    \line_buffer.n525\ <= \line_buffer.mem13_physical_RDATA_wire\(11);
    \line_buffer.n524\ <= \line_buffer.mem13_physical_RDATA_wire\(3);
    \line_buffer.mem13_physical_RADDR_wire\ <= \N__13810\&\N__12298\&\N__10159\&\N__11179\&\N__11464\&\N__12031\&\N__11719\&\N__19423\&\N__20467\&\N__8917\&\N__14053\;
    \line_buffer.mem13_physical_WADDR_wire\ <= \N__17755\&\N__16309\&\N__15964\&\N__16600\&\N__16861\&\N__17116\&\N__17377\&\N__17986\&\N__15424\&\N__15676\&\N__18235\;
    \line_buffer.mem13_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem13_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__10600\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__10716\&'0'&'0'&'0';
    \line_buffer.n468\ <= \line_buffer.mem19_physical_RDATA_wire\(11);
    \line_buffer.n467\ <= \line_buffer.mem19_physical_RDATA_wire\(3);
    \line_buffer.mem19_physical_RADDR_wire\ <= \N__13738\&\N__12226\&\N__10087\&\N__11107\&\N__11392\&\N__11959\&\N__11647\&\N__19351\&\N__20395\&\N__8845\&\N__13981\;
    \line_buffer.mem19_physical_WADDR_wire\ <= \N__17683\&\N__16237\&\N__15892\&\N__16528\&\N__16789\&\N__17044\&\N__17305\&\N__17914\&\N__15352\&\N__15604\&\N__18163\;
    \line_buffer.mem19_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem19_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__10602\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__10728\&'0'&'0'&'0';
    \line_buffer.n537\ <= \line_buffer.mem23_physical_RDATA_wire\(11);
    \line_buffer.n536\ <= \line_buffer.mem23_physical_RDATA_wire\(3);
    \line_buffer.mem23_physical_RADDR_wire\ <= \N__13874\&\N__12355\&\N__10220\&\N__11243\&\N__11503\&\N__12095\&\N__11780\&\N__19480\&\N__20528\&\N__8968\&\N__14114\;
    \line_buffer.mem23_physical_WADDR_wire\ <= \N__17806\&\N__16354\&\N__16021\&\N__16657\&\N__16918\&\N__17177\&\N__17438\&\N__18043\&\N__15481\&\N__15733\&\N__18280\;
    \line_buffer.mem23_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem23_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__22523\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19006\&'0'&'0'&'0';
    \line_buffer.n531\ <= \line_buffer.mem0_physical_RDATA_wire\(11);
    \line_buffer.n530\ <= \line_buffer.mem0_physical_RDATA_wire\(3);
    \line_buffer.mem0_physical_RADDR_wire\ <= \N__13870\&\N__12356\&\N__10219\&\N__11239\&\N__11513\&\N__12091\&\N__11779\&\N__19481\&\N__20527\&\N__8972\&\N__14113\;
    \line_buffer.mem0_physical_WADDR_wire\ <= \N__17810\&\N__16361\&\N__16022\&\N__16658\&\N__16919\&\N__17176\&\N__17437\&\N__18044\&\N__15482\&\N__15734\&\N__18287\;
    \line_buffer.mem0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__18579\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19120\&'0'&'0'&'0';
    \line_buffer.n569\ <= \line_buffer.mem26_physical_RDATA_wire\(11);
    \line_buffer.n568\ <= \line_buffer.mem26_physical_RDATA_wire\(3);
    \line_buffer.mem26_physical_RADDR_wire\ <= \N__13843\&\N__12319\&\N__10186\&\N__11212\&\N__11467\&\N__12064\&\N__11746\&\N__19444\&\N__20494\&\N__8932\&\N__14080\;
    \line_buffer.mem26_physical_WADDR_wire\ <= \N__17770\&\N__16318\&\N__15985\&\N__16621\&\N__16882\&\N__17143\&\N__17404\&\N__18007\&\N__15445\&\N__15697\&\N__18244\;
    \line_buffer.mem26_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem26_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__22513\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19021\&'0'&'0'&'0';
    \line_buffer.n595\ <= \line_buffer.mem3_physical_RDATA_wire\(11);
    \line_buffer.n594\ <= \line_buffer.mem3_physical_RDATA_wire\(3);
    \line_buffer.mem3_physical_RADDR_wire\ <= \N__13795\&\N__12271\&\N__10138\&\N__11164\&\N__11419\&\N__12016\&\N__11698\&\N__19396\&\N__20446\&\N__8884\&\N__14032\;
    \line_buffer.mem3_physical_WADDR_wire\ <= \N__17722\&\N__16270\&\N__15937\&\N__16573\&\N__16834\&\N__17095\&\N__17356\&\N__17959\&\N__15397\&\N__15649\&\N__18196\;
    \line_buffer.mem3_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem3_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__18556\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19111\&'0'&'0'&'0';
    \line_buffer.n472\ <= \line_buffer.mem17_physical_RDATA_wire\(11);
    \line_buffer.n471\ <= \line_buffer.mem17_physical_RDATA_wire\(3);
    \line_buffer.mem17_physical_RADDR_wire\ <= \N__13762\&\N__12250\&\N__10111\&\N__11131\&\N__11416\&\N__11983\&\N__11671\&\N__19375\&\N__20419\&\N__8869\&\N__14005\;
    \line_buffer.mem17_physical_WADDR_wire\ <= \N__17707\&\N__16261\&\N__15916\&\N__16552\&\N__16813\&\N__17068\&\N__17329\&\N__17938\&\N__15376\&\N__15628\&\N__18187\;
    \line_buffer.mem17_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem17_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__22483\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19036\&'0'&'0'&'0';
    \line_buffer.n597\ <= \line_buffer.mem31_physical_RDATA_wire\(11);
    \line_buffer.n596\ <= \line_buffer.mem31_physical_RDATA_wire\(3);
    \line_buffer.mem31_physical_RADDR_wire\ <= \N__13771\&\N__12247\&\N__10114\&\N__11140\&\N__11395\&\N__11992\&\N__11674\&\N__19372\&\N__20422\&\N__8860\&\N__14008\;
    \line_buffer.mem31_physical_WADDR_wire\ <= \N__17698\&\N__16246\&\N__15913\&\N__16549\&\N__16810\&\N__17071\&\N__17332\&\N__17935\&\N__15373\&\N__15625\&\N__18172\;
    \line_buffer.mem31_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem31_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__10610\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__10736\&'0'&'0'&'0';
    \line_buffer.n462\ <= \line_buffer.mem9_physical_RDATA_wire\(11);
    \line_buffer.n461\ <= \line_buffer.mem9_physical_RDATA_wire\(3);
    \line_buffer.mem9_physical_RADDR_wire\ <= \N__13699\&\N__12175\&\N__10042\&\N__11068\&\N__11323\&\N__11920\&\N__11602\&\N__19300\&\N__20350\&\N__8788\&\N__13936\;
    \line_buffer.mem9_physical_WADDR_wire\ <= \N__17626\&\N__16174\&\N__15841\&\N__16477\&\N__16738\&\N__16999\&\N__17260\&\N__17863\&\N__15301\&\N__15553\&\N__18100\;
    \line_buffer.mem9_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem9_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__9058\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__10517\&'0'&'0'&'0';
    \line_buffer.n601\ <= \line_buffer.mem29_physical_RDATA_wire\(11);
    \line_buffer.n600\ <= \line_buffer.mem29_physical_RDATA_wire\(3);
    \line_buffer.mem29_physical_RADDR_wire\ <= \N__13807\&\N__12283\&\N__10150\&\N__11176\&\N__11431\&\N__12028\&\N__11710\&\N__19408\&\N__20458\&\N__8896\&\N__14044\;
    \line_buffer.mem29_physical_WADDR_wire\ <= \N__17734\&\N__16282\&\N__15949\&\N__16585\&\N__16846\&\N__17107\&\N__17368\&\N__17971\&\N__15409\&\N__15661\&\N__18208\;
    \line_buffer.mem29_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem29_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__22519\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19001\&'0'&'0'&'0';
    \line_buffer.n603\ <= \line_buffer.mem6_physical_RDATA_wire\(11);
    \line_buffer.n602\ <= \line_buffer.mem6_physical_RDATA_wire\(3);
    \line_buffer.mem6_physical_RADDR_wire\ <= \N__13735\&\N__12211\&\N__10078\&\N__11104\&\N__11359\&\N__11956\&\N__11638\&\N__19336\&\N__20386\&\N__8824\&\N__13972\;
    \line_buffer.mem6_physical_WADDR_wire\ <= \N__17662\&\N__16210\&\N__15877\&\N__16513\&\N__16774\&\N__17035\&\N__17296\&\N__17899\&\N__15337\&\N__15589\&\N__18136\;
    \line_buffer.mem6_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem6_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__18592\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19147\&'0'&'0'&'0';
    \line_buffer.n460\ <= \line_buffer.mem10_physical_RDATA_wire\(11);
    \line_buffer.n459\ <= \line_buffer.mem10_physical_RDATA_wire\(3);
    \line_buffer.mem10_physical_RADDR_wire\ <= \N__13846\&\N__12334\&\N__10195\&\N__11215\&\N__11500\&\N__12067\&\N__11755\&\N__19459\&\N__20503\&\N__8953\&\N__14089\;
    \line_buffer.mem10_physical_WADDR_wire\ <= \N__17791\&\N__16345\&\N__16000\&\N__16636\&\N__16897\&\N__17152\&\N__17413\&\N__18022\&\N__15460\&\N__15712\&\N__18271\;
    \line_buffer.mem10_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem10_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__10599\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__10715\&'0'&'0'&'0';
    \line_buffer.n589\ <= \line_buffer.mem22_physical_RDATA_wire\(11);
    \line_buffer.n588\ <= \line_buffer.mem22_physical_RDATA_wire\(3);
    \line_buffer.mem22_physical_RADDR_wire\ <= \N__13690\&\N__12178\&\N__10039\&\N__11059\&\N__11344\&\N__11911\&\N__11599\&\N__19303\&\N__20347\&\N__8797\&\N__13933\;
    \line_buffer.mem22_physical_WADDR_wire\ <= \N__17635\&\N__16189\&\N__15844\&\N__16480\&\N__16741\&\N__16996\&\N__17257\&\N__17866\&\N__15304\&\N__15556\&\N__18115\;
    \line_buffer.mem22_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem22_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__10609\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__10735\&'0'&'0'&'0';
    \line_buffer.n533\ <= \line_buffer.mem25_physical_RDATA_wire\(11);
    \line_buffer.n532\ <= \line_buffer.mem25_physical_RDATA_wire\(3);
    \line_buffer.mem25_physical_RADDR_wire\ <= \N__13855\&\N__12331\&\N__10198\&\N__11224\&\N__11479\&\N__12076\&\N__11758\&\N__19456\&\N__20506\&\N__8944\&\N__14092\;
    \line_buffer.mem25_physical_WADDR_wire\ <= \N__17782\&\N__16330\&\N__15997\&\N__16633\&\N__16894\&\N__17155\&\N__17416\&\N__18019\&\N__15457\&\N__15709\&\N__18256\;
    \line_buffer.mem25_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem25_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__10594\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__10708\&'0'&'0'&'0';
    \line_buffer.n464\ <= \line_buffer.mem8_physical_RDATA_wire\(11);
    \line_buffer.n463\ <= \line_buffer.mem8_physical_RDATA_wire\(3);
    \line_buffer.mem8_physical_RADDR_wire\ <= \N__13711\&\N__12187\&\N__10054\&\N__11080\&\N__11335\&\N__11932\&\N__11614\&\N__19312\&\N__20362\&\N__8800\&\N__13948\;
    \line_buffer.mem8_physical_WADDR_wire\ <= \N__17638\&\N__16186\&\N__15853\&\N__16489\&\N__16750\&\N__17011\&\N__17272\&\N__17875\&\N__15313\&\N__15565\&\N__18112\;
    \line_buffer.mem8_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem8_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__22496\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__19035\&'0'&'0'&'0';
    \line_buffer.n565\ <= \line_buffer.mem28_physical_RDATA_wire\(11);
    \line_buffer.n564\ <= \line_buffer.mem28_physical_RDATA_wire\(3);
    \line_buffer.mem28_physical_RADDR_wire\ <= \N__13819\&\N__12295\&\N__10162\&\N__11188\&\N__11443\&\N__12040\&\N__11722\&\N__19420\&\N__20470\&\N__8908\&\N__14056\;
    \line_buffer.mem28_physical_WADDR_wire\ <= \N__17746\&\N__16294\&\N__15961\&\N__16597\&\N__16858\&\N__17119\&\N__17380\&\N__17983\&\N__15421\&\N__15673\&\N__18220\;
    \line_buffer.mem28_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem28_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__10595\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__10724\&'0'&'0'&'0';
    \line_buffer.n470\ <= \line_buffer.mem18_physical_RDATA_wire\(11);
    \line_buffer.n469\ <= \line_buffer.mem18_physical_RDATA_wire\(3);
    \line_buffer.mem18_physical_RADDR_wire\ <= \N__13750\&\N__12238\&\N__10099\&\N__11119\&\N__11404\&\N__11971\&\N__11659\&\N__19363\&\N__20407\&\N__8857\&\N__13993\;
    \line_buffer.mem18_physical_WADDR_wire\ <= \N__17695\&\N__16249\&\N__15904\&\N__16540\&\N__16801\&\N__17056\&\N__17317\&\N__17926\&\N__15364\&\N__15616\&\N__18175\;
    \line_buffer.mem18_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \line_buffer.mem18_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__9070\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__10500\&'0'&'0'&'0';

    \tx_pll.TX_PLL_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "010",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "100",
            DIVF => "0100110",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            LATCHINPUTVALUE => '0',
            SCLK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => \ADV_CLK_c\,
            REFERENCECLK => \N__16120\,
            RESETB => \N__24513\,
            BYPASS => \GNDG0\,
            SDI => '0',
            DYNAMICDELAY => \tx_pll.TX_PLL_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => OPEN
        );

    \line_buffer.mem2_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_E => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_D => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_C => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_B => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_A => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_9 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_8 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_7 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_6 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_5 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_4 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_3 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_2 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_1 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_0 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001"
        )
    port map (
            RDATA => \line_buffer.mem2_physical_RDATA_wire\,
            RADDR => \line_buffer.mem2_physical_RADDR_wire\,
            WADDR => \line_buffer.mem2_physical_WADDR_wire\,
            MASK => \line_buffer.mem2_physical_MASK_wire\,
            WDATA => \line_buffer.mem2_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23413\,
            RE => \N__24378\,
            WCLKE => 'H',
            WCLK => \N__24162\,
            WE => \N__13076\
        );

    \line_buffer.mem14_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_E => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_D => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_C => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_B => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_A => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_9 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_8 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_7 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_6 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_5 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_4 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_3 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011",
            INIT_2 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011",
            INIT_1 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011",
            INIT_0 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011"
        )
    port map (
            RDATA => \line_buffer.mem14_physical_RDATA_wire\,
            RADDR => \line_buffer.mem14_physical_RADDR_wire\,
            WADDR => \line_buffer.mem14_physical_WADDR_wire\,
            MASK => \line_buffer.mem14_physical_MASK_wire\,
            WDATA => \line_buffer.mem14_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23510\,
            RE => \N__24363\,
            WCLKE => 'H',
            WCLK => \N__24142\,
            WE => \N__12890\
        );

    \line_buffer.mem5_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_E => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_D => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_C => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_B => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_A => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_9 => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_8 => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_7 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_6 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_5 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_4 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_3 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110",
            INIT_2 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110",
            INIT_1 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110",
            INIT_0 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110"
        )
    port map (
            RDATA => \line_buffer.mem5_physical_RDATA_wire\,
            RADDR => \line_buffer.mem5_physical_RADDR_wire\,
            WADDR => \line_buffer.mem5_physical_WADDR_wire\,
            MASK => \line_buffer.mem5_physical_MASK_wire\,
            WDATA => \line_buffer.mem5_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22912\,
            RE => \N__24409\,
            WCLKE => 'H',
            WCLK => \N__24160\,
            WE => \N__14753\
        );

    \line_buffer.mem11_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_E => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_D => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_C => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_B => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_A => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_9 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_8 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_7 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_6 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_5 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_4 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_3 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_2 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_1 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_0 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100"
        )
    port map (
            RDATA => \line_buffer.mem11_physical_RDATA_wire\,
            RADDR => \line_buffer.mem11_physical_RADDR_wire\,
            WADDR => \line_buffer.mem11_physical_WADDR_wire\,
            MASK => \line_buffer.mem11_physical_MASK_wire\,
            WDATA => \line_buffer.mem11_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23688\,
            RE => \N__24454\,
            WCLKE => 'H',
            WCLK => \N__24130\,
            WE => \N__13024\
        );

    \line_buffer.mem21_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_E => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_D => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_C => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_B => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_A => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_9 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_8 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_7 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_6 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_5 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_4 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_3 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_2 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_1 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_0 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011"
        )
    port map (
            RDATA => \line_buffer.mem21_physical_RDATA_wire\,
            RADDR => \line_buffer.mem21_physical_RADDR_wire\,
            WADDR => \line_buffer.mem21_physical_WADDR_wire\,
            MASK => \line_buffer.mem21_physical_MASK_wire\,
            WDATA => \line_buffer.mem21_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23249\,
            RE => \N__24425\,
            WCLKE => 'H',
            WCLK => \N__24166\,
            WE => \N__13414\
        );

    \line_buffer.mem12_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_E => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_D => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_C => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_B => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_A => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_9 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_8 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_7 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_6 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_5 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_4 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_3 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_2 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_1 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_0 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100"
        )
    port map (
            RDATA => \line_buffer.mem12_physical_RDATA_wire\,
            RADDR => \line_buffer.mem12_physical_RADDR_wire\,
            WADDR => \line_buffer.mem12_physical_WADDR_wire\,
            MASK => \line_buffer.mem12_physical_MASK_wire\,
            WDATA => \line_buffer.mem12_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23621\,
            RE => \N__24412\,
            WCLKE => 'H',
            WCLK => \N__24136\,
            WE => \N__13017\
        );

    \line_buffer.mem24_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_E => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_D => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_C => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_B => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_A => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_9 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_8 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_7 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_6 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_5 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_4 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_3 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_2 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_1 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_0 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001"
        )
    port map (
            RDATA => \line_buffer.mem24_physical_RDATA_wire\,
            RADDR => \line_buffer.mem24_physical_RADDR_wire\,
            WADDR => \line_buffer.mem24_physical_WADDR_wire\,
            MASK => \line_buffer.mem24_physical_MASK_wire\,
            WDATA => \line_buffer.mem24_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23734\,
            RE => \N__24523\,
            WCLKE => 'H',
            WCLK => \N__24117\,
            WE => \N__12639\
        );

    \line_buffer.mem1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_E => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_D => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_C => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_B => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_A => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_9 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_8 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_7 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_6 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_5 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_4 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_3 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011",
            INIT_2 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011",
            INIT_1 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011",
            INIT_0 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011"
        )
    port map (
            RDATA => \line_buffer.mem1_physical_RDATA_wire\,
            RADDR => \line_buffer.mem1_physical_RADDR_wire\,
            WADDR => \line_buffer.mem1_physical_WADDR_wire\,
            MASK => \line_buffer.mem1_physical_MASK_wire\,
            WDATA => \line_buffer.mem1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23722\,
            RE => \N__24488\,
            WCLKE => 'H',
            WCLK => \N__24113\,
            WE => \N__12902\
        );

    \line_buffer.mem15_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_E => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_D => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_C => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_B => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_A => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_9 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_8 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_7 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_6 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_5 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_4 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_3 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011",
            INIT_2 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011",
            INIT_1 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011",
            INIT_0 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011"
        )
    port map (
            RDATA => \line_buffer.mem15_physical_RDATA_wire\,
            RADDR => \line_buffer.mem15_physical_RADDR_wire\,
            WADDR => \line_buffer.mem15_physical_WADDR_wire\,
            MASK => \line_buffer.mem15_physical_MASK_wire\,
            WDATA => \line_buffer.mem15_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23509\,
            RE => \N__24342\,
            WCLKE => 'H',
            WCLK => \N__24144\,
            WE => \N__12900\
        );

    \line_buffer.mem27_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_E => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_D => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_C => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_B => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_A => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_9 => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_8 => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_7 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_6 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_5 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_4 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_3 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110",
            INIT_2 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110",
            INIT_1 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110",
            INIT_0 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110"
        )
    port map (
            RDATA => \line_buffer.mem27_physical_RDATA_wire\,
            RADDR => \line_buffer.mem27_physical_RADDR_wire\,
            WADDR => \line_buffer.mem27_physical_WADDR_wire\,
            MASK => \line_buffer.mem27_physical_MASK_wire\,
            WDATA => \line_buffer.mem27_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23696\,
            RE => \N__24496\,
            WCLKE => 'H',
            WCLK => \N__24137\,
            WE => \N__14748\
        );

    \line_buffer.mem4_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_E => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_D => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_C => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_B => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_A => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_9 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_8 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_7 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_6 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_5 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_4 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_3 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_2 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_1 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_0 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001"
        )
    port map (
            RDATA => \line_buffer.mem4_physical_RDATA_wire\,
            RADDR => \line_buffer.mem4_physical_RADDR_wire\,
            WADDR => \line_buffer.mem4_physical_WADDR_wire\,
            MASK => \line_buffer.mem4_physical_MASK_wire\,
            WDATA => \line_buffer.mem4_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23403\,
            RE => \N__24468\,
            WCLKE => 'H',
            WCLK => \N__24158\,
            WE => \N__12640\
        );

    \line_buffer.mem16_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_E => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_D => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_C => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_B => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_A => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_9 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_8 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_7 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_6 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_5 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_4 => "0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011",
            INIT_3 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011",
            INIT_2 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011",
            INIT_1 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011",
            INIT_0 => "0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011"
        )
    port map (
            RDATA => \line_buffer.mem16_physical_RDATA_wire\,
            RADDR => \line_buffer.mem16_physical_RADDR_wire\,
            WADDR => \line_buffer.mem16_physical_WADDR_wire\,
            MASK => \line_buffer.mem16_physical_MASK_wire\,
            WDATA => \line_buffer.mem16_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23358\,
            RE => \N__24322\,
            WCLKE => 'H',
            WCLK => \N__24147\,
            WE => \N__12901\
        );

    \line_buffer.mem30_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_E => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_D => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_C => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_B => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_A => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_9 => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_8 => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_7 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_6 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_5 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_4 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_3 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110",
            INIT_2 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110",
            INIT_1 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110",
            INIT_0 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110"
        )
    port map (
            RDATA => \line_buffer.mem30_physical_RDATA_wire\,
            RADDR => \line_buffer.mem30_physical_RADDR_wire\,
            WADDR => \line_buffer.mem30_physical_WADDR_wire\,
            MASK => \line_buffer.mem30_physical_MASK_wire\,
            WDATA => \line_buffer.mem30_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23527\,
            RE => \N__24435\,
            WCLKE => 'H',
            WCLK => \N__24152\,
            WE => \N__15024\
        );

    \line_buffer.mem7_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_E => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_D => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_C => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_B => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_A => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_9 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_8 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_7 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_6 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_5 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_4 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_3 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_2 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_1 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_0 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000"
        )
    port map (
            RDATA => \line_buffer.mem7_physical_RDATA_wire\,
            RADDR => \line_buffer.mem7_physical_RADDR_wire\,
            WADDR => \line_buffer.mem7_physical_WADDR_wire\,
            MASK => \line_buffer.mem7_physical_MASK_wire\,
            WDATA => \line_buffer.mem7_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23298\,
            RE => \N__24521\,
            WCLKE => 'H',
            WCLK => \N__24165\,
            WE => \N__14987\
        );

    \line_buffer.mem20_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_E => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_D => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_C => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_B => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_A => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_9 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_8 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_7 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_6 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_5 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_4 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_3 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_2 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_1 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_0 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011"
        )
    port map (
            RDATA => \line_buffer.mem20_physical_RDATA_wire\,
            RADDR => \line_buffer.mem20_physical_RADDR_wire\,
            WADDR => \line_buffer.mem20_physical_WADDR_wire\,
            MASK => \line_buffer.mem20_physical_MASK_wire\,
            WDATA => \line_buffer.mem20_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23552\,
            RE => \N__24424\,
            WCLKE => 'H',
            WCLK => \N__24164\,
            WE => \N__13413\
        );

    \line_buffer.mem13_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_E => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_D => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_C => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_B => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_A => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_9 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_8 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_7 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_6 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_5 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_4 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_3 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_2 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_1 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_0 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100"
        )
    port map (
            RDATA => \line_buffer.mem13_physical_RDATA_wire\,
            RADDR => \line_buffer.mem13_physical_RADDR_wire\,
            WADDR => \line_buffer.mem13_physical_WADDR_wire\,
            MASK => \line_buffer.mem13_physical_MASK_wire\,
            WDATA => \line_buffer.mem13_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23620\,
            RE => \N__24411\,
            WCLKE => 'H',
            WCLK => \N__24138\,
            WE => \N__13016\
        );

    \line_buffer.mem19_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_E => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_D => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_C => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_B => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_A => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_9 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_8 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_7 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_6 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_5 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_4 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_3 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_2 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_1 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_0 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001"
        )
    port map (
            RDATA => \line_buffer.mem19_physical_RDATA_wire\,
            RADDR => \line_buffer.mem19_physical_RADDR_wire\,
            WADDR => \line_buffer.mem19_physical_WADDR_wire\,
            MASK => \line_buffer.mem19_physical_MASK_wire\,
            WDATA => \line_buffer.mem19_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23023\,
            RE => \N__24377\,
            WCLKE => 'H',
            WCLK => \N__24159\,
            WE => \N__13072\
        );

    \line_buffer.mem23_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_E => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_D => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_C => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_B => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_A => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_9 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_8 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_7 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_6 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_5 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_4 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_3 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_2 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_1 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_0 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001"
        )
    port map (
            RDATA => \line_buffer.mem23_physical_RDATA_wire\,
            RADDR => \line_buffer.mem23_physical_RADDR_wire\,
            WADDR => \line_buffer.mem23_physical_WADDR_wire\,
            MASK => \line_buffer.mem23_physical_MASK_wire\,
            WDATA => \line_buffer.mem23_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23735\,
            RE => \N__24524\,
            WCLKE => 'H',
            WCLK => \N__24109\,
            WE => \N__12641\
        );

    \line_buffer.mem0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_E => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_D => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_C => "1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110",
            INIT_B => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_A => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_9 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_8 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_7 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_6 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_5 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_4 => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_3 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_2 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_1 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_0 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100"
        )
    port map (
            RDATA => \line_buffer.mem0_physical_RDATA_wire\,
            RADDR => \line_buffer.mem0_physical_RADDR_wire\,
            WADDR => \line_buffer.mem0_physical_WADDR_wire\,
            MASK => \line_buffer.mem0_physical_MASK_wire\,
            WDATA => \line_buffer.mem0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23723\,
            RE => \N__24489\,
            WCLKE => 'H',
            WCLK => \N__24104\,
            WE => \N__13028\
        );

    \line_buffer.mem26_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_E => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_D => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_C => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_B => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_A => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_9 => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_8 => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_7 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_6 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_5 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_4 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_3 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110",
            INIT_2 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110",
            INIT_1 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110",
            INIT_0 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110"
        )
    port map (
            RDATA => \line_buffer.mem26_physical_RDATA_wire\,
            RADDR => \line_buffer.mem26_physical_RADDR_wire\,
            WADDR => \line_buffer.mem26_physical_WADDR_wire\,
            MASK => \line_buffer.mem26_physical_MASK_wire\,
            WDATA => \line_buffer.mem26_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23724\,
            RE => \N__24408\,
            WCLKE => 'H',
            WCLK => \N__24134\,
            WE => \N__14749\
        );

    \line_buffer.mem3_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_E => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_D => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_C => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_B => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_A => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_9 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_8 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_7 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_6 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_5 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_4 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_3 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_2 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_1 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_0 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011"
        )
    port map (
            RDATA => \line_buffer.mem3_physical_RDATA_wire\,
            RADDR => \line_buffer.mem3_physical_RADDR_wire\,
            WADDR => \line_buffer.mem3_physical_WADDR_wire\,
            MASK => \line_buffer.mem3_physical_MASK_wire\,
            WDATA => \line_buffer.mem3_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23478\,
            RE => \N__24469\,
            WCLKE => 'H',
            WCLK => \N__24145\,
            WE => \N__13403\
        );

    \line_buffer.mem17_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_E => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_D => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_C => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_B => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_A => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_9 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_8 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_7 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_6 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_5 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_4 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_3 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_2 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_1 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_0 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001"
        )
    port map (
            RDATA => \line_buffer.mem17_physical_RDATA_wire\,
            RADDR => \line_buffer.mem17_physical_RADDR_wire\,
            WADDR => \line_buffer.mem17_physical_WADDR_wire\,
            MASK => \line_buffer.mem17_physical_MASK_wire\,
            WDATA => \line_buffer.mem17_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23357\,
            RE => \N__24269\,
            WCLKE => 'H',
            WCLK => \N__24153\,
            WE => \N__13061\
        );

    \line_buffer.mem31_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_E => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_D => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_C => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_B => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_A => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_9 => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_8 => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_7 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_6 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_5 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_4 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_3 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110",
            INIT_2 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110",
            INIT_1 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110",
            INIT_0 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110"
        )
    port map (
            RDATA => \line_buffer.mem31_physical_RDATA_wire\,
            RADDR => \line_buffer.mem31_physical_RADDR_wire\,
            WADDR => \line_buffer.mem31_physical_WADDR_wire\,
            MASK => \line_buffer.mem31_physical_MASK_wire\,
            WDATA => \line_buffer.mem31_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23331\,
            RE => \N__24343\,
            WCLKE => 'H',
            WCLK => \N__24154\,
            WE => \N__15031\
        );

    \line_buffer.mem9_physical\ : SB_RAM40_4K
    generic map (
            INIT_0 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_E => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_D => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_C => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_B => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_A => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_9 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_8 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_7 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_6 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_5 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_4 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_3 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_2 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_1 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000"
        )
    port map (
            RDATA => \line_buffer.mem9_physical_RDATA_wire\,
            RADDR => \line_buffer.mem9_physical_RADDR_wire\,
            WADDR => \line_buffer.mem9_physical_WADDR_wire\,
            MASK => \line_buffer.mem9_physical_MASK_wire\,
            WDATA => \line_buffer.mem9_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__22955\,
            RE => \N__24407\,
            WCLKE => 'H',
            WCLK => \N__24169\,
            WE => \N__14993\
        );

    \line_buffer.mem29_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_E => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_D => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_C => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_B => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_A => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_9 => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_8 => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_7 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_6 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_5 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_4 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_3 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110",
            INIT_2 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110",
            INIT_1 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110",
            INIT_0 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110"
        )
    port map (
            RDATA => \line_buffer.mem29_physical_RDATA_wire\,
            RADDR => \line_buffer.mem29_physical_RADDR_wire\,
            WADDR => \line_buffer.mem29_physical_WADDR_wire\,
            MASK => \line_buffer.mem29_physical_MASK_wire\,
            WDATA => \line_buffer.mem29_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23636\,
            RE => \N__24470\,
            WCLKE => 'H',
            WCLK => \N__24143\,
            WE => \N__15015\
        );

    \line_buffer.mem6_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_E => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_D => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_C => "1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011",
            INIT_B => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_A => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_9 => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_8 => "1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011",
            INIT_7 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_6 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_5 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_4 => "1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111",
            INIT_3 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110",
            INIT_2 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110",
            INIT_1 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110",
            INIT_0 => "1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110"
        )
    port map (
            RDATA => \line_buffer.mem6_physical_RDATA_wire\,
            RADDR => \line_buffer.mem6_physical_RADDR_wire\,
            WADDR => \line_buffer.mem6_physical_WADDR_wire\,
            MASK => \line_buffer.mem6_physical_MASK_wire\,
            WDATA => \line_buffer.mem6_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23466\,
            RE => \N__24505\,
            WCLKE => 'H',
            WCLK => \N__24163\,
            WE => \N__15035\
        );

    \line_buffer.mem10_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_E => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_D => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_C => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_B => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_A => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_9 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_8 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_7 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_6 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_5 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_4 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_3 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_2 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_1 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_0 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000"
        )
    port map (
            RDATA => \line_buffer.mem10_physical_RDATA_wire\,
            RADDR => \line_buffer.mem10_physical_RADDR_wire\,
            WADDR => \line_buffer.mem10_physical_WADDR_wire\,
            MASK => \line_buffer.mem10_physical_MASK_wire\,
            WDATA => \line_buffer.mem10_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23689\,
            RE => \N__24455\,
            WCLKE => 'H',
            WCLK => \N__24120\,
            WE => \N__14992\
        );

    \line_buffer.mem22_physical\ : SB_RAM40_4K
    generic map (
            INIT_0 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_E => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_D => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_C => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_B => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_A => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_9 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_8 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_7 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_6 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_5 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_4 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_3 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_2 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011",
            INIT_1 => "0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011"
        )
    port map (
            RDATA => \line_buffer.mem22_physical_RDATA_wire\,
            RADDR => \line_buffer.mem22_physical_RADDR_wire\,
            WADDR => \line_buffer.mem22_physical_WADDR_wire\,
            MASK => \line_buffer.mem22_physical_MASK_wire\,
            WDATA => \line_buffer.mem22_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23253\,
            RE => \N__24462\,
            WCLKE => 'H',
            WCLK => \N__24168\,
            WE => \N__13418\
        );

    \line_buffer.mem25_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_E => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_D => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_C => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_B => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_A => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_9 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_8 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_7 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_6 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_5 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_4 => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_3 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_2 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_1 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_0 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001"
        )
    port map (
            RDATA => \line_buffer.mem25_physical_RDATA_wire\,
            RADDR => \line_buffer.mem25_physical_RADDR_wire\,
            WADDR => \line_buffer.mem25_physical_WADDR_wire\,
            MASK => \line_buffer.mem25_physical_MASK_wire\,
            WDATA => \line_buffer.mem25_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23730\,
            RE => \N__24514\,
            WCLKE => 'H',
            WCLK => \N__24126\,
            WE => \N__12626\
        );

    \line_buffer.mem8_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_E => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_D => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_C => "1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100",
            INIT_B => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_A => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_9 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_8 => "1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100",
            INIT_7 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_6 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_5 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_4 => "1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100",
            INIT_3 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_2 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_1 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000",
            INIT_0 => "1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000"
        )
    port map (
            RDATA => \line_buffer.mem8_physical_RDATA_wire\,
            RADDR => \line_buffer.mem8_physical_RADDR_wire\,
            WADDR => \line_buffer.mem8_physical_WADDR_wire\,
            MASK => \line_buffer.mem8_physical_MASK_wire\,
            WDATA => \line_buffer.mem8_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23083\,
            RE => \N__24522\,
            WCLKE => 'H',
            WCLK => \N__24167\,
            WE => \N__14988\
        );

    \line_buffer.mem28_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_E => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_D => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_C => "0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111",
            INIT_B => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_A => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_9 => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_8 => "0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110",
            INIT_7 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_6 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_5 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_4 => "1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110",
            INIT_3 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110",
            INIT_2 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110",
            INIT_1 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110",
            INIT_0 => "1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110"
        )
    port map (
            RDATA => \line_buffer.mem28_physical_RDATA_wire\,
            RADDR => \line_buffer.mem28_physical_RADDR_wire\,
            WADDR => \line_buffer.mem28_physical_WADDR_wire\,
            MASK => \line_buffer.mem28_physical_MASK_wire\,
            WDATA => \line_buffer.mem28_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23037\,
            RE => \N__24410\,
            WCLKE => 'H',
            WCLK => \N__24140\,
            WE => \N__14741\
        );

    \line_buffer.mem18_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_F => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_E => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_D => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_C => "1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001",
            INIT_B => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_A => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_9 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_8 => "0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001",
            INIT_7 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_6 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_5 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_4 => "0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001",
            INIT_3 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_2 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_1 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001",
            INIT_0 => "0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001"
        )
    port map (
            RDATA => \line_buffer.mem18_physical_RDATA_wire\,
            RADDR => \line_buffer.mem18_physical_RADDR_wire\,
            WADDR => \line_buffer.mem18_physical_WADDR_wire\,
            MASK => \line_buffer.mem18_physical_MASK_wire\,
            WDATA => \line_buffer.mem18_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__23184\,
            RE => \N__24323\,
            WCLKE => 'H',
            WCLK => \N__24156\,
            WE => \N__13071\
        );

    \DEBUG_c_3_pad_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__25263\,
            GLOBALBUFFEROUTPUT => \DEBUG_c_3_c\
        );

    \DEBUG_c_3_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__25265\,
            DIN => \N__25264\,
            DOUT => \N__25263\,
            PACKAGEPIN => \TVP_CLK_wire\
        );

    \DEBUG_c_3_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25265\,
            PADOUT => \N__25264\,
            PADIN => \N__25263\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_CLK_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25254\,
            DIN => \N__25253\,
            DOUT => \N__25252\,
            PACKAGEPIN => \ADV_CLK_wire\
        );

    \ADV_CLK_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25254\,
            PADOUT => \N__25253\,
            PADIN => \N__25252\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__23278\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_c_2_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__25245\,
            DIN => \N__25244\,
            DOUT => \N__25243\,
            PACKAGEPIN => \TVP_HSYNC_wire\
        );

    \DEBUG_c_2_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25245\,
            PADOUT => \N__25244\,
            PADIN => \N__25243\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DEBUG_c_2_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__25236\,
            DIN => \N__25235\,
            DOUT => \N__25234\,
            PACKAGEPIN => DEBUG(3)
        );

    \DEBUG_pad_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25236\,
            PADOUT => \N__25235\,
            PADIN => \N__25234\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__16121\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_VIDEO_pad_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__25227\,
            DIN => \N__25226\,
            DOUT => \N__25225\,
            PACKAGEPIN => \TVP_VIDEO_wire\(2)
        );

    \TVP_VIDEO_pad_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25227\,
            PADOUT => \N__25226\,
            PADIN => \N__25225\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_VIDEO_c_2\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25218\,
            DIN => \N__25217\,
            DOUT => \N__25216\,
            PACKAGEPIN => \ADV_G_wire\(5)
        );

    \ADV_G_pad_5_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25218\,
            PADOUT => \N__25217\,
            PADIN => \N__25216\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__21994\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25209\,
            DIN => \N__25208\,
            DOUT => \N__25207\,
            PACKAGEPIN => \ADV_R_wire\(3)
        );

    \ADV_R_pad_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25209\,
            PADOUT => \N__25208\,
            PADIN => \N__25207\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__19263\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25200\,
            DIN => \N__25199\,
            DOUT => \N__25198\,
            PACKAGEPIN => \ADV_R_wire\(0)
        );

    \ADV_R_pad_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25200\,
            PADOUT => \N__25199\,
            PADIN => \N__25198\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__16084\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__25191\,
            DIN => \N__25190\,
            DOUT => \N__25189\,
            PACKAGEPIN => DEBUG(2)
        );

    \DEBUG_pad_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25191\,
            PADOUT => \N__25190\,
            PADIN => \N__25189\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__21644\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_VIDEO_pad_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__25182\,
            DIN => \N__25181\,
            DOUT => \N__25180\,
            PACKAGEPIN => \TVP_VIDEO_wire\(3)
        );

    \TVP_VIDEO_pad_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25182\,
            PADOUT => \N__25181\,
            PADIN => \N__25180\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_VIDEO_c_3\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25173\,
            DIN => \N__25172\,
            DOUT => \N__25171\,
            PACKAGEPIN => \ADV_G_wire\(4)
        );

    \ADV_G_pad_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25173\,
            PADOUT => \N__25172\,
            PADIN => \N__25171\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__20969\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25164\,
            DIN => \N__25163\,
            DOUT => \N__25162\,
            PACKAGEPIN => \ADV_R_wire\(5)
        );

    \ADV_R_pad_5_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25164\,
            PADOUT => \N__25163\,
            PADIN => \N__25162\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__21984\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_VIDEO_pad_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__25155\,
            DIN => \N__25154\,
            DOUT => \N__25153\,
            PACKAGEPIN => \TVP_VIDEO_wire\(9)
        );

    \TVP_VIDEO_pad_9_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25155\,
            PADOUT => \N__25154\,
            PADIN => \N__25153\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_VIDEO_c_9\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__25146\,
            DIN => \N__25145\,
            DOUT => \N__25144\,
            PACKAGEPIN => DEBUG(1)
        );

    \DEBUG_pad_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25146\,
            PADOUT => \N__25145\,
            PADIN => \N__25144\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__14426\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_c_6_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__25137\,
            DIN => \N__25136\,
            DOUT => \N__25135\,
            PACKAGEPIN => \TVP_VIDEO_wire\(6)
        );

    \DEBUG_c_6_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25137\,
            PADOUT => \N__25136\,
            PADIN => \N__25135\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DEBUG_c_6_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25128\,
            DIN => \N__25127\,
            DOUT => \N__25126\,
            PACKAGEPIN => \ADV_B_wire\(1)
        );

    \ADV_B_pad_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25128\,
            PADOUT => \N__25127\,
            PADIN => \N__25126\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__20875\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_SYNC_N_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__25119\,
            DIN => \N__25118\,
            DOUT => \N__25117\,
            PACKAGEPIN => \ADV_SYNC_N_wire\
        );

    \ADV_SYNC_N_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25119\,
            PADOUT => \N__25118\,
            PADIN => \N__25117\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25110\,
            DIN => \N__25109\,
            DOUT => \N__25108\,
            PACKAGEPIN => \ADV_B_wire\(6)
        );

    \ADV_B_pad_6_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25110\,
            PADOUT => \N__25109\,
            PADIN => \N__25108\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__23791\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__25101\,
            DIN => \N__25100\,
            DOUT => \N__25099\,
            PACKAGEPIN => DEBUG(6)
        );

    \DEBUG_pad_6_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25101\,
            PADOUT => \N__25100\,
            PADIN => \N__25099\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__14399\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25092\,
            DIN => \N__25091\,
            DOUT => \N__25090\,
            PACKAGEPIN => \ADV_G_wire\(0)
        );

    \ADV_G_pad_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25092\,
            PADOUT => \N__25091\,
            PADIN => \N__25090\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__16085\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25083\,
            DIN => \N__25082\,
            DOUT => \N__25081\,
            PACKAGEPIN => \ADV_R_wire\(1)
        );

    \ADV_R_pad_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25083\,
            PADOUT => \N__25082\,
            PADIN => \N__25081\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__20890\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__25074\,
            DIN => \N__25073\,
            DOUT => \N__25072\,
            PACKAGEPIN => DEBUG(5)
        );

    \DEBUG_pad_5_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25074\,
            PADOUT => \N__25073\,
            PADIN => \N__25072\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__9107\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25065\,
            DIN => \N__25064\,
            DOUT => \N__25063\,
            PACKAGEPIN => \ADV_G_wire\(7)
        );

    \ADV_G_pad_7_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25065\,
            PADOUT => \N__25064\,
            PADIN => \N__25063\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12727\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25056\,
            DIN => \N__25055\,
            DOUT => \N__25054\,
            PACKAGEPIN => \ADV_R_wire\(6)
        );

    \ADV_R_pad_6_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25056\,
            PADOUT => \N__25055\,
            PADIN => \N__25054\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__23795\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_BLANK_N_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__25047\,
            DIN => \N__25046\,
            DOUT => \N__25045\,
            PACKAGEPIN => \ADV_BLANK_N_wire\
        );

    \ADV_BLANK_N_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25047\,
            PADOUT => \N__25046\,
            PADIN => \N__25045\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__24512\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__25038\,
            DIN => \N__25037\,
            DOUT => \N__25036\,
            PACKAGEPIN => DEBUG(0)
        );

    \DEBUG_pad_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25038\,
            PADOUT => \N__25037\,
            PADIN => \N__25036\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__18818\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__25029\,
            DIN => \N__25028\,
            DOUT => \N__25027\,
            PACKAGEPIN => \ADV_B_wire\(2)
        );

    \ADV_B_pad_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25029\,
            PADOUT => \N__25028\,
            PADIN => \N__25027\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__21747\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_c_7_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__25020\,
            DIN => \N__25019\,
            DOUT => \N__25018\,
            PACKAGEPIN => \TVP_VIDEO_wire\(7)
        );

    \DEBUG_c_7_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25020\,
            PADOUT => \N__25019\,
            PADIN => \N__25018\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DEBUG_c_7_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_c_1_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__25011\,
            DIN => \N__25010\,
            DOUT => \N__25009\,
            PACKAGEPIN => \TVP_VSYNC_wire\
        );

    \DEBUG_c_1_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25011\,
            PADOUT => \N__25010\,
            PADIN => \N__25009\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DEBUG_c_1_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_c_5_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__25002\,
            DIN => \N__25001\,
            DOUT => \N__25000\,
            PACKAGEPIN => \TVP_VIDEO_wire\(5)
        );

    \DEBUG_c_5_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__25002\,
            PADOUT => \N__25001\,
            PADIN => \N__25000\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \DEBUG_c_5_c\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24993\,
            DIN => \N__24992\,
            DOUT => \N__24991\,
            PACKAGEPIN => \ADV_B_wire\(7)
        );

    \ADV_B_pad_7_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24993\,
            PADOUT => \N__24992\,
            PADIN => \N__24991\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12726\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LED_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24984\,
            DIN => \N__24983\,
            DOUT => \N__24982\,
            PACKAGEPIN => \LED_wire\
        );

    \LED_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24984\,
            PADOUT => \N__24983\,
            PADIN => \N__24982\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__17495\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_VIDEO_pad_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24975\,
            DIN => \N__24974\,
            DOUT => \N__24973\,
            PACKAGEPIN => \TVP_VIDEO_wire\(4)
        );

    \TVP_VIDEO_pad_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24975\,
            PADOUT => \N__24974\,
            PADIN => \N__24973\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_VIDEO_c_4\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24966\,
            DIN => \N__24965\,
            DOUT => \N__24964\,
            PACKAGEPIN => \ADV_G_wire\(3)
        );

    \ADV_G_pad_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24966\,
            PADOUT => \N__24965\,
            PADIN => \N__24964\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__19268\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_HSYNC_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24957\,
            DIN => \N__24956\,
            DOUT => \N__24955\,
            PACKAGEPIN => \ADV_HSYNC_wire\
        );

    \ADV_HSYNC_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24957\,
            PADOUT => \N__24956\,
            PADIN => \N__24955\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10829\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24948\,
            DIN => \N__24947\,
            DOUT => \N__24946\,
            PACKAGEPIN => \ADV_R_wire\(2)
        );

    \ADV_R_pad_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24948\,
            PADOUT => \N__24947\,
            PADIN => \N__24946\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__21760\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24939\,
            DIN => \N__24938\,
            DOUT => \N__24937\,
            PACKAGEPIN => \ADV_B_wire\(4)
        );

    \ADV_B_pad_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24939\,
            PADOUT => \N__24938\,
            PADIN => \N__24937\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__20964\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24930\,
            DIN => \N__24929\,
            DOUT => \N__24928\,
            PACKAGEPIN => DEBUG(4)
        );

    \DEBUG_pad_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24930\,
            PADOUT => \N__24929\,
            PADIN => \N__24928\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__18767\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24921\,
            DIN => \N__24920\,
            DOUT => \N__24919\,
            PACKAGEPIN => \ADV_G_wire\(6)
        );

    \ADV_G_pad_6_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24921\,
            PADOUT => \N__24920\,
            PADIN => \N__24919\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__23790\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24912\,
            DIN => \N__24911\,
            DOUT => \N__24910\,
            PACKAGEPIN => \ADV_R_wire\(7)
        );

    \ADV_R_pad_7_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24912\,
            PADOUT => \N__24911\,
            PADIN => \N__24910\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12728\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24903\,
            DIN => \N__24902\,
            DOUT => \N__24901\,
            PACKAGEPIN => \ADV_B_wire\(3)
        );

    \ADV_B_pad_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24903\,
            PADOUT => \N__24902\,
            PADIN => \N__24901\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__19264\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_R_pad_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24894\,
            DIN => \N__24893\,
            DOUT => \N__24892\,
            PACKAGEPIN => \ADV_R_wire\(4)
        );

    \ADV_R_pad_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24894\,
            PADOUT => \N__24893\,
            PADIN => \N__24892\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__20965\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \TVP_VIDEO_pad_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24885\,
            DIN => \N__24884\,
            DOUT => \N__24883\,
            PACKAGEPIN => \TVP_VIDEO_wire\(8)
        );

    \TVP_VIDEO_pad_8_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24885\,
            PADOUT => \N__24884\,
            PADIN => \N__24883\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \TVP_VIDEO_c_8\,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24876\,
            DIN => \N__24875\,
            DOUT => \N__24874\,
            PACKAGEPIN => \ADV_B_wire\(0)
        );

    \ADV_B_pad_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24876\,
            PADOUT => \N__24875\,
            PADIN => \N__24874\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__16074\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24867\,
            DIN => \N__24866\,
            DOUT => \N__24865\,
            PACKAGEPIN => \ADV_G_wire\(2)
        );

    \ADV_G_pad_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24867\,
            PADOUT => \N__24866\,
            PADIN => \N__24865\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__21764\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_VSYNC_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24858\,
            DIN => \N__24857\,
            DOUT => \N__24856\,
            PACKAGEPIN => \ADV_VSYNC_wire\
        );

    \ADV_VSYNC_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24858\,
            PADOUT => \N__24857\,
            PADIN => \N__24856\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__19996\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_B_pad_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24849\,
            DIN => \N__24848\,
            DOUT => \N__24847\,
            PACKAGEPIN => \ADV_B_wire\(5)
        );

    \ADV_B_pad_5_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24849\,
            PADOUT => \N__24848\,
            PADIN => \N__24847\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__21995\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \DEBUG_pad_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '1'
        )
    port map (
            OE => \N__24840\,
            DIN => \N__24839\,
            DOUT => \N__24838\,
            PACKAGEPIN => DEBUG(7)
        );

    \DEBUG_pad_7_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24840\,
            PADOUT => \N__24839\,
            PADIN => \N__24838\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__22169\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \ADV_G_pad_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__24831\,
            DIN => \N__24830\,
            DOUT => \N__24829\,
            PACKAGEPIN => \ADV_G_wire\(1)
        );

    \ADV_G_pad_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__24831\,
            PADOUT => \N__24830\,
            PADIN => \N__24829\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__20894\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__6001\ : InMux
    port map (
            O => \N__24812\,
            I => \N__24809\
        );

    \I__6000\ : LocalMux
    port map (
            O => \N__24809\,
            I => \tvp_video_buffer.BUFFER_0_7\
        );

    \I__5999\ : InMux
    port map (
            O => \N__24806\,
            I => \N__24803\
        );

    \I__5998\ : LocalMux
    port map (
            O => \N__24803\,
            I => \tvp_video_buffer.BUFFER_1_7\
        );

    \I__5997\ : InMux
    port map (
            O => \N__24800\,
            I => \N__24790\
        );

    \I__5996\ : InMux
    port map (
            O => \N__24799\,
            I => \N__24787\
        );

    \I__5995\ : InMux
    port map (
            O => \N__24798\,
            I => \N__24781\
        );

    \I__5994\ : InMux
    port map (
            O => \N__24797\,
            I => \N__24776\
        );

    \I__5993\ : InMux
    port map (
            O => \N__24796\,
            I => \N__24773\
        );

    \I__5992\ : InMux
    port map (
            O => \N__24795\,
            I => \N__24769\
        );

    \I__5991\ : InMux
    port map (
            O => \N__24794\,
            I => \N__24766\
        );

    \I__5990\ : InMux
    port map (
            O => \N__24793\,
            I => \N__24760\
        );

    \I__5989\ : LocalMux
    port map (
            O => \N__24790\,
            I => \N__24757\
        );

    \I__5988\ : LocalMux
    port map (
            O => \N__24787\,
            I => \N__24754\
        );

    \I__5987\ : InMux
    port map (
            O => \N__24786\,
            I => \N__24749\
        );

    \I__5986\ : InMux
    port map (
            O => \N__24785\,
            I => \N__24749\
        );

    \I__5985\ : InMux
    port map (
            O => \N__24784\,
            I => \N__24746\
        );

    \I__5984\ : LocalMux
    port map (
            O => \N__24781\,
            I => \N__24740\
        );

    \I__5983\ : InMux
    port map (
            O => \N__24780\,
            I => \N__24737\
        );

    \I__5982\ : InMux
    port map (
            O => \N__24779\,
            I => \N__24734\
        );

    \I__5981\ : LocalMux
    port map (
            O => \N__24776\,
            I => \N__24727\
        );

    \I__5980\ : LocalMux
    port map (
            O => \N__24773\,
            I => \N__24727\
        );

    \I__5979\ : InMux
    port map (
            O => \N__24772\,
            I => \N__24724\
        );

    \I__5978\ : LocalMux
    port map (
            O => \N__24769\,
            I => \N__24719\
        );

    \I__5977\ : LocalMux
    port map (
            O => \N__24766\,
            I => \N__24719\
        );

    \I__5976\ : InMux
    port map (
            O => \N__24765\,
            I => \N__24716\
        );

    \I__5975\ : InMux
    port map (
            O => \N__24764\,
            I => \N__24711\
        );

    \I__5974\ : InMux
    port map (
            O => \N__24763\,
            I => \N__24708\
        );

    \I__5973\ : LocalMux
    port map (
            O => \N__24760\,
            I => \N__24705\
        );

    \I__5972\ : Span4Mux_h
    port map (
            O => \N__24757\,
            I => \N__24696\
        );

    \I__5971\ : Span4Mux_v
    port map (
            O => \N__24754\,
            I => \N__24696\
        );

    \I__5970\ : LocalMux
    port map (
            O => \N__24749\,
            I => \N__24696\
        );

    \I__5969\ : LocalMux
    port map (
            O => \N__24746\,
            I => \N__24696\
        );

    \I__5968\ : InMux
    port map (
            O => \N__24745\,
            I => \N__24693\
        );

    \I__5967\ : InMux
    port map (
            O => \N__24744\,
            I => \N__24690\
        );

    \I__5966\ : InMux
    port map (
            O => \N__24743\,
            I => \N__24687\
        );

    \I__5965\ : Span4Mux_v
    port map (
            O => \N__24740\,
            I => \N__24681\
        );

    \I__5964\ : LocalMux
    port map (
            O => \N__24737\,
            I => \N__24681\
        );

    \I__5963\ : LocalMux
    port map (
            O => \N__24734\,
            I => \N__24678\
        );

    \I__5962\ : InMux
    port map (
            O => \N__24733\,
            I => \N__24675\
        );

    \I__5961\ : InMux
    port map (
            O => \N__24732\,
            I => \N__24672\
        );

    \I__5960\ : Span4Mux_v
    port map (
            O => \N__24727\,
            I => \N__24669\
        );

    \I__5959\ : LocalMux
    port map (
            O => \N__24724\,
            I => \N__24666\
        );

    \I__5958\ : Span4Mux_v
    port map (
            O => \N__24719\,
            I => \N__24663\
        );

    \I__5957\ : LocalMux
    port map (
            O => \N__24716\,
            I => \N__24660\
        );

    \I__5956\ : InMux
    port map (
            O => \N__24715\,
            I => \N__24657\
        );

    \I__5955\ : InMux
    port map (
            O => \N__24714\,
            I => \N__24654\
        );

    \I__5954\ : LocalMux
    port map (
            O => \N__24711\,
            I => \N__24651\
        );

    \I__5953\ : LocalMux
    port map (
            O => \N__24708\,
            I => \N__24642\
        );

    \I__5952\ : Span4Mux_h
    port map (
            O => \N__24705\,
            I => \N__24642\
        );

    \I__5951\ : Span4Mux_v
    port map (
            O => \N__24696\,
            I => \N__24642\
        );

    \I__5950\ : LocalMux
    port map (
            O => \N__24693\,
            I => \N__24642\
        );

    \I__5949\ : LocalMux
    port map (
            O => \N__24690\,
            I => \N__24636\
        );

    \I__5948\ : LocalMux
    port map (
            O => \N__24687\,
            I => \N__24636\
        );

    \I__5947\ : InMux
    port map (
            O => \N__24686\,
            I => \N__24633\
        );

    \I__5946\ : Span4Mux_v
    port map (
            O => \N__24681\,
            I => \N__24630\
        );

    \I__5945\ : Span4Mux_v
    port map (
            O => \N__24678\,
            I => \N__24625\
        );

    \I__5944\ : LocalMux
    port map (
            O => \N__24675\,
            I => \N__24625\
        );

    \I__5943\ : LocalMux
    port map (
            O => \N__24672\,
            I => \N__24618\
        );

    \I__5942\ : Span4Mux_v
    port map (
            O => \N__24669\,
            I => \N__24618\
        );

    \I__5941\ : Span4Mux_v
    port map (
            O => \N__24666\,
            I => \N__24618\
        );

    \I__5940\ : Span4Mux_v
    port map (
            O => \N__24663\,
            I => \N__24613\
        );

    \I__5939\ : Span4Mux_v
    port map (
            O => \N__24660\,
            I => \N__24613\
        );

    \I__5938\ : LocalMux
    port map (
            O => \N__24657\,
            I => \N__24606\
        );

    \I__5937\ : LocalMux
    port map (
            O => \N__24654\,
            I => \N__24606\
        );

    \I__5936\ : Span4Mux_h
    port map (
            O => \N__24651\,
            I => \N__24606\
        );

    \I__5935\ : Span4Mux_h
    port map (
            O => \N__24642\,
            I => \N__24603\
        );

    \I__5934\ : InMux
    port map (
            O => \N__24641\,
            I => \N__24600\
        );

    \I__5933\ : Span12Mux_h
    port map (
            O => \N__24636\,
            I => \N__24597\
        );

    \I__5932\ : LocalMux
    port map (
            O => \N__24633\,
            I => \N__24594\
        );

    \I__5931\ : Span4Mux_v
    port map (
            O => \N__24630\,
            I => \N__24585\
        );

    \I__5930\ : Span4Mux_v
    port map (
            O => \N__24625\,
            I => \N__24585\
        );

    \I__5929\ : Span4Mux_h
    port map (
            O => \N__24618\,
            I => \N__24585\
        );

    \I__5928\ : Span4Mux_h
    port map (
            O => \N__24613\,
            I => \N__24585\
        );

    \I__5927\ : Span4Mux_h
    port map (
            O => \N__24606\,
            I => \N__24582\
        );

    \I__5926\ : Span4Mux_h
    port map (
            O => \N__24603\,
            I => \N__24579\
        );

    \I__5925\ : LocalMux
    port map (
            O => \N__24600\,
            I => \TX_ADDR_11\
        );

    \I__5924\ : Odrv12
    port map (
            O => \N__24597\,
            I => \TX_ADDR_11\
        );

    \I__5923\ : Odrv12
    port map (
            O => \N__24594\,
            I => \TX_ADDR_11\
        );

    \I__5922\ : Odrv4
    port map (
            O => \N__24585\,
            I => \TX_ADDR_11\
        );

    \I__5921\ : Odrv4
    port map (
            O => \N__24582\,
            I => \TX_ADDR_11\
        );

    \I__5920\ : Odrv4
    port map (
            O => \N__24579\,
            I => \TX_ADDR_11\
        );

    \I__5919\ : InMux
    port map (
            O => \N__24566\,
            I => \N__24563\
        );

    \I__5918\ : LocalMux
    port map (
            O => \N__24563\,
            I => \N__24560\
        );

    \I__5917\ : Span4Mux_v
    port map (
            O => \N__24560\,
            I => \N__24557\
        );

    \I__5916\ : Sp12to4
    port map (
            O => \N__24557\,
            I => \N__24554\
        );

    \I__5915\ : Odrv12
    port map (
            O => \N__24554\,
            I => \line_buffer.n538\
        );

    \I__5914\ : InMux
    port map (
            O => \N__24551\,
            I => \N__24548\
        );

    \I__5913\ : LocalMux
    port map (
            O => \N__24548\,
            I => \N__24545\
        );

    \I__5912\ : Span4Mux_v
    port map (
            O => \N__24545\,
            I => \N__24542\
        );

    \I__5911\ : Span4Mux_h
    port map (
            O => \N__24542\,
            I => \N__24539\
        );

    \I__5910\ : Sp12to4
    port map (
            O => \N__24539\,
            I => \N__24536\
        );

    \I__5909\ : Span12Mux_v
    port map (
            O => \N__24536\,
            I => \N__24533\
        );

    \I__5908\ : Odrv12
    port map (
            O => \N__24533\,
            I => \line_buffer.n530\
        );

    \I__5907\ : InMux
    port map (
            O => \N__24530\,
            I => \N__24527\
        );

    \I__5906\ : LocalMux
    port map (
            O => \N__24527\,
            I => \line_buffer.n3542\
        );

    \I__5905\ : SRMux
    port map (
            O => \N__24524\,
            I => \N__24518\
        );

    \I__5904\ : SRMux
    port map (
            O => \N__24523\,
            I => \N__24515\
        );

    \I__5903\ : SRMux
    port map (
            O => \N__24522\,
            I => \N__24509\
        );

    \I__5902\ : SRMux
    port map (
            O => \N__24521\,
            I => \N__24506\
        );

    \I__5901\ : LocalMux
    port map (
            O => \N__24518\,
            I => \N__24500\
        );

    \I__5900\ : LocalMux
    port map (
            O => \N__24515\,
            I => \N__24500\
        );

    \I__5899\ : SRMux
    port map (
            O => \N__24514\,
            I => \N__24497\
        );

    \I__5898\ : IoInMux
    port map (
            O => \N__24513\,
            I => \N__24493\
        );

    \I__5897\ : IoInMux
    port map (
            O => \N__24512\,
            I => \N__24490\
        );

    \I__5896\ : LocalMux
    port map (
            O => \N__24509\,
            I => \N__24485\
        );

    \I__5895\ : LocalMux
    port map (
            O => \N__24506\,
            I => \N__24482\
        );

    \I__5894\ : SRMux
    port map (
            O => \N__24505\,
            I => \N__24479\
        );

    \I__5893\ : Span4Mux_s2_v
    port map (
            O => \N__24500\,
            I => \N__24474\
        );

    \I__5892\ : LocalMux
    port map (
            O => \N__24497\,
            I => \N__24474\
        );

    \I__5891\ : SRMux
    port map (
            O => \N__24496\,
            I => \N__24471\
        );

    \I__5890\ : LocalMux
    port map (
            O => \N__24493\,
            I => \N__24463\
        );

    \I__5889\ : LocalMux
    port map (
            O => \N__24490\,
            I => \N__24463\
        );

    \I__5888\ : SRMux
    port map (
            O => \N__24489\,
            I => \N__24459\
        );

    \I__5887\ : SRMux
    port map (
            O => \N__24488\,
            I => \N__24456\
        );

    \I__5886\ : Span4Mux_v
    port map (
            O => \N__24485\,
            I => \N__24447\
        );

    \I__5885\ : Span4Mux_h
    port map (
            O => \N__24482\,
            I => \N__24447\
        );

    \I__5884\ : LocalMux
    port map (
            O => \N__24479\,
            I => \N__24447\
        );

    \I__5883\ : Span4Mux_v
    port map (
            O => \N__24474\,
            I => \N__24442\
        );

    \I__5882\ : LocalMux
    port map (
            O => \N__24471\,
            I => \N__24442\
        );

    \I__5881\ : SRMux
    port map (
            O => \N__24470\,
            I => \N__24439\
        );

    \I__5880\ : SRMux
    port map (
            O => \N__24469\,
            I => \N__24436\
        );

    \I__5879\ : SRMux
    port map (
            O => \N__24468\,
            I => \N__24432\
        );

    \I__5878\ : IoSpan4Mux
    port map (
            O => \N__24463\,
            I => \N__24429\
        );

    \I__5877\ : SRMux
    port map (
            O => \N__24462\,
            I => \N__24426\
        );

    \I__5876\ : LocalMux
    port map (
            O => \N__24459\,
            I => \N__24419\
        );

    \I__5875\ : LocalMux
    port map (
            O => \N__24456\,
            I => \N__24419\
        );

    \I__5874\ : SRMux
    port map (
            O => \N__24455\,
            I => \N__24416\
        );

    \I__5873\ : SRMux
    port map (
            O => \N__24454\,
            I => \N__24413\
        );

    \I__5872\ : Span4Mux_v
    port map (
            O => \N__24447\,
            I => \N__24404\
        );

    \I__5871\ : Span4Mux_v
    port map (
            O => \N__24442\,
            I => \N__24397\
        );

    \I__5870\ : LocalMux
    port map (
            O => \N__24439\,
            I => \N__24397\
        );

    \I__5869\ : LocalMux
    port map (
            O => \N__24436\,
            I => \N__24397\
        );

    \I__5868\ : SRMux
    port map (
            O => \N__24435\,
            I => \N__24394\
        );

    \I__5867\ : LocalMux
    port map (
            O => \N__24432\,
            I => \N__24391\
        );

    \I__5866\ : IoSpan4Mux
    port map (
            O => \N__24429\,
            I => \N__24388\
        );

    \I__5865\ : LocalMux
    port map (
            O => \N__24426\,
            I => \N__24385\
        );

    \I__5864\ : SRMux
    port map (
            O => \N__24425\,
            I => \N__24382\
        );

    \I__5863\ : SRMux
    port map (
            O => \N__24424\,
            I => \N__24379\
        );

    \I__5862\ : Span4Mux_s2_v
    port map (
            O => \N__24419\,
            I => \N__24370\
        );

    \I__5861\ : LocalMux
    port map (
            O => \N__24416\,
            I => \N__24370\
        );

    \I__5860\ : LocalMux
    port map (
            O => \N__24413\,
            I => \N__24370\
        );

    \I__5859\ : SRMux
    port map (
            O => \N__24412\,
            I => \N__24367\
        );

    \I__5858\ : SRMux
    port map (
            O => \N__24411\,
            I => \N__24364\
        );

    \I__5857\ : SRMux
    port map (
            O => \N__24410\,
            I => \N__24360\
        );

    \I__5856\ : SRMux
    port map (
            O => \N__24409\,
            I => \N__24357\
        );

    \I__5855\ : SRMux
    port map (
            O => \N__24408\,
            I => \N__24354\
        );

    \I__5854\ : SRMux
    port map (
            O => \N__24407\,
            I => \N__24351\
        );

    \I__5853\ : Span4Mux_v
    port map (
            O => \N__24404\,
            I => \N__24344\
        );

    \I__5852\ : Span4Mux_v
    port map (
            O => \N__24397\,
            I => \N__24344\
        );

    \I__5851\ : LocalMux
    port map (
            O => \N__24394\,
            I => \N__24344\
        );

    \I__5850\ : Span4Mux_h
    port map (
            O => \N__24391\,
            I => \N__24339\
        );

    \I__5849\ : Span4Mux_s3_v
    port map (
            O => \N__24388\,
            I => \N__24330\
        );

    \I__5848\ : Span4Mux_s3_v
    port map (
            O => \N__24385\,
            I => \N__24330\
        );

    \I__5847\ : LocalMux
    port map (
            O => \N__24382\,
            I => \N__24330\
        );

    \I__5846\ : LocalMux
    port map (
            O => \N__24379\,
            I => \N__24330\
        );

    \I__5845\ : SRMux
    port map (
            O => \N__24378\,
            I => \N__24327\
        );

    \I__5844\ : SRMux
    port map (
            O => \N__24377\,
            I => \N__24324\
        );

    \I__5843\ : Span4Mux_v
    port map (
            O => \N__24370\,
            I => \N__24315\
        );

    \I__5842\ : LocalMux
    port map (
            O => \N__24367\,
            I => \N__24315\
        );

    \I__5841\ : LocalMux
    port map (
            O => \N__24364\,
            I => \N__24315\
        );

    \I__5840\ : SRMux
    port map (
            O => \N__24363\,
            I => \N__24312\
        );

    \I__5839\ : LocalMux
    port map (
            O => \N__24360\,
            I => \N__24309\
        );

    \I__5838\ : LocalMux
    port map (
            O => \N__24357\,
            I => \N__24306\
        );

    \I__5837\ : LocalMux
    port map (
            O => \N__24354\,
            I => \N__24303\
        );

    \I__5836\ : LocalMux
    port map (
            O => \N__24351\,
            I => \N__24300\
        );

    \I__5835\ : Span4Mux_v
    port map (
            O => \N__24344\,
            I => \N__24297\
        );

    \I__5834\ : SRMux
    port map (
            O => \N__24343\,
            I => \N__24294\
        );

    \I__5833\ : SRMux
    port map (
            O => \N__24342\,
            I => \N__24291\
        );

    \I__5832\ : Span4Mux_h
    port map (
            O => \N__24339\,
            I => \N__24288\
        );

    \I__5831\ : Span4Mux_v
    port map (
            O => \N__24330\,
            I => \N__24281\
        );

    \I__5830\ : LocalMux
    port map (
            O => \N__24327\,
            I => \N__24281\
        );

    \I__5829\ : LocalMux
    port map (
            O => \N__24324\,
            I => \N__24281\
        );

    \I__5828\ : SRMux
    port map (
            O => \N__24323\,
            I => \N__24278\
        );

    \I__5827\ : SRMux
    port map (
            O => \N__24322\,
            I => \N__24275\
        );

    \I__5826\ : Span4Mux_v
    port map (
            O => \N__24315\,
            I => \N__24270\
        );

    \I__5825\ : LocalMux
    port map (
            O => \N__24312\,
            I => \N__24270\
        );

    \I__5824\ : Span12Mux_s9_h
    port map (
            O => \N__24309\,
            I => \N__24266\
        );

    \I__5823\ : Span12Mux_s9_h
    port map (
            O => \N__24306\,
            I => \N__24263\
        );

    \I__5822\ : Span12Mux_h
    port map (
            O => \N__24303\,
            I => \N__24260\
        );

    \I__5821\ : Span12Mux_h
    port map (
            O => \N__24300\,
            I => \N__24257\
        );

    \I__5820\ : Sp12to4
    port map (
            O => \N__24297\,
            I => \N__24252\
        );

    \I__5819\ : LocalMux
    port map (
            O => \N__24294\,
            I => \N__24252\
        );

    \I__5818\ : LocalMux
    port map (
            O => \N__24291\,
            I => \N__24249\
        );

    \I__5817\ : Span4Mux_h
    port map (
            O => \N__24288\,
            I => \N__24246\
        );

    \I__5816\ : Span4Mux_v
    port map (
            O => \N__24281\,
            I => \N__24241\
        );

    \I__5815\ : LocalMux
    port map (
            O => \N__24278\,
            I => \N__24241\
        );

    \I__5814\ : LocalMux
    port map (
            O => \N__24275\,
            I => \N__24238\
        );

    \I__5813\ : Span4Mux_v
    port map (
            O => \N__24270\,
            I => \N__24235\
        );

    \I__5812\ : SRMux
    port map (
            O => \N__24269\,
            I => \N__24232\
        );

    \I__5811\ : Span12Mux_h
    port map (
            O => \N__24266\,
            I => \N__24227\
        );

    \I__5810\ : Span12Mux_h
    port map (
            O => \N__24263\,
            I => \N__24227\
        );

    \I__5809\ : Span12Mux_v
    port map (
            O => \N__24260\,
            I => \N__24220\
        );

    \I__5808\ : Span12Mux_v
    port map (
            O => \N__24257\,
            I => \N__24220\
        );

    \I__5807\ : Span12Mux_h
    port map (
            O => \N__24252\,
            I => \N__24220\
        );

    \I__5806\ : Span4Mux_h
    port map (
            O => \N__24249\,
            I => \N__24217\
        );

    \I__5805\ : Span4Mux_h
    port map (
            O => \N__24246\,
            I => \N__24210\
        );

    \I__5804\ : Span4Mux_h
    port map (
            O => \N__24241\,
            I => \N__24210\
        );

    \I__5803\ : Span4Mux_h
    port map (
            O => \N__24238\,
            I => \N__24210\
        );

    \I__5802\ : Span4Mux_v
    port map (
            O => \N__24235\,
            I => \N__24205\
        );

    \I__5801\ : LocalMux
    port map (
            O => \N__24232\,
            I => \N__24205\
        );

    \I__5800\ : Odrv12
    port map (
            O => \N__24227\,
            I => \CONSTANT_ONE_NET\
        );

    \I__5799\ : Odrv12
    port map (
            O => \N__24220\,
            I => \CONSTANT_ONE_NET\
        );

    \I__5798\ : Odrv4
    port map (
            O => \N__24217\,
            I => \CONSTANT_ONE_NET\
        );

    \I__5797\ : Odrv4
    port map (
            O => \N__24210\,
            I => \CONSTANT_ONE_NET\
        );

    \I__5796\ : Odrv4
    port map (
            O => \N__24205\,
            I => \CONSTANT_ONE_NET\
        );

    \I__5795\ : InMux
    port map (
            O => \N__24194\,
            I => \N__24191\
        );

    \I__5794\ : LocalMux
    port map (
            O => \N__24191\,
            I => \N__24188\
        );

    \I__5793\ : Odrv12
    port map (
            O => \N__24188\,
            I => \TVP_VIDEO_c_9\
        );

    \I__5792\ : InMux
    port map (
            O => \N__24185\,
            I => \N__24182\
        );

    \I__5791\ : LocalMux
    port map (
            O => \N__24182\,
            I => \N__24179\
        );

    \I__5790\ : Span4Mux_v
    port map (
            O => \N__24179\,
            I => \N__24176\
        );

    \I__5789\ : Odrv4
    port map (
            O => \N__24176\,
            I => \tvp_video_buffer.BUFFER_0_9\
        );

    \I__5788\ : InMux
    port map (
            O => \N__24173\,
            I => \N__24170\
        );

    \I__5787\ : LocalMux
    port map (
            O => \N__24170\,
            I => \N__24149\
        );

    \I__5786\ : ClkMux
    port map (
            O => \N__24169\,
            I => \N__23957\
        );

    \I__5785\ : ClkMux
    port map (
            O => \N__24168\,
            I => \N__23957\
        );

    \I__5784\ : ClkMux
    port map (
            O => \N__24167\,
            I => \N__23957\
        );

    \I__5783\ : ClkMux
    port map (
            O => \N__24166\,
            I => \N__23957\
        );

    \I__5782\ : ClkMux
    port map (
            O => \N__24165\,
            I => \N__23957\
        );

    \I__5781\ : ClkMux
    port map (
            O => \N__24164\,
            I => \N__23957\
        );

    \I__5780\ : ClkMux
    port map (
            O => \N__24163\,
            I => \N__23957\
        );

    \I__5779\ : ClkMux
    port map (
            O => \N__24162\,
            I => \N__23957\
        );

    \I__5778\ : ClkMux
    port map (
            O => \N__24161\,
            I => \N__23957\
        );

    \I__5777\ : ClkMux
    port map (
            O => \N__24160\,
            I => \N__23957\
        );

    \I__5776\ : ClkMux
    port map (
            O => \N__24159\,
            I => \N__23957\
        );

    \I__5775\ : ClkMux
    port map (
            O => \N__24158\,
            I => \N__23957\
        );

    \I__5774\ : ClkMux
    port map (
            O => \N__24157\,
            I => \N__23957\
        );

    \I__5773\ : ClkMux
    port map (
            O => \N__24156\,
            I => \N__23957\
        );

    \I__5772\ : ClkMux
    port map (
            O => \N__24155\,
            I => \N__23957\
        );

    \I__5771\ : ClkMux
    port map (
            O => \N__24154\,
            I => \N__23957\
        );

    \I__5770\ : ClkMux
    port map (
            O => \N__24153\,
            I => \N__23957\
        );

    \I__5769\ : ClkMux
    port map (
            O => \N__24152\,
            I => \N__23957\
        );

    \I__5768\ : Glb2LocalMux
    port map (
            O => \N__24149\,
            I => \N__23957\
        );

    \I__5767\ : ClkMux
    port map (
            O => \N__24148\,
            I => \N__23957\
        );

    \I__5766\ : ClkMux
    port map (
            O => \N__24147\,
            I => \N__23957\
        );

    \I__5765\ : ClkMux
    port map (
            O => \N__24146\,
            I => \N__23957\
        );

    \I__5764\ : ClkMux
    port map (
            O => \N__24145\,
            I => \N__23957\
        );

    \I__5763\ : ClkMux
    port map (
            O => \N__24144\,
            I => \N__23957\
        );

    \I__5762\ : ClkMux
    port map (
            O => \N__24143\,
            I => \N__23957\
        );

    \I__5761\ : ClkMux
    port map (
            O => \N__24142\,
            I => \N__23957\
        );

    \I__5760\ : ClkMux
    port map (
            O => \N__24141\,
            I => \N__23957\
        );

    \I__5759\ : ClkMux
    port map (
            O => \N__24140\,
            I => \N__23957\
        );

    \I__5758\ : ClkMux
    port map (
            O => \N__24139\,
            I => \N__23957\
        );

    \I__5757\ : ClkMux
    port map (
            O => \N__24138\,
            I => \N__23957\
        );

    \I__5756\ : ClkMux
    port map (
            O => \N__24137\,
            I => \N__23957\
        );

    \I__5755\ : ClkMux
    port map (
            O => \N__24136\,
            I => \N__23957\
        );

    \I__5754\ : ClkMux
    port map (
            O => \N__24135\,
            I => \N__23957\
        );

    \I__5753\ : ClkMux
    port map (
            O => \N__24134\,
            I => \N__23957\
        );

    \I__5752\ : ClkMux
    port map (
            O => \N__24133\,
            I => \N__23957\
        );

    \I__5751\ : ClkMux
    port map (
            O => \N__24132\,
            I => \N__23957\
        );

    \I__5750\ : ClkMux
    port map (
            O => \N__24131\,
            I => \N__23957\
        );

    \I__5749\ : ClkMux
    port map (
            O => \N__24130\,
            I => \N__23957\
        );

    \I__5748\ : ClkMux
    port map (
            O => \N__24129\,
            I => \N__23957\
        );

    \I__5747\ : ClkMux
    port map (
            O => \N__24128\,
            I => \N__23957\
        );

    \I__5746\ : ClkMux
    port map (
            O => \N__24127\,
            I => \N__23957\
        );

    \I__5745\ : ClkMux
    port map (
            O => \N__24126\,
            I => \N__23957\
        );

    \I__5744\ : ClkMux
    port map (
            O => \N__24125\,
            I => \N__23957\
        );

    \I__5743\ : ClkMux
    port map (
            O => \N__24124\,
            I => \N__23957\
        );

    \I__5742\ : ClkMux
    port map (
            O => \N__24123\,
            I => \N__23957\
        );

    \I__5741\ : ClkMux
    port map (
            O => \N__24122\,
            I => \N__23957\
        );

    \I__5740\ : ClkMux
    port map (
            O => \N__24121\,
            I => \N__23957\
        );

    \I__5739\ : ClkMux
    port map (
            O => \N__24120\,
            I => \N__23957\
        );

    \I__5738\ : ClkMux
    port map (
            O => \N__24119\,
            I => \N__23957\
        );

    \I__5737\ : ClkMux
    port map (
            O => \N__24118\,
            I => \N__23957\
        );

    \I__5736\ : ClkMux
    port map (
            O => \N__24117\,
            I => \N__23957\
        );

    \I__5735\ : ClkMux
    port map (
            O => \N__24116\,
            I => \N__23957\
        );

    \I__5734\ : ClkMux
    port map (
            O => \N__24115\,
            I => \N__23957\
        );

    \I__5733\ : ClkMux
    port map (
            O => \N__24114\,
            I => \N__23957\
        );

    \I__5732\ : ClkMux
    port map (
            O => \N__24113\,
            I => \N__23957\
        );

    \I__5731\ : ClkMux
    port map (
            O => \N__24112\,
            I => \N__23957\
        );

    \I__5730\ : ClkMux
    port map (
            O => \N__24111\,
            I => \N__23957\
        );

    \I__5729\ : ClkMux
    port map (
            O => \N__24110\,
            I => \N__23957\
        );

    \I__5728\ : ClkMux
    port map (
            O => \N__24109\,
            I => \N__23957\
        );

    \I__5727\ : ClkMux
    port map (
            O => \N__24108\,
            I => \N__23957\
        );

    \I__5726\ : ClkMux
    port map (
            O => \N__24107\,
            I => \N__23957\
        );

    \I__5725\ : ClkMux
    port map (
            O => \N__24106\,
            I => \N__23957\
        );

    \I__5724\ : ClkMux
    port map (
            O => \N__24105\,
            I => \N__23957\
        );

    \I__5723\ : ClkMux
    port map (
            O => \N__24104\,
            I => \N__23957\
        );

    \I__5722\ : ClkMux
    port map (
            O => \N__24103\,
            I => \N__23957\
        );

    \I__5721\ : ClkMux
    port map (
            O => \N__24102\,
            I => \N__23957\
        );

    \I__5720\ : ClkMux
    port map (
            O => \N__24101\,
            I => \N__23957\
        );

    \I__5719\ : ClkMux
    port map (
            O => \N__24100\,
            I => \N__23957\
        );

    \I__5718\ : ClkMux
    port map (
            O => \N__24099\,
            I => \N__23957\
        );

    \I__5717\ : ClkMux
    port map (
            O => \N__24098\,
            I => \N__23957\
        );

    \I__5716\ : GlobalMux
    port map (
            O => \N__23957\,
            I => \N__23954\
        );

    \I__5715\ : gio2CtrlBuf
    port map (
            O => \N__23954\,
            I => \DEBUG_c_3_c\
        );

    \I__5714\ : CascadeMux
    port map (
            O => \N__23951\,
            I => \N__23945\
        );

    \I__5713\ : CascadeMux
    port map (
            O => \N__23950\,
            I => \N__23941\
        );

    \I__5712\ : CascadeMux
    port map (
            O => \N__23949\,
            I => \N__23934\
        );

    \I__5711\ : InMux
    port map (
            O => \N__23948\,
            I => \N__23929\
        );

    \I__5710\ : InMux
    port map (
            O => \N__23945\,
            I => \N__23926\
        );

    \I__5709\ : InMux
    port map (
            O => \N__23944\,
            I => \N__23923\
        );

    \I__5708\ : InMux
    port map (
            O => \N__23941\,
            I => \N__23920\
        );

    \I__5707\ : InMux
    port map (
            O => \N__23940\,
            I => \N__23914\
        );

    \I__5706\ : InMux
    port map (
            O => \N__23939\,
            I => \N__23911\
        );

    \I__5705\ : InMux
    port map (
            O => \N__23938\,
            I => \N__23908\
        );

    \I__5704\ : InMux
    port map (
            O => \N__23937\,
            I => \N__23905\
        );

    \I__5703\ : InMux
    port map (
            O => \N__23934\,
            I => \N__23902\
        );

    \I__5702\ : CascadeMux
    port map (
            O => \N__23933\,
            I => \N__23899\
        );

    \I__5701\ : InMux
    port map (
            O => \N__23932\,
            I => \N__23896\
        );

    \I__5700\ : LocalMux
    port map (
            O => \N__23929\,
            I => \N__23891\
        );

    \I__5699\ : LocalMux
    port map (
            O => \N__23926\,
            I => \N__23891\
        );

    \I__5698\ : LocalMux
    port map (
            O => \N__23923\,
            I => \N__23886\
        );

    \I__5697\ : LocalMux
    port map (
            O => \N__23920\,
            I => \N__23886\
        );

    \I__5696\ : CascadeMux
    port map (
            O => \N__23919\,
            I => \N__23883\
        );

    \I__5695\ : InMux
    port map (
            O => \N__23918\,
            I => \N__23880\
        );

    \I__5694\ : InMux
    port map (
            O => \N__23917\,
            I => \N__23877\
        );

    \I__5693\ : LocalMux
    port map (
            O => \N__23914\,
            I => \N__23874\
        );

    \I__5692\ : LocalMux
    port map (
            O => \N__23911\,
            I => \N__23871\
        );

    \I__5691\ : LocalMux
    port map (
            O => \N__23908\,
            I => \N__23864\
        );

    \I__5690\ : LocalMux
    port map (
            O => \N__23905\,
            I => \N__23864\
        );

    \I__5689\ : LocalMux
    port map (
            O => \N__23902\,
            I => \N__23864\
        );

    \I__5688\ : InMux
    port map (
            O => \N__23899\,
            I => \N__23861\
        );

    \I__5687\ : LocalMux
    port map (
            O => \N__23896\,
            I => \N__23856\
        );

    \I__5686\ : Span4Mux_h
    port map (
            O => \N__23891\,
            I => \N__23856\
        );

    \I__5685\ : Span4Mux_h
    port map (
            O => \N__23886\,
            I => \N__23853\
        );

    \I__5684\ : InMux
    port map (
            O => \N__23883\,
            I => \N__23850\
        );

    \I__5683\ : LocalMux
    port map (
            O => \N__23880\,
            I => \N__23847\
        );

    \I__5682\ : LocalMux
    port map (
            O => \N__23877\,
            I => \N__23844\
        );

    \I__5681\ : Span4Mux_v
    port map (
            O => \N__23874\,
            I => \N__23839\
        );

    \I__5680\ : Span4Mux_h
    port map (
            O => \N__23871\,
            I => \N__23839\
        );

    \I__5679\ : Span12Mux_h
    port map (
            O => \N__23864\,
            I => \N__23836\
        );

    \I__5678\ : LocalMux
    port map (
            O => \N__23861\,
            I => \N__23827\
        );

    \I__5677\ : Span4Mux_h
    port map (
            O => \N__23856\,
            I => \N__23827\
        );

    \I__5676\ : Span4Mux_h
    port map (
            O => \N__23853\,
            I => \N__23827\
        );

    \I__5675\ : LocalMux
    port map (
            O => \N__23850\,
            I => \N__23827\
        );

    \I__5674\ : Span4Mux_h
    port map (
            O => \N__23847\,
            I => \N__23822\
        );

    \I__5673\ : Span4Mux_h
    port map (
            O => \N__23844\,
            I => \N__23822\
        );

    \I__5672\ : Odrv4
    port map (
            O => \N__23839\,
            I => \TX_ADDR_13\
        );

    \I__5671\ : Odrv12
    port map (
            O => \N__23836\,
            I => \TX_ADDR_13\
        );

    \I__5670\ : Odrv4
    port map (
            O => \N__23827\,
            I => \TX_ADDR_13\
        );

    \I__5669\ : Odrv4
    port map (
            O => \N__23822\,
            I => \TX_ADDR_13\
        );

    \I__5668\ : CascadeMux
    port map (
            O => \N__23813\,
            I => \line_buffer.n3608_cascade_\
        );

    \I__5667\ : InMux
    port map (
            O => \N__23810\,
            I => \N__23807\
        );

    \I__5666\ : LocalMux
    port map (
            O => \N__23807\,
            I => \N__23804\
        );

    \I__5665\ : Odrv4
    port map (
            O => \N__23804\,
            I => \line_buffer.n3576\
        );

    \I__5664\ : InMux
    port map (
            O => \N__23801\,
            I => \N__23798\
        );

    \I__5663\ : LocalMux
    port map (
            O => \N__23798\,
            I => \TX_DATA_6\
        );

    \I__5662\ : IoInMux
    port map (
            O => \N__23795\,
            I => \N__23792\
        );

    \I__5661\ : LocalMux
    port map (
            O => \N__23792\,
            I => \N__23787\
        );

    \I__5660\ : IoInMux
    port map (
            O => \N__23791\,
            I => \N__23784\
        );

    \I__5659\ : IoInMux
    port map (
            O => \N__23790\,
            I => \N__23781\
        );

    \I__5658\ : Span4Mux_s3_h
    port map (
            O => \N__23787\,
            I => \N__23778\
        );

    \I__5657\ : LocalMux
    port map (
            O => \N__23784\,
            I => \N__23775\
        );

    \I__5656\ : LocalMux
    port map (
            O => \N__23781\,
            I => \N__23772\
        );

    \I__5655\ : Span4Mux_v
    port map (
            O => \N__23778\,
            I => \N__23769\
        );

    \I__5654\ : Span4Mux_s3_v
    port map (
            O => \N__23775\,
            I => \N__23766\
        );

    \I__5653\ : IoSpan4Mux
    port map (
            O => \N__23772\,
            I => \N__23763\
        );

    \I__5652\ : Span4Mux_v
    port map (
            O => \N__23769\,
            I => \N__23760\
        );

    \I__5651\ : Span4Mux_h
    port map (
            O => \N__23766\,
            I => \N__23757\
        );

    \I__5650\ : Span4Mux_s3_v
    port map (
            O => \N__23763\,
            I => \N__23754\
        );

    \I__5649\ : Sp12to4
    port map (
            O => \N__23760\,
            I => \N__23751\
        );

    \I__5648\ : Sp12to4
    port map (
            O => \N__23757\,
            I => \N__23748\
        );

    \I__5647\ : Sp12to4
    port map (
            O => \N__23754\,
            I => \N__23745\
        );

    \I__5646\ : Span12Mux_h
    port map (
            O => \N__23751\,
            I => \N__23738\
        );

    \I__5645\ : Span12Mux_s10_v
    port map (
            O => \N__23748\,
            I => \N__23738\
        );

    \I__5644\ : Span12Mux_s10_v
    port map (
            O => \N__23745\,
            I => \N__23738\
        );

    \I__5643\ : Odrv12
    port map (
            O => \N__23738\,
            I => n1815
        );

    \I__5642\ : ClkMux
    port map (
            O => \N__23735\,
            I => \N__23731\
        );

    \I__5641\ : ClkMux
    port map (
            O => \N__23734\,
            I => \N__23725\
        );

    \I__5640\ : LocalMux
    port map (
            O => \N__23731\,
            I => \N__23719\
        );

    \I__5639\ : ClkMux
    port map (
            O => \N__23730\,
            I => \N__23716\
        );

    \I__5638\ : ClkMux
    port map (
            O => \N__23729\,
            I => \N__23711\
        );

    \I__5637\ : ClkMux
    port map (
            O => \N__23728\,
            I => \N__23705\
        );

    \I__5636\ : LocalMux
    port map (
            O => \N__23725\,
            I => \N__23700\
        );

    \I__5635\ : ClkMux
    port map (
            O => \N__23724\,
            I => \N__23697\
        );

    \I__5634\ : ClkMux
    port map (
            O => \N__23723\,
            I => \N__23693\
        );

    \I__5633\ : ClkMux
    port map (
            O => \N__23722\,
            I => \N__23690\
        );

    \I__5632\ : Span4Mux_s2_v
    port map (
            O => \N__23719\,
            I => \N__23681\
        );

    \I__5631\ : LocalMux
    port map (
            O => \N__23716\,
            I => \N__23681\
        );

    \I__5630\ : ClkMux
    port map (
            O => \N__23715\,
            I => \N__23678\
        );

    \I__5629\ : ClkMux
    port map (
            O => \N__23714\,
            I => \N__23674\
        );

    \I__5628\ : LocalMux
    port map (
            O => \N__23711\,
            I => \N__23671\
        );

    \I__5627\ : ClkMux
    port map (
            O => \N__23710\,
            I => \N__23668\
        );

    \I__5626\ : ClkMux
    port map (
            O => \N__23709\,
            I => \N__23663\
        );

    \I__5625\ : ClkMux
    port map (
            O => \N__23708\,
            I => \N__23660\
        );

    \I__5624\ : LocalMux
    port map (
            O => \N__23705\,
            I => \N__23657\
        );

    \I__5623\ : ClkMux
    port map (
            O => \N__23704\,
            I => \N__23653\
        );

    \I__5622\ : ClkMux
    port map (
            O => \N__23703\,
            I => \N__23650\
        );

    \I__5621\ : Span4Mux_v
    port map (
            O => \N__23700\,
            I => \N__23641\
        );

    \I__5620\ : LocalMux
    port map (
            O => \N__23697\,
            I => \N__23641\
        );

    \I__5619\ : ClkMux
    port map (
            O => \N__23696\,
            I => \N__23638\
        );

    \I__5618\ : LocalMux
    port map (
            O => \N__23693\,
            I => \N__23631\
        );

    \I__5617\ : LocalMux
    port map (
            O => \N__23690\,
            I => \N__23628\
        );

    \I__5616\ : ClkMux
    port map (
            O => \N__23689\,
            I => \N__23625\
        );

    \I__5615\ : ClkMux
    port map (
            O => \N__23688\,
            I => \N__23622\
        );

    \I__5614\ : ClkMux
    port map (
            O => \N__23687\,
            I => \N__23617\
        );

    \I__5613\ : ClkMux
    port map (
            O => \N__23686\,
            I => \N__23614\
        );

    \I__5612\ : Span4Mux_v
    port map (
            O => \N__23681\,
            I => \N__23608\
        );

    \I__5611\ : LocalMux
    port map (
            O => \N__23678\,
            I => \N__23608\
        );

    \I__5610\ : ClkMux
    port map (
            O => \N__23677\,
            I => \N__23605\
        );

    \I__5609\ : LocalMux
    port map (
            O => \N__23674\,
            I => \N__23595\
        );

    \I__5608\ : Span4Mux_h
    port map (
            O => \N__23671\,
            I => \N__23590\
        );

    \I__5607\ : LocalMux
    port map (
            O => \N__23668\,
            I => \N__23590\
        );

    \I__5606\ : ClkMux
    port map (
            O => \N__23667\,
            I => \N__23587\
        );

    \I__5605\ : ClkMux
    port map (
            O => \N__23666\,
            I => \N__23584\
        );

    \I__5604\ : LocalMux
    port map (
            O => \N__23663\,
            I => \N__23581\
        );

    \I__5603\ : LocalMux
    port map (
            O => \N__23660\,
            I => \N__23578\
        );

    \I__5602\ : Span4Mux_h
    port map (
            O => \N__23657\,
            I => \N__23575\
        );

    \I__5601\ : ClkMux
    port map (
            O => \N__23656\,
            I => \N__23572\
        );

    \I__5600\ : LocalMux
    port map (
            O => \N__23653\,
            I => \N__23567\
        );

    \I__5599\ : LocalMux
    port map (
            O => \N__23650\,
            I => \N__23564\
        );

    \I__5598\ : ClkMux
    port map (
            O => \N__23649\,
            I => \N__23561\
        );

    \I__5597\ : ClkMux
    port map (
            O => \N__23648\,
            I => \N__23557\
        );

    \I__5596\ : ClkMux
    port map (
            O => \N__23647\,
            I => \N__23554\
        );

    \I__5595\ : ClkMux
    port map (
            O => \N__23646\,
            I => \N__23547\
        );

    \I__5594\ : Span4Mux_v
    port map (
            O => \N__23641\,
            I => \N__23542\
        );

    \I__5593\ : LocalMux
    port map (
            O => \N__23638\,
            I => \N__23542\
        );

    \I__5592\ : ClkMux
    port map (
            O => \N__23637\,
            I => \N__23539\
        );

    \I__5591\ : ClkMux
    port map (
            O => \N__23636\,
            I => \N__23536\
        );

    \I__5590\ : ClkMux
    port map (
            O => \N__23635\,
            I => \N__23533\
        );

    \I__5589\ : ClkMux
    port map (
            O => \N__23634\,
            I => \N__23528\
        );

    \I__5588\ : Span4Mux_s2_v
    port map (
            O => \N__23631\,
            I => \N__23520\
        );

    \I__5587\ : Span4Mux_h
    port map (
            O => \N__23628\,
            I => \N__23520\
        );

    \I__5586\ : LocalMux
    port map (
            O => \N__23625\,
            I => \N__23520\
        );

    \I__5585\ : LocalMux
    port map (
            O => \N__23622\,
            I => \N__23517\
        );

    \I__5584\ : ClkMux
    port map (
            O => \N__23621\,
            I => \N__23514\
        );

    \I__5583\ : ClkMux
    port map (
            O => \N__23620\,
            I => \N__23511\
        );

    \I__5582\ : LocalMux
    port map (
            O => \N__23617\,
            I => \N__23506\
        );

    \I__5581\ : LocalMux
    port map (
            O => \N__23614\,
            I => \N__23503\
        );

    \I__5580\ : ClkMux
    port map (
            O => \N__23613\,
            I => \N__23500\
        );

    \I__5579\ : Span4Mux_v
    port map (
            O => \N__23608\,
            I => \N__23495\
        );

    \I__5578\ : LocalMux
    port map (
            O => \N__23605\,
            I => \N__23495\
        );

    \I__5577\ : ClkMux
    port map (
            O => \N__23604\,
            I => \N__23492\
        );

    \I__5576\ : ClkMux
    port map (
            O => \N__23603\,
            I => \N__23489\
        );

    \I__5575\ : ClkMux
    port map (
            O => \N__23602\,
            I => \N__23483\
        );

    \I__5574\ : ClkMux
    port map (
            O => \N__23601\,
            I => \N__23479\
        );

    \I__5573\ : ClkMux
    port map (
            O => \N__23600\,
            I => \N__23475\
        );

    \I__5572\ : ClkMux
    port map (
            O => \N__23599\,
            I => \N__23471\
        );

    \I__5571\ : ClkMux
    port map (
            O => \N__23598\,
            I => \N__23468\
        );

    \I__5570\ : Span4Mux_h
    port map (
            O => \N__23595\,
            I => \N__23457\
        );

    \I__5569\ : Span4Mux_h
    port map (
            O => \N__23590\,
            I => \N__23457\
        );

    \I__5568\ : LocalMux
    port map (
            O => \N__23587\,
            I => \N__23457\
        );

    \I__5567\ : LocalMux
    port map (
            O => \N__23584\,
            I => \N__23457\
        );

    \I__5566\ : Span4Mux_v
    port map (
            O => \N__23581\,
            I => \N__23452\
        );

    \I__5565\ : Span4Mux_h
    port map (
            O => \N__23578\,
            I => \N__23452\
        );

    \I__5564\ : Span4Mux_v
    port map (
            O => \N__23575\,
            I => \N__23447\
        );

    \I__5563\ : LocalMux
    port map (
            O => \N__23572\,
            I => \N__23447\
        );

    \I__5562\ : ClkMux
    port map (
            O => \N__23571\,
            I => \N__23444\
        );

    \I__5561\ : ClkMux
    port map (
            O => \N__23570\,
            I => \N__23441\
        );

    \I__5560\ : Span4Mux_h
    port map (
            O => \N__23567\,
            I => \N__23436\
        );

    \I__5559\ : Span4Mux_v
    port map (
            O => \N__23564\,
            I => \N__23431\
        );

    \I__5558\ : LocalMux
    port map (
            O => \N__23561\,
            I => \N__23431\
        );

    \I__5557\ : ClkMux
    port map (
            O => \N__23560\,
            I => \N__23428\
        );

    \I__5556\ : LocalMux
    port map (
            O => \N__23557\,
            I => \N__23425\
        );

    \I__5555\ : LocalMux
    port map (
            O => \N__23554\,
            I => \N__23422\
        );

    \I__5554\ : ClkMux
    port map (
            O => \N__23553\,
            I => \N__23419\
        );

    \I__5553\ : ClkMux
    port map (
            O => \N__23552\,
            I => \N__23414\
        );

    \I__5552\ : ClkMux
    port map (
            O => \N__23551\,
            I => \N__23410\
        );

    \I__5551\ : ClkMux
    port map (
            O => \N__23550\,
            I => \N__23406\
        );

    \I__5550\ : LocalMux
    port map (
            O => \N__23547\,
            I => \N__23400\
        );

    \I__5549\ : Span4Mux_h
    port map (
            O => \N__23542\,
            I => \N__23395\
        );

    \I__5548\ : LocalMux
    port map (
            O => \N__23539\,
            I => \N__23395\
        );

    \I__5547\ : LocalMux
    port map (
            O => \N__23536\,
            I => \N__23390\
        );

    \I__5546\ : LocalMux
    port map (
            O => \N__23533\,
            I => \N__23390\
        );

    \I__5545\ : ClkMux
    port map (
            O => \N__23532\,
            I => \N__23387\
        );

    \I__5544\ : ClkMux
    port map (
            O => \N__23531\,
            I => \N__23384\
        );

    \I__5543\ : LocalMux
    port map (
            O => \N__23528\,
            I => \N__23380\
        );

    \I__5542\ : ClkMux
    port map (
            O => \N__23527\,
            I => \N__23377\
        );

    \I__5541\ : Span4Mux_v
    port map (
            O => \N__23520\,
            I => \N__23368\
        );

    \I__5540\ : Span4Mux_h
    port map (
            O => \N__23517\,
            I => \N__23368\
        );

    \I__5539\ : LocalMux
    port map (
            O => \N__23514\,
            I => \N__23368\
        );

    \I__5538\ : LocalMux
    port map (
            O => \N__23511\,
            I => \N__23365\
        );

    \I__5537\ : ClkMux
    port map (
            O => \N__23510\,
            I => \N__23362\
        );

    \I__5536\ : ClkMux
    port map (
            O => \N__23509\,
            I => \N__23359\
        );

    \I__5535\ : Span4Mux_v
    port map (
            O => \N__23506\,
            I => \N__23350\
        );

    \I__5534\ : Span4Mux_h
    port map (
            O => \N__23503\,
            I => \N__23350\
        );

    \I__5533\ : LocalMux
    port map (
            O => \N__23500\,
            I => \N__23350\
        );

    \I__5532\ : Span4Mux_h
    port map (
            O => \N__23495\,
            I => \N__23343\
        );

    \I__5531\ : LocalMux
    port map (
            O => \N__23492\,
            I => \N__23343\
        );

    \I__5530\ : LocalMux
    port map (
            O => \N__23489\,
            I => \N__23343\
        );

    \I__5529\ : ClkMux
    port map (
            O => \N__23488\,
            I => \N__23340\
        );

    \I__5528\ : ClkMux
    port map (
            O => \N__23487\,
            I => \N__23337\
        );

    \I__5527\ : ClkMux
    port map (
            O => \N__23486\,
            I => \N__23332\
        );

    \I__5526\ : LocalMux
    port map (
            O => \N__23483\,
            I => \N__23328\
        );

    \I__5525\ : ClkMux
    port map (
            O => \N__23482\,
            I => \N__23325\
        );

    \I__5524\ : LocalMux
    port map (
            O => \N__23479\,
            I => \N__23321\
        );

    \I__5523\ : ClkMux
    port map (
            O => \N__23478\,
            I => \N__23318\
        );

    \I__5522\ : LocalMux
    port map (
            O => \N__23475\,
            I => \N__23315\
        );

    \I__5521\ : ClkMux
    port map (
            O => \N__23474\,
            I => \N__23312\
        );

    \I__5520\ : LocalMux
    port map (
            O => \N__23471\,
            I => \N__23309\
        );

    \I__5519\ : LocalMux
    port map (
            O => \N__23468\,
            I => \N__23306\
        );

    \I__5518\ : ClkMux
    port map (
            O => \N__23467\,
            I => \N__23303\
        );

    \I__5517\ : ClkMux
    port map (
            O => \N__23466\,
            I => \N__23299\
        );

    \I__5516\ : Span4Mux_h
    port map (
            O => \N__23457\,
            I => \N__23295\
        );

    \I__5515\ : Span4Mux_h
    port map (
            O => \N__23452\,
            I => \N__23288\
        );

    \I__5514\ : Span4Mux_v
    port map (
            O => \N__23447\,
            I => \N__23288\
        );

    \I__5513\ : LocalMux
    port map (
            O => \N__23444\,
            I => \N__23288\
        );

    \I__5512\ : LocalMux
    port map (
            O => \N__23441\,
            I => \N__23285\
        );

    \I__5511\ : ClkMux
    port map (
            O => \N__23440\,
            I => \N__23282\
        );

    \I__5510\ : ClkMux
    port map (
            O => \N__23439\,
            I => \N__23279\
        );

    \I__5509\ : Span4Mux_v
    port map (
            O => \N__23436\,
            I => \N__23271\
        );

    \I__5508\ : Span4Mux_h
    port map (
            O => \N__23431\,
            I => \N__23271\
        );

    \I__5507\ : LocalMux
    port map (
            O => \N__23428\,
            I => \N__23271\
        );

    \I__5506\ : Span4Mux_v
    port map (
            O => \N__23425\,
            I => \N__23264\
        );

    \I__5505\ : Span4Mux_v
    port map (
            O => \N__23422\,
            I => \N__23264\
        );

    \I__5504\ : LocalMux
    port map (
            O => \N__23419\,
            I => \N__23264\
        );

    \I__5503\ : ClkMux
    port map (
            O => \N__23418\,
            I => \N__23261\
        );

    \I__5502\ : ClkMux
    port map (
            O => \N__23417\,
            I => \N__23258\
        );

    \I__5501\ : LocalMux
    port map (
            O => \N__23414\,
            I => \N__23254\
        );

    \I__5500\ : ClkMux
    port map (
            O => \N__23413\,
            I => \N__23250\
        );

    \I__5499\ : LocalMux
    port map (
            O => \N__23410\,
            I => \N__23245\
        );

    \I__5498\ : ClkMux
    port map (
            O => \N__23409\,
            I => \N__23242\
        );

    \I__5497\ : LocalMux
    port map (
            O => \N__23406\,
            I => \N__23239\
        );

    \I__5496\ : ClkMux
    port map (
            O => \N__23405\,
            I => \N__23236\
        );

    \I__5495\ : ClkMux
    port map (
            O => \N__23404\,
            I => \N__23233\
        );

    \I__5494\ : ClkMux
    port map (
            O => \N__23403\,
            I => \N__23229\
        );

    \I__5493\ : Span4Mux_h
    port map (
            O => \N__23400\,
            I => \N__23216\
        );

    \I__5492\ : Span4Mux_v
    port map (
            O => \N__23395\,
            I => \N__23216\
        );

    \I__5491\ : Span4Mux_h
    port map (
            O => \N__23390\,
            I => \N__23216\
        );

    \I__5490\ : LocalMux
    port map (
            O => \N__23387\,
            I => \N__23216\
        );

    \I__5489\ : LocalMux
    port map (
            O => \N__23384\,
            I => \N__23216\
        );

    \I__5488\ : ClkMux
    port map (
            O => \N__23383\,
            I => \N__23213\
        );

    \I__5487\ : Span4Mux_v
    port map (
            O => \N__23380\,
            I => \N__23208\
        );

    \I__5486\ : LocalMux
    port map (
            O => \N__23377\,
            I => \N__23208\
        );

    \I__5485\ : ClkMux
    port map (
            O => \N__23376\,
            I => \N__23205\
        );

    \I__5484\ : ClkMux
    port map (
            O => \N__23375\,
            I => \N__23202\
        );

    \I__5483\ : Span4Mux_v
    port map (
            O => \N__23368\,
            I => \N__23194\
        );

    \I__5482\ : Span4Mux_h
    port map (
            O => \N__23365\,
            I => \N__23194\
        );

    \I__5481\ : LocalMux
    port map (
            O => \N__23362\,
            I => \N__23194\
        );

    \I__5480\ : LocalMux
    port map (
            O => \N__23359\,
            I => \N__23191\
        );

    \I__5479\ : ClkMux
    port map (
            O => \N__23358\,
            I => \N__23188\
        );

    \I__5478\ : ClkMux
    port map (
            O => \N__23357\,
            I => \N__23185\
        );

    \I__5477\ : Span4Mux_h
    port map (
            O => \N__23350\,
            I => \N__23177\
        );

    \I__5476\ : Span4Mux_v
    port map (
            O => \N__23343\,
            I => \N__23177\
        );

    \I__5475\ : LocalMux
    port map (
            O => \N__23340\,
            I => \N__23177\
        );

    \I__5474\ : LocalMux
    port map (
            O => \N__23337\,
            I => \N__23174\
        );

    \I__5473\ : ClkMux
    port map (
            O => \N__23336\,
            I => \N__23171\
        );

    \I__5472\ : ClkMux
    port map (
            O => \N__23335\,
            I => \N__23168\
        );

    \I__5471\ : LocalMux
    port map (
            O => \N__23332\,
            I => \N__23165\
        );

    \I__5470\ : ClkMux
    port map (
            O => \N__23331\,
            I => \N__23162\
        );

    \I__5469\ : Span4Mux_v
    port map (
            O => \N__23328\,
            I => \N__23157\
        );

    \I__5468\ : LocalMux
    port map (
            O => \N__23325\,
            I => \N__23157\
        );

    \I__5467\ : ClkMux
    port map (
            O => \N__23324\,
            I => \N__23154\
        );

    \I__5466\ : Span4Mux_v
    port map (
            O => \N__23321\,
            I => \N__23149\
        );

    \I__5465\ : LocalMux
    port map (
            O => \N__23318\,
            I => \N__23149\
        );

    \I__5464\ : Span4Mux_h
    port map (
            O => \N__23315\,
            I => \N__23144\
        );

    \I__5463\ : LocalMux
    port map (
            O => \N__23312\,
            I => \N__23144\
        );

    \I__5462\ : Span4Mux_v
    port map (
            O => \N__23309\,
            I => \N__23137\
        );

    \I__5461\ : Span4Mux_h
    port map (
            O => \N__23306\,
            I => \N__23137\
        );

    \I__5460\ : LocalMux
    port map (
            O => \N__23303\,
            I => \N__23137\
        );

    \I__5459\ : ClkMux
    port map (
            O => \N__23302\,
            I => \N__23134\
        );

    \I__5458\ : LocalMux
    port map (
            O => \N__23299\,
            I => \N__23129\
        );

    \I__5457\ : ClkMux
    port map (
            O => \N__23298\,
            I => \N__23126\
        );

    \I__5456\ : Span4Mux_v
    port map (
            O => \N__23295\,
            I => \N__23118\
        );

    \I__5455\ : Span4Mux_h
    port map (
            O => \N__23288\,
            I => \N__23118\
        );

    \I__5454\ : Span4Mux_h
    port map (
            O => \N__23285\,
            I => \N__23118\
        );

    \I__5453\ : LocalMux
    port map (
            O => \N__23282\,
            I => \N__23115\
        );

    \I__5452\ : LocalMux
    port map (
            O => \N__23279\,
            I => \N__23112\
        );

    \I__5451\ : IoInMux
    port map (
            O => \N__23278\,
            I => \N__23109\
        );

    \I__5450\ : Span4Mux_h
    port map (
            O => \N__23271\,
            I => \N__23106\
        );

    \I__5449\ : Span4Mux_h
    port map (
            O => \N__23264\,
            I => \N__23099\
        );

    \I__5448\ : LocalMux
    port map (
            O => \N__23261\,
            I => \N__23099\
        );

    \I__5447\ : LocalMux
    port map (
            O => \N__23258\,
            I => \N__23099\
        );

    \I__5446\ : ClkMux
    port map (
            O => \N__23257\,
            I => \N__23096\
        );

    \I__5445\ : Span4Mux_h
    port map (
            O => \N__23254\,
            I => \N__23093\
        );

    \I__5444\ : ClkMux
    port map (
            O => \N__23253\,
            I => \N__23090\
        );

    \I__5443\ : LocalMux
    port map (
            O => \N__23250\,
            I => \N__23087\
        );

    \I__5442\ : ClkMux
    port map (
            O => \N__23249\,
            I => \N__23084\
        );

    \I__5441\ : ClkMux
    port map (
            O => \N__23248\,
            I => \N__23080\
        );

    \I__5440\ : Span4Mux_v
    port map (
            O => \N__23245\,
            I => \N__23075\
        );

    \I__5439\ : LocalMux
    port map (
            O => \N__23242\,
            I => \N__23075\
        );

    \I__5438\ : Span4Mux_v
    port map (
            O => \N__23239\,
            I => \N__23068\
        );

    \I__5437\ : LocalMux
    port map (
            O => \N__23236\,
            I => \N__23068\
        );

    \I__5436\ : LocalMux
    port map (
            O => \N__23233\,
            I => \N__23068\
        );

    \I__5435\ : ClkMux
    port map (
            O => \N__23232\,
            I => \N__23065\
        );

    \I__5434\ : LocalMux
    port map (
            O => \N__23229\,
            I => \N__23062\
        );

    \I__5433\ : ClkMux
    port map (
            O => \N__23228\,
            I => \N__23059\
        );

    \I__5432\ : ClkMux
    port map (
            O => \N__23227\,
            I => \N__23056\
        );

    \I__5431\ : Span4Mux_h
    port map (
            O => \N__23216\,
            I => \N__23051\
        );

    \I__5430\ : LocalMux
    port map (
            O => \N__23213\,
            I => \N__23051\
        );

    \I__5429\ : Span4Mux_h
    port map (
            O => \N__23208\,
            I => \N__23046\
        );

    \I__5428\ : LocalMux
    port map (
            O => \N__23205\,
            I => \N__23046\
        );

    \I__5427\ : LocalMux
    port map (
            O => \N__23202\,
            I => \N__23043\
        );

    \I__5426\ : ClkMux
    port map (
            O => \N__23201\,
            I => \N__23040\
        );

    \I__5425\ : Span4Mux_v
    port map (
            O => \N__23194\,
            I => \N__23030\
        );

    \I__5424\ : Span4Mux_h
    port map (
            O => \N__23191\,
            I => \N__23030\
        );

    \I__5423\ : LocalMux
    port map (
            O => \N__23188\,
            I => \N__23030\
        );

    \I__5422\ : LocalMux
    port map (
            O => \N__23185\,
            I => \N__23027\
        );

    \I__5421\ : ClkMux
    port map (
            O => \N__23184\,
            I => \N__23024\
        );

    \I__5420\ : Span4Mux_v
    port map (
            O => \N__23177\,
            I => \N__23020\
        );

    \I__5419\ : Span4Mux_v
    port map (
            O => \N__23174\,
            I => \N__23015\
        );

    \I__5418\ : LocalMux
    port map (
            O => \N__23171\,
            I => \N__23015\
        );

    \I__5417\ : LocalMux
    port map (
            O => \N__23168\,
            I => \N__23012\
        );

    \I__5416\ : Span4Mux_v
    port map (
            O => \N__23165\,
            I => \N__23003\
        );

    \I__5415\ : LocalMux
    port map (
            O => \N__23162\,
            I => \N__23003\
        );

    \I__5414\ : Span4Mux_v
    port map (
            O => \N__23157\,
            I => \N__23003\
        );

    \I__5413\ : LocalMux
    port map (
            O => \N__23154\,
            I => \N__23003\
        );

    \I__5412\ : Span4Mux_h
    port map (
            O => \N__23149\,
            I => \N__22994\
        );

    \I__5411\ : Span4Mux_v
    port map (
            O => \N__23144\,
            I => \N__22994\
        );

    \I__5410\ : Span4Mux_h
    port map (
            O => \N__23137\,
            I => \N__22994\
        );

    \I__5409\ : LocalMux
    port map (
            O => \N__23134\,
            I => \N__22994\
        );

    \I__5408\ : ClkMux
    port map (
            O => \N__23133\,
            I => \N__22991\
        );

    \I__5407\ : ClkMux
    port map (
            O => \N__23132\,
            I => \N__22988\
        );

    \I__5406\ : Span4Mux_v
    port map (
            O => \N__23129\,
            I => \N__22982\
        );

    \I__5405\ : LocalMux
    port map (
            O => \N__23126\,
            I => \N__22982\
        );

    \I__5404\ : ClkMux
    port map (
            O => \N__23125\,
            I => \N__22979\
        );

    \I__5403\ : Span4Mux_v
    port map (
            O => \N__23118\,
            I => \N__22972\
        );

    \I__5402\ : Span4Mux_h
    port map (
            O => \N__23115\,
            I => \N__22972\
        );

    \I__5401\ : Span4Mux_h
    port map (
            O => \N__23112\,
            I => \N__22972\
        );

    \I__5400\ : LocalMux
    port map (
            O => \N__23109\,
            I => \N__22969\
        );

    \I__5399\ : Span4Mux_v
    port map (
            O => \N__23106\,
            I => \N__22964\
        );

    \I__5398\ : Span4Mux_h
    port map (
            O => \N__23099\,
            I => \N__22964\
        );

    \I__5397\ : LocalMux
    port map (
            O => \N__23096\,
            I => \N__22961\
        );

    \I__5396\ : Span4Mux_v
    port map (
            O => \N__23093\,
            I => \N__22956\
        );

    \I__5395\ : LocalMux
    port map (
            O => \N__23090\,
            I => \N__22956\
        );

    \I__5394\ : Span4Mux_h
    port map (
            O => \N__23087\,
            I => \N__22952\
        );

    \I__5393\ : LocalMux
    port map (
            O => \N__23084\,
            I => \N__22949\
        );

    \I__5392\ : ClkMux
    port map (
            O => \N__23083\,
            I => \N__22946\
        );

    \I__5391\ : LocalMux
    port map (
            O => \N__23080\,
            I => \N__22943\
        );

    \I__5390\ : Span4Mux_v
    port map (
            O => \N__23075\,
            I => \N__22936\
        );

    \I__5389\ : Span4Mux_h
    port map (
            O => \N__23068\,
            I => \N__22936\
        );

    \I__5388\ : LocalMux
    port map (
            O => \N__23065\,
            I => \N__22936\
        );

    \I__5387\ : Span4Mux_h
    port map (
            O => \N__23062\,
            I => \N__22931\
        );

    \I__5386\ : LocalMux
    port map (
            O => \N__23059\,
            I => \N__22931\
        );

    \I__5385\ : LocalMux
    port map (
            O => \N__23056\,
            I => \N__22928\
        );

    \I__5384\ : Span4Mux_v
    port map (
            O => \N__23051\,
            I => \N__22919\
        );

    \I__5383\ : Span4Mux_h
    port map (
            O => \N__23046\,
            I => \N__22919\
        );

    \I__5382\ : Span4Mux_h
    port map (
            O => \N__23043\,
            I => \N__22919\
        );

    \I__5381\ : LocalMux
    port map (
            O => \N__23040\,
            I => \N__22919\
        );

    \I__5380\ : ClkMux
    port map (
            O => \N__23039\,
            I => \N__22916\
        );

    \I__5379\ : ClkMux
    port map (
            O => \N__23038\,
            I => \N__22913\
        );

    \I__5378\ : ClkMux
    port map (
            O => \N__23037\,
            I => \N__22909\
        );

    \I__5377\ : Span4Mux_v
    port map (
            O => \N__23030\,
            I => \N__22901\
        );

    \I__5376\ : Span4Mux_h
    port map (
            O => \N__23027\,
            I => \N__22901\
        );

    \I__5375\ : LocalMux
    port map (
            O => \N__23024\,
            I => \N__22901\
        );

    \I__5374\ : ClkMux
    port map (
            O => \N__23023\,
            I => \N__22898\
        );

    \I__5373\ : Span4Mux_v
    port map (
            O => \N__23020\,
            I => \N__22895\
        );

    \I__5372\ : Span4Mux_v
    port map (
            O => \N__23015\,
            I => \N__22892\
        );

    \I__5371\ : Span4Mux_v
    port map (
            O => \N__23012\,
            I => \N__22887\
        );

    \I__5370\ : Span4Mux_h
    port map (
            O => \N__23003\,
            I => \N__22887\
        );

    \I__5369\ : Span4Mux_h
    port map (
            O => \N__22994\,
            I => \N__22880\
        );

    \I__5368\ : LocalMux
    port map (
            O => \N__22991\,
            I => \N__22880\
        );

    \I__5367\ : LocalMux
    port map (
            O => \N__22988\,
            I => \N__22880\
        );

    \I__5366\ : ClkMux
    port map (
            O => \N__22987\,
            I => \N__22877\
        );

    \I__5365\ : Span4Mux_h
    port map (
            O => \N__22982\,
            I => \N__22873\
        );

    \I__5364\ : LocalMux
    port map (
            O => \N__22979\,
            I => \N__22870\
        );

    \I__5363\ : Span4Mux_v
    port map (
            O => \N__22972\,
            I => \N__22866\
        );

    \I__5362\ : IoSpan4Mux
    port map (
            O => \N__22969\,
            I => \N__22863\
        );

    \I__5361\ : Span4Mux_v
    port map (
            O => \N__22964\,
            I => \N__22858\
        );

    \I__5360\ : Span4Mux_h
    port map (
            O => \N__22961\,
            I => \N__22858\
        );

    \I__5359\ : Span4Mux_h
    port map (
            O => \N__22956\,
            I => \N__22855\
        );

    \I__5358\ : ClkMux
    port map (
            O => \N__22955\,
            I => \N__22852\
        );

    \I__5357\ : Span4Mux_v
    port map (
            O => \N__22952\,
            I => \N__22847\
        );

    \I__5356\ : Span4Mux_h
    port map (
            O => \N__22949\,
            I => \N__22847\
        );

    \I__5355\ : LocalMux
    port map (
            O => \N__22946\,
            I => \N__22844\
        );

    \I__5354\ : Span4Mux_h
    port map (
            O => \N__22943\,
            I => \N__22841\
        );

    \I__5353\ : Span4Mux_v
    port map (
            O => \N__22936\,
            I => \N__22830\
        );

    \I__5352\ : Span4Mux_h
    port map (
            O => \N__22931\,
            I => \N__22830\
        );

    \I__5351\ : Span4Mux_h
    port map (
            O => \N__22928\,
            I => \N__22830\
        );

    \I__5350\ : Span4Mux_v
    port map (
            O => \N__22919\,
            I => \N__22830\
        );

    \I__5349\ : LocalMux
    port map (
            O => \N__22916\,
            I => \N__22830\
        );

    \I__5348\ : LocalMux
    port map (
            O => \N__22913\,
            I => \N__22827\
        );

    \I__5347\ : ClkMux
    port map (
            O => \N__22912\,
            I => \N__22824\
        );

    \I__5346\ : LocalMux
    port map (
            O => \N__22909\,
            I => \N__22821\
        );

    \I__5345\ : ClkMux
    port map (
            O => \N__22908\,
            I => \N__22818\
        );

    \I__5344\ : Span4Mux_v
    port map (
            O => \N__22901\,
            I => \N__22815\
        );

    \I__5343\ : LocalMux
    port map (
            O => \N__22898\,
            I => \N__22812\
        );

    \I__5342\ : Span4Mux_h
    port map (
            O => \N__22895\,
            I => \N__22807\
        );

    \I__5341\ : Span4Mux_v
    port map (
            O => \N__22892\,
            I => \N__22807\
        );

    \I__5340\ : Span4Mux_h
    port map (
            O => \N__22887\,
            I => \N__22800\
        );

    \I__5339\ : Span4Mux_v
    port map (
            O => \N__22880\,
            I => \N__22800\
        );

    \I__5338\ : LocalMux
    port map (
            O => \N__22877\,
            I => \N__22800\
        );

    \I__5337\ : ClkMux
    port map (
            O => \N__22876\,
            I => \N__22797\
        );

    \I__5336\ : Span4Mux_h
    port map (
            O => \N__22873\,
            I => \N__22792\
        );

    \I__5335\ : Span4Mux_v
    port map (
            O => \N__22870\,
            I => \N__22792\
        );

    \I__5334\ : ClkMux
    port map (
            O => \N__22869\,
            I => \N__22789\
        );

    \I__5333\ : Span4Mux_v
    port map (
            O => \N__22866\,
            I => \N__22786\
        );

    \I__5332\ : IoSpan4Mux
    port map (
            O => \N__22863\,
            I => \N__22783\
        );

    \I__5331\ : Span4Mux_v
    port map (
            O => \N__22858\,
            I => \N__22780\
        );

    \I__5330\ : Span4Mux_h
    port map (
            O => \N__22855\,
            I => \N__22777\
        );

    \I__5329\ : LocalMux
    port map (
            O => \N__22852\,
            I => \N__22774\
        );

    \I__5328\ : Span4Mux_h
    port map (
            O => \N__22847\,
            I => \N__22771\
        );

    \I__5327\ : Span4Mux_h
    port map (
            O => \N__22844\,
            I => \N__22768\
        );

    \I__5326\ : Span4Mux_v
    port map (
            O => \N__22841\,
            I => \N__22761\
        );

    \I__5325\ : Span4Mux_v
    port map (
            O => \N__22830\,
            I => \N__22761\
        );

    \I__5324\ : Span4Mux_h
    port map (
            O => \N__22827\,
            I => \N__22761\
        );

    \I__5323\ : LocalMux
    port map (
            O => \N__22824\,
            I => \N__22758\
        );

    \I__5322\ : Span12Mux_h
    port map (
            O => \N__22821\,
            I => \N__22753\
        );

    \I__5321\ : LocalMux
    port map (
            O => \N__22818\,
            I => \N__22753\
        );

    \I__5320\ : Sp12to4
    port map (
            O => \N__22815\,
            I => \N__22746\
        );

    \I__5319\ : Sp12to4
    port map (
            O => \N__22812\,
            I => \N__22746\
        );

    \I__5318\ : Sp12to4
    port map (
            O => \N__22807\,
            I => \N__22746\
        );

    \I__5317\ : Span4Mux_v
    port map (
            O => \N__22800\,
            I => \N__22737\
        );

    \I__5316\ : LocalMux
    port map (
            O => \N__22797\,
            I => \N__22737\
        );

    \I__5315\ : Span4Mux_v
    port map (
            O => \N__22792\,
            I => \N__22737\
        );

    \I__5314\ : LocalMux
    port map (
            O => \N__22789\,
            I => \N__22737\
        );

    \I__5313\ : IoSpan4Mux
    port map (
            O => \N__22786\,
            I => \N__22732\
        );

    \I__5312\ : IoSpan4Mux
    port map (
            O => \N__22783\,
            I => \N__22732\
        );

    \I__5311\ : Span4Mux_v
    port map (
            O => \N__22780\,
            I => \N__22729\
        );

    \I__5310\ : Span4Mux_h
    port map (
            O => \N__22777\,
            I => \N__22726\
        );

    \I__5309\ : Span12Mux_h
    port map (
            O => \N__22774\,
            I => \N__22723\
        );

    \I__5308\ : Span4Mux_h
    port map (
            O => \N__22771\,
            I => \N__22716\
        );

    \I__5307\ : Span4Mux_h
    port map (
            O => \N__22768\,
            I => \N__22716\
        );

    \I__5306\ : Span4Mux_v
    port map (
            O => \N__22761\,
            I => \N__22716\
        );

    \I__5305\ : Span12Mux_h
    port map (
            O => \N__22758\,
            I => \N__22707\
        );

    \I__5304\ : Span12Mux_v
    port map (
            O => \N__22753\,
            I => \N__22707\
        );

    \I__5303\ : Span12Mux_h
    port map (
            O => \N__22746\,
            I => \N__22707\
        );

    \I__5302\ : Sp12to4
    port map (
            O => \N__22737\,
            I => \N__22707\
        );

    \I__5301\ : Odrv4
    port map (
            O => \N__22732\,
            I => \ADV_CLK_c\
        );

    \I__5300\ : Odrv4
    port map (
            O => \N__22729\,
            I => \ADV_CLK_c\
        );

    \I__5299\ : Odrv4
    port map (
            O => \N__22726\,
            I => \ADV_CLK_c\
        );

    \I__5298\ : Odrv12
    port map (
            O => \N__22723\,
            I => \ADV_CLK_c\
        );

    \I__5297\ : Odrv4
    port map (
            O => \N__22716\,
            I => \ADV_CLK_c\
        );

    \I__5296\ : Odrv12
    port map (
            O => \N__22707\,
            I => \ADV_CLK_c\
        );

    \I__5295\ : SRMux
    port map (
            O => \N__22694\,
            I => \N__22689\
        );

    \I__5294\ : SRMux
    port map (
            O => \N__22693\,
            I => \N__22684\
        );

    \I__5293\ : SRMux
    port map (
            O => \N__22692\,
            I => \N__22681\
        );

    \I__5292\ : LocalMux
    port map (
            O => \N__22689\,
            I => \N__22677\
        );

    \I__5291\ : SRMux
    port map (
            O => \N__22688\,
            I => \N__22674\
        );

    \I__5290\ : SRMux
    port map (
            O => \N__22687\,
            I => \N__22671\
        );

    \I__5289\ : LocalMux
    port map (
            O => \N__22684\,
            I => \N__22667\
        );

    \I__5288\ : LocalMux
    port map (
            O => \N__22681\,
            I => \N__22664\
        );

    \I__5287\ : SRMux
    port map (
            O => \N__22680\,
            I => \N__22661\
        );

    \I__5286\ : Span4Mux_h
    port map (
            O => \N__22677\,
            I => \N__22656\
        );

    \I__5285\ : LocalMux
    port map (
            O => \N__22674\,
            I => \N__22656\
        );

    \I__5284\ : LocalMux
    port map (
            O => \N__22671\,
            I => \N__22653\
        );

    \I__5283\ : SRMux
    port map (
            O => \N__22670\,
            I => \N__22650\
        );

    \I__5282\ : Span4Mux_v
    port map (
            O => \N__22667\,
            I => \N__22646\
        );

    \I__5281\ : Span4Mux_v
    port map (
            O => \N__22664\,
            I => \N__22641\
        );

    \I__5280\ : LocalMux
    port map (
            O => \N__22661\,
            I => \N__22641\
        );

    \I__5279\ : Span4Mux_h
    port map (
            O => \N__22656\,
            I => \N__22634\
        );

    \I__5278\ : Span4Mux_h
    port map (
            O => \N__22653\,
            I => \N__22634\
        );

    \I__5277\ : LocalMux
    port map (
            O => \N__22650\,
            I => \N__22634\
        );

    \I__5276\ : SRMux
    port map (
            O => \N__22649\,
            I => \N__22631\
        );

    \I__5275\ : Span4Mux_h
    port map (
            O => \N__22646\,
            I => \N__22626\
        );

    \I__5274\ : Span4Mux_v
    port map (
            O => \N__22641\,
            I => \N__22626\
        );

    \I__5273\ : Span4Mux_v
    port map (
            O => \N__22634\,
            I => \N__22623\
        );

    \I__5272\ : LocalMux
    port map (
            O => \N__22631\,
            I => \N__22620\
        );

    \I__5271\ : Odrv4
    port map (
            O => \N__22626\,
            I => \transmit_module.n2388\
        );

    \I__5270\ : Odrv4
    port map (
            O => \N__22623\,
            I => \transmit_module.n2388\
        );

    \I__5269\ : Odrv12
    port map (
            O => \N__22620\,
            I => \transmit_module.n2388\
        );

    \I__5268\ : InMux
    port map (
            O => \N__22613\,
            I => \N__22610\
        );

    \I__5267\ : LocalMux
    port map (
            O => \N__22610\,
            I => \N__22607\
        );

    \I__5266\ : Span4Mux_v
    port map (
            O => \N__22607\,
            I => \N__22604\
        );

    \I__5265\ : Sp12to4
    port map (
            O => \N__22604\,
            I => \N__22601\
        );

    \I__5264\ : Odrv12
    port map (
            O => \N__22601\,
            I => \line_buffer.n596\
        );

    \I__5263\ : InMux
    port map (
            O => \N__22598\,
            I => \N__22595\
        );

    \I__5262\ : LocalMux
    port map (
            O => \N__22595\,
            I => \N__22592\
        );

    \I__5261\ : Span4Mux_h
    port map (
            O => \N__22592\,
            I => \N__22589\
        );

    \I__5260\ : Span4Mux_v
    port map (
            O => \N__22589\,
            I => \N__22586\
        );

    \I__5259\ : Span4Mux_v
    port map (
            O => \N__22586\,
            I => \N__22583\
        );

    \I__5258\ : Span4Mux_h
    port map (
            O => \N__22583\,
            I => \N__22580\
        );

    \I__5257\ : Odrv4
    port map (
            O => \N__22580\,
            I => \line_buffer.n588\
        );

    \I__5256\ : InMux
    port map (
            O => \N__22577\,
            I => \N__22574\
        );

    \I__5255\ : LocalMux
    port map (
            O => \N__22574\,
            I => \line_buffer.n3644\
        );

    \I__5254\ : InMux
    port map (
            O => \N__22571\,
            I => \N__22568\
        );

    \I__5253\ : LocalMux
    port map (
            O => \N__22568\,
            I => \N__22565\
        );

    \I__5252\ : Span4Mux_h
    port map (
            O => \N__22565\,
            I => \N__22562\
        );

    \I__5251\ : Span4Mux_h
    port map (
            O => \N__22562\,
            I => \N__22559\
        );

    \I__5250\ : Odrv4
    port map (
            O => \N__22559\,
            I => \line_buffer.n473\
        );

    \I__5249\ : InMux
    port map (
            O => \N__22556\,
            I => \N__22553\
        );

    \I__5248\ : LocalMux
    port map (
            O => \N__22553\,
            I => \N__22550\
        );

    \I__5247\ : Span4Mux_v
    port map (
            O => \N__22550\,
            I => \N__22547\
        );

    \I__5246\ : Sp12to4
    port map (
            O => \N__22547\,
            I => \N__22544\
        );

    \I__5245\ : Odrv12
    port map (
            O => \N__22544\,
            I => \line_buffer.n465\
        );

    \I__5244\ : InMux
    port map (
            O => \N__22541\,
            I => \N__22538\
        );

    \I__5243\ : LocalMux
    port map (
            O => \N__22538\,
            I => \N__22535\
        );

    \I__5242\ : Odrv12
    port map (
            O => \N__22535\,
            I => \line_buffer.n3575\
        );

    \I__5241\ : InMux
    port map (
            O => \N__22532\,
            I => \N__22529\
        );

    \I__5240\ : LocalMux
    port map (
            O => \N__22529\,
            I => \N__22526\
        );

    \I__5239\ : Odrv12
    port map (
            O => \N__22526\,
            I => \tvp_video_buffer.BUFFER_1_9\
        );

    \I__5238\ : InMux
    port map (
            O => \N__22523\,
            I => \N__22520\
        );

    \I__5237\ : LocalMux
    port map (
            O => \N__22520\,
            I => \N__22514\
        );

    \I__5236\ : InMux
    port map (
            O => \N__22519\,
            I => \N__22510\
        );

    \I__5235\ : InMux
    port map (
            O => \N__22518\,
            I => \N__22507\
        );

    \I__5234\ : InMux
    port map (
            O => \N__22517\,
            I => \N__22503\
        );

    \I__5233\ : Span4Mux_s2_v
    port map (
            O => \N__22514\,
            I => \N__22500\
        );

    \I__5232\ : InMux
    port map (
            O => \N__22513\,
            I => \N__22497\
        );

    \I__5231\ : LocalMux
    port map (
            O => \N__22510\,
            I => \N__22493\
        );

    \I__5230\ : LocalMux
    port map (
            O => \N__22507\,
            I => \N__22490\
        );

    \I__5229\ : InMux
    port map (
            O => \N__22506\,
            I => \N__22487\
        );

    \I__5228\ : LocalMux
    port map (
            O => \N__22503\,
            I => \N__22484\
        );

    \I__5227\ : Span4Mux_v
    port map (
            O => \N__22500\,
            I => \N__22478\
        );

    \I__5226\ : LocalMux
    port map (
            O => \N__22497\,
            I => \N__22478\
        );

    \I__5225\ : InMux
    port map (
            O => \N__22496\,
            I => \N__22475\
        );

    \I__5224\ : Span4Mux_h
    port map (
            O => \N__22493\,
            I => \N__22472\
        );

    \I__5223\ : Span4Mux_v
    port map (
            O => \N__22490\,
            I => \N__22469\
        );

    \I__5222\ : LocalMux
    port map (
            O => \N__22487\,
            I => \N__22466\
        );

    \I__5221\ : Span4Mux_v
    port map (
            O => \N__22484\,
            I => \N__22463\
        );

    \I__5220\ : InMux
    port map (
            O => \N__22483\,
            I => \N__22460\
        );

    \I__5219\ : Span4Mux_h
    port map (
            O => \N__22478\,
            I => \N__22457\
        );

    \I__5218\ : LocalMux
    port map (
            O => \N__22475\,
            I => \N__22453\
        );

    \I__5217\ : Span4Mux_v
    port map (
            O => \N__22472\,
            I => \N__22450\
        );

    \I__5216\ : Span4Mux_v
    port map (
            O => \N__22469\,
            I => \N__22445\
        );

    \I__5215\ : Span4Mux_h
    port map (
            O => \N__22466\,
            I => \N__22445\
        );

    \I__5214\ : Span4Mux_v
    port map (
            O => \N__22463\,
            I => \N__22440\
        );

    \I__5213\ : LocalMux
    port map (
            O => \N__22460\,
            I => \N__22440\
        );

    \I__5212\ : Span4Mux_h
    port map (
            O => \N__22457\,
            I => \N__22437\
        );

    \I__5211\ : InMux
    port map (
            O => \N__22456\,
            I => \N__22434\
        );

    \I__5210\ : Span12Mux_h
    port map (
            O => \N__22453\,
            I => \N__22431\
        );

    \I__5209\ : Sp12to4
    port map (
            O => \N__22450\,
            I => \N__22428\
        );

    \I__5208\ : Span4Mux_v
    port map (
            O => \N__22445\,
            I => \N__22423\
        );

    \I__5207\ : Span4Mux_v
    port map (
            O => \N__22440\,
            I => \N__22423\
        );

    \I__5206\ : Sp12to4
    port map (
            O => \N__22437\,
            I => \N__22418\
        );

    \I__5205\ : LocalMux
    port map (
            O => \N__22434\,
            I => \N__22418\
        );

    \I__5204\ : Span12Mux_v
    port map (
            O => \N__22431\,
            I => \N__22409\
        );

    \I__5203\ : Span12Mux_h
    port map (
            O => \N__22428\,
            I => \N__22409\
        );

    \I__5202\ : Sp12to4
    port map (
            O => \N__22423\,
            I => \N__22409\
        );

    \I__5201\ : Span12Mux_v
    port map (
            O => \N__22418\,
            I => \N__22409\
        );

    \I__5200\ : Odrv12
    port map (
            O => \N__22409\,
            I => \RX_DATA_5\
        );

    \I__5199\ : InMux
    port map (
            O => \N__22406\,
            I => \N__22403\
        );

    \I__5198\ : LocalMux
    port map (
            O => \N__22403\,
            I => \N__22400\
        );

    \I__5197\ : Span12Mux_v
    port map (
            O => \N__22400\,
            I => \N__22397\
        );

    \I__5196\ : Odrv12
    port map (
            O => \N__22397\,
            I => \line_buffer.n601\
        );

    \I__5195\ : CascadeMux
    port map (
            O => \N__22394\,
            I => \N__22385\
        );

    \I__5194\ : CascadeMux
    port map (
            O => \N__22393\,
            I => \N__22382\
        );

    \I__5193\ : CascadeMux
    port map (
            O => \N__22392\,
            I => \N__22378\
        );

    \I__5192\ : InMux
    port map (
            O => \N__22391\,
            I => \N__22369\
        );

    \I__5191\ : InMux
    port map (
            O => \N__22390\,
            I => \N__22366\
        );

    \I__5190\ : InMux
    port map (
            O => \N__22389\,
            I => \N__22363\
        );

    \I__5189\ : InMux
    port map (
            O => \N__22388\,
            I => \N__22360\
        );

    \I__5188\ : InMux
    port map (
            O => \N__22385\,
            I => \N__22357\
        );

    \I__5187\ : InMux
    port map (
            O => \N__22382\,
            I => \N__22354\
        );

    \I__5186\ : CascadeMux
    port map (
            O => \N__22381\,
            I => \N__22351\
        );

    \I__5185\ : InMux
    port map (
            O => \N__22378\,
            I => \N__22347\
        );

    \I__5184\ : CascadeMux
    port map (
            O => \N__22377\,
            I => \N__22343\
        );

    \I__5183\ : CascadeMux
    port map (
            O => \N__22376\,
            I => \N__22340\
        );

    \I__5182\ : InMux
    port map (
            O => \N__22375\,
            I => \N__22334\
        );

    \I__5181\ : InMux
    port map (
            O => \N__22374\,
            I => \N__22331\
        );

    \I__5180\ : CascadeMux
    port map (
            O => \N__22373\,
            I => \N__22328\
        );

    \I__5179\ : CascadeMux
    port map (
            O => \N__22372\,
            I => \N__22325\
        );

    \I__5178\ : LocalMux
    port map (
            O => \N__22369\,
            I => \N__22322\
        );

    \I__5177\ : LocalMux
    port map (
            O => \N__22366\,
            I => \N__22313\
        );

    \I__5176\ : LocalMux
    port map (
            O => \N__22363\,
            I => \N__22313\
        );

    \I__5175\ : LocalMux
    port map (
            O => \N__22360\,
            I => \N__22313\
        );

    \I__5174\ : LocalMux
    port map (
            O => \N__22357\,
            I => \N__22313\
        );

    \I__5173\ : LocalMux
    port map (
            O => \N__22354\,
            I => \N__22310\
        );

    \I__5172\ : InMux
    port map (
            O => \N__22351\,
            I => \N__22307\
        );

    \I__5171\ : InMux
    port map (
            O => \N__22350\,
            I => \N__22302\
        );

    \I__5170\ : LocalMux
    port map (
            O => \N__22347\,
            I => \N__22299\
        );

    \I__5169\ : InMux
    port map (
            O => \N__22346\,
            I => \N__22296\
        );

    \I__5168\ : InMux
    port map (
            O => \N__22343\,
            I => \N__22293\
        );

    \I__5167\ : InMux
    port map (
            O => \N__22340\,
            I => \N__22290\
        );

    \I__5166\ : InMux
    port map (
            O => \N__22339\,
            I => \N__22287\
        );

    \I__5165\ : InMux
    port map (
            O => \N__22338\,
            I => \N__22284\
        );

    \I__5164\ : InMux
    port map (
            O => \N__22337\,
            I => \N__22281\
        );

    \I__5163\ : LocalMux
    port map (
            O => \N__22334\,
            I => \N__22276\
        );

    \I__5162\ : LocalMux
    port map (
            O => \N__22331\,
            I => \N__22276\
        );

    \I__5161\ : InMux
    port map (
            O => \N__22328\,
            I => \N__22273\
        );

    \I__5160\ : InMux
    port map (
            O => \N__22325\,
            I => \N__22270\
        );

    \I__5159\ : Span4Mux_v
    port map (
            O => \N__22322\,
            I => \N__22260\
        );

    \I__5158\ : Span4Mux_v
    port map (
            O => \N__22313\,
            I => \N__22260\
        );

    \I__5157\ : Span4Mux_h
    port map (
            O => \N__22310\,
            I => \N__22260\
        );

    \I__5156\ : LocalMux
    port map (
            O => \N__22307\,
            I => \N__22260\
        );

    \I__5155\ : InMux
    port map (
            O => \N__22306\,
            I => \N__22257\
        );

    \I__5154\ : InMux
    port map (
            O => \N__22305\,
            I => \N__22254\
        );

    \I__5153\ : LocalMux
    port map (
            O => \N__22302\,
            I => \N__22249\
        );

    \I__5152\ : Span4Mux_v
    port map (
            O => \N__22299\,
            I => \N__22249\
        );

    \I__5151\ : LocalMux
    port map (
            O => \N__22296\,
            I => \N__22242\
        );

    \I__5150\ : LocalMux
    port map (
            O => \N__22293\,
            I => \N__22242\
        );

    \I__5149\ : LocalMux
    port map (
            O => \N__22290\,
            I => \N__22242\
        );

    \I__5148\ : LocalMux
    port map (
            O => \N__22287\,
            I => \N__22229\
        );

    \I__5147\ : LocalMux
    port map (
            O => \N__22284\,
            I => \N__22229\
        );

    \I__5146\ : LocalMux
    port map (
            O => \N__22281\,
            I => \N__22229\
        );

    \I__5145\ : Span4Mux_v
    port map (
            O => \N__22276\,
            I => \N__22229\
        );

    \I__5144\ : LocalMux
    port map (
            O => \N__22273\,
            I => \N__22229\
        );

    \I__5143\ : LocalMux
    port map (
            O => \N__22270\,
            I => \N__22229\
        );

    \I__5142\ : InMux
    port map (
            O => \N__22269\,
            I => \N__22226\
        );

    \I__5141\ : Span4Mux_h
    port map (
            O => \N__22260\,
            I => \N__22223\
        );

    \I__5140\ : LocalMux
    port map (
            O => \N__22257\,
            I => \N__22220\
        );

    \I__5139\ : LocalMux
    port map (
            O => \N__22254\,
            I => \N__22211\
        );

    \I__5138\ : Span4Mux_h
    port map (
            O => \N__22249\,
            I => \N__22211\
        );

    \I__5137\ : Span4Mux_v
    port map (
            O => \N__22242\,
            I => \N__22211\
        );

    \I__5136\ : Span4Mux_v
    port map (
            O => \N__22229\,
            I => \N__22211\
        );

    \I__5135\ : LocalMux
    port map (
            O => \N__22226\,
            I => \N__22208\
        );

    \I__5134\ : Span4Mux_h
    port map (
            O => \N__22223\,
            I => \N__22205\
        );

    \I__5133\ : Span4Mux_v
    port map (
            O => \N__22220\,
            I => \N__22200\
        );

    \I__5132\ : Span4Mux_h
    port map (
            O => \N__22211\,
            I => \N__22200\
        );

    \I__5131\ : Odrv4
    port map (
            O => \N__22208\,
            I => \TX_ADDR_12\
        );

    \I__5130\ : Odrv4
    port map (
            O => \N__22205\,
            I => \TX_ADDR_12\
        );

    \I__5129\ : Odrv4
    port map (
            O => \N__22200\,
            I => \TX_ADDR_12\
        );

    \I__5128\ : InMux
    port map (
            O => \N__22193\,
            I => \N__22190\
        );

    \I__5127\ : LocalMux
    port map (
            O => \N__22190\,
            I => \N__22187\
        );

    \I__5126\ : Span4Mux_v
    port map (
            O => \N__22187\,
            I => \N__22184\
        );

    \I__5125\ : Span4Mux_v
    port map (
            O => \N__22184\,
            I => \N__22181\
        );

    \I__5124\ : Span4Mux_h
    port map (
            O => \N__22181\,
            I => \N__22178\
        );

    \I__5123\ : Odrv4
    port map (
            O => \N__22178\,
            I => \line_buffer.n593\
        );

    \I__5122\ : InMux
    port map (
            O => \N__22175\,
            I => \N__22172\
        );

    \I__5121\ : LocalMux
    port map (
            O => \N__22172\,
            I => \line_buffer.n3596\
        );

    \I__5120\ : IoInMux
    port map (
            O => \N__22169\,
            I => \N__22166\
        );

    \I__5119\ : LocalMux
    port map (
            O => \N__22166\,
            I => \N__22162\
        );

    \I__5118\ : InMux
    port map (
            O => \N__22165\,
            I => \N__22159\
        );

    \I__5117\ : IoSpan4Mux
    port map (
            O => \N__22162\,
            I => \N__22156\
        );

    \I__5116\ : LocalMux
    port map (
            O => \N__22159\,
            I => \N__22153\
        );

    \I__5115\ : Span4Mux_s2_h
    port map (
            O => \N__22156\,
            I => \N__22150\
        );

    \I__5114\ : Span4Mux_v
    port map (
            O => \N__22153\,
            I => \N__22147\
        );

    \I__5113\ : Sp12to4
    port map (
            O => \N__22150\,
            I => \N__22144\
        );

    \I__5112\ : Sp12to4
    port map (
            O => \N__22147\,
            I => \N__22141\
        );

    \I__5111\ : Span12Mux_v
    port map (
            O => \N__22144\,
            I => \N__22138\
        );

    \I__5110\ : Span12Mux_h
    port map (
            O => \N__22141\,
            I => \N__22135\
        );

    \I__5109\ : Span12Mux_h
    port map (
            O => \N__22138\,
            I => \N__22132\
        );

    \I__5108\ : Span12Mux_v
    port map (
            O => \N__22135\,
            I => \N__22129\
        );

    \I__5107\ : Odrv12
    port map (
            O => \N__22132\,
            I => \DEBUG_c_7_c\
        );

    \I__5106\ : Odrv12
    port map (
            O => \N__22129\,
            I => \DEBUG_c_7_c\
        );

    \I__5105\ : InMux
    port map (
            O => \N__22124\,
            I => \N__22121\
        );

    \I__5104\ : LocalMux
    port map (
            O => \N__22121\,
            I => \N__22118\
        );

    \I__5103\ : Span4Mux_v
    port map (
            O => \N__22118\,
            I => \N__22115\
        );

    \I__5102\ : Span4Mux_h
    port map (
            O => \N__22115\,
            I => \N__22112\
        );

    \I__5101\ : Odrv4
    port map (
            O => \N__22112\,
            I => \line_buffer.n467\
        );

    \I__5100\ : CascadeMux
    port map (
            O => \N__22109\,
            I => \N__22106\
        );

    \I__5099\ : InMux
    port map (
            O => \N__22106\,
            I => \N__22103\
        );

    \I__5098\ : LocalMux
    port map (
            O => \N__22103\,
            I => \N__22100\
        );

    \I__5097\ : Span4Mux_v
    port map (
            O => \N__22100\,
            I => \N__22097\
        );

    \I__5096\ : Sp12to4
    port map (
            O => \N__22097\,
            I => \N__22094\
        );

    \I__5095\ : Span12Mux_h
    port map (
            O => \N__22094\,
            I => \N__22091\
        );

    \I__5094\ : Span12Mux_v
    port map (
            O => \N__22091\,
            I => \N__22088\
        );

    \I__5093\ : Odrv12
    port map (
            O => \N__22088\,
            I => \line_buffer.n459\
        );

    \I__5092\ : InMux
    port map (
            O => \N__22085\,
            I => \N__22082\
        );

    \I__5091\ : LocalMux
    port map (
            O => \N__22082\,
            I => \N__22079\
        );

    \I__5090\ : Odrv4
    port map (
            O => \N__22079\,
            I => \line_buffer.n3638\
        );

    \I__5089\ : InMux
    port map (
            O => \N__22076\,
            I => \N__22073\
        );

    \I__5088\ : LocalMux
    port map (
            O => \N__22073\,
            I => \line_buffer.n3641\
        );

    \I__5087\ : InMux
    port map (
            O => \N__22070\,
            I => \N__22067\
        );

    \I__5086\ : LocalMux
    port map (
            O => \N__22067\,
            I => \N__22064\
        );

    \I__5085\ : Span4Mux_v
    port map (
            O => \N__22064\,
            I => \N__22061\
        );

    \I__5084\ : Odrv4
    port map (
            O => \N__22061\,
            I => \TX_DATA_0\
        );

    \I__5083\ : InMux
    port map (
            O => \N__22058\,
            I => \N__22055\
        );

    \I__5082\ : LocalMux
    port map (
            O => \N__22055\,
            I => \N__22052\
        );

    \I__5081\ : Span4Mux_v
    port map (
            O => \N__22052\,
            I => \N__22049\
        );

    \I__5080\ : Span4Mux_v
    port map (
            O => \N__22049\,
            I => \N__22046\
        );

    \I__5079\ : Sp12to4
    port map (
            O => \N__22046\,
            I => \N__22043\
        );

    \I__5078\ : Span12Mux_h
    port map (
            O => \N__22043\,
            I => \N__22040\
        );

    \I__5077\ : Span12Mux_v
    port map (
            O => \N__22040\,
            I => \N__22037\
        );

    \I__5076\ : Odrv12
    port map (
            O => \N__22037\,
            I => \line_buffer.n532\
        );

    \I__5075\ : CascadeMux
    port map (
            O => \N__22034\,
            I => \N__22031\
        );

    \I__5074\ : InMux
    port map (
            O => \N__22031\,
            I => \N__22028\
        );

    \I__5073\ : LocalMux
    port map (
            O => \N__22028\,
            I => \N__22025\
        );

    \I__5072\ : Span4Mux_h
    port map (
            O => \N__22025\,
            I => \N__22022\
        );

    \I__5071\ : Span4Mux_h
    port map (
            O => \N__22022\,
            I => \N__22019\
        );

    \I__5070\ : Span4Mux_v
    port map (
            O => \N__22019\,
            I => \N__22016\
        );

    \I__5069\ : Span4Mux_v
    port map (
            O => \N__22016\,
            I => \N__22013\
        );

    \I__5068\ : Odrv4
    port map (
            O => \N__22013\,
            I => \line_buffer.n524\
        );

    \I__5067\ : InMux
    port map (
            O => \N__22010\,
            I => \N__22007\
        );

    \I__5066\ : LocalMux
    port map (
            O => \N__22007\,
            I => \line_buffer.n3647\
        );

    \I__5065\ : InMux
    port map (
            O => \N__22004\,
            I => \N__22001\
        );

    \I__5064\ : LocalMux
    port map (
            O => \N__22001\,
            I => \N__21998\
        );

    \I__5063\ : Odrv12
    port map (
            O => \N__21998\,
            I => \TX_DATA_5\
        );

    \I__5062\ : IoInMux
    port map (
            O => \N__21995\,
            I => \N__21991\
        );

    \I__5061\ : IoInMux
    port map (
            O => \N__21994\,
            I => \N__21988\
        );

    \I__5060\ : LocalMux
    port map (
            O => \N__21991\,
            I => \N__21985\
        );

    \I__5059\ : LocalMux
    port map (
            O => \N__21988\,
            I => \N__21981\
        );

    \I__5058\ : Span4Mux_s0_v
    port map (
            O => \N__21985\,
            I => \N__21978\
        );

    \I__5057\ : IoInMux
    port map (
            O => \N__21984\,
            I => \N__21975\
        );

    \I__5056\ : Span4Mux_s3_v
    port map (
            O => \N__21981\,
            I => \N__21972\
        );

    \I__5055\ : Sp12to4
    port map (
            O => \N__21978\,
            I => \N__21969\
        );

    \I__5054\ : LocalMux
    port map (
            O => \N__21975\,
            I => \N__21966\
        );

    \I__5053\ : Span4Mux_v
    port map (
            O => \N__21972\,
            I => \N__21963\
        );

    \I__5052\ : Span12Mux_h
    port map (
            O => \N__21969\,
            I => \N__21960\
        );

    \I__5051\ : Span12Mux_s6_h
    port map (
            O => \N__21966\,
            I => \N__21955\
        );

    \I__5050\ : Sp12to4
    port map (
            O => \N__21963\,
            I => \N__21955\
        );

    \I__5049\ : Odrv12
    port map (
            O => \N__21960\,
            I => n1816
        );

    \I__5048\ : Odrv12
    port map (
            O => \N__21955\,
            I => n1816
        );

    \I__5047\ : InMux
    port map (
            O => \N__21950\,
            I => \N__21947\
        );

    \I__5046\ : LocalMux
    port map (
            O => \N__21947\,
            I => \N__21944\
        );

    \I__5045\ : Span4Mux_v
    port map (
            O => \N__21944\,
            I => \N__21941\
        );

    \I__5044\ : Sp12to4
    port map (
            O => \N__21941\,
            I => \N__21938\
        );

    \I__5043\ : Span12Mux_v
    port map (
            O => \N__21938\,
            I => \N__21935\
        );

    \I__5042\ : Odrv12
    port map (
            O => \N__21935\,
            I => \line_buffer.n537\
        );

    \I__5041\ : CascadeMux
    port map (
            O => \N__21932\,
            I => \N__21929\
        );

    \I__5040\ : InMux
    port map (
            O => \N__21929\,
            I => \N__21926\
        );

    \I__5039\ : LocalMux
    port map (
            O => \N__21926\,
            I => \N__21923\
        );

    \I__5038\ : Span4Mux_h
    port map (
            O => \N__21923\,
            I => \N__21920\
        );

    \I__5037\ : Span4Mux_h
    port map (
            O => \N__21920\,
            I => \N__21917\
        );

    \I__5036\ : Span4Mux_v
    port map (
            O => \N__21917\,
            I => \N__21914\
        );

    \I__5035\ : Span4Mux_v
    port map (
            O => \N__21914\,
            I => \N__21911\
        );

    \I__5034\ : Odrv4
    port map (
            O => \N__21911\,
            I => \line_buffer.n529\
        );

    \I__5033\ : InMux
    port map (
            O => \N__21908\,
            I => \N__21905\
        );

    \I__5032\ : LocalMux
    port map (
            O => \N__21905\,
            I => \line_buffer.n3599\
        );

    \I__5031\ : InMux
    port map (
            O => \N__21902\,
            I => \N__21899\
        );

    \I__5030\ : LocalMux
    port map (
            O => \N__21899\,
            I => \N__21896\
        );

    \I__5029\ : Odrv12
    port map (
            O => \N__21896\,
            I => \line_buffer.n597\
        );

    \I__5028\ : InMux
    port map (
            O => \N__21893\,
            I => \N__21890\
        );

    \I__5027\ : LocalMux
    port map (
            O => \N__21890\,
            I => \N__21887\
        );

    \I__5026\ : Span12Mux_h
    port map (
            O => \N__21887\,
            I => \N__21884\
        );

    \I__5025\ : Span12Mux_v
    port map (
            O => \N__21884\,
            I => \N__21881\
        );

    \I__5024\ : Odrv12
    port map (
            O => \N__21881\,
            I => \line_buffer.n589\
        );

    \I__5023\ : InMux
    port map (
            O => \N__21878\,
            I => \N__21875\
        );

    \I__5022\ : LocalMux
    port map (
            O => \N__21875\,
            I => \N__21872\
        );

    \I__5021\ : Span4Mux_h
    port map (
            O => \N__21872\,
            I => \N__21869\
        );

    \I__5020\ : Odrv4
    port map (
            O => \N__21869\,
            I => \line_buffer.n3650\
        );

    \I__5019\ : InMux
    port map (
            O => \N__21866\,
            I => \N__21863\
        );

    \I__5018\ : LocalMux
    port map (
            O => \N__21863\,
            I => \N__21860\
        );

    \I__5017\ : Span4Mux_v
    port map (
            O => \N__21860\,
            I => \N__21857\
        );

    \I__5016\ : Span4Mux_v
    port map (
            O => \N__21857\,
            I => \N__21854\
        );

    \I__5015\ : Sp12to4
    port map (
            O => \N__21854\,
            I => \N__21851\
        );

    \I__5014\ : Odrv12
    port map (
            O => \N__21851\,
            I => \line_buffer.n570\
        );

    \I__5013\ : InMux
    port map (
            O => \N__21848\,
            I => \N__21845\
        );

    \I__5012\ : LocalMux
    port map (
            O => \N__21845\,
            I => \N__21842\
        );

    \I__5011\ : Span4Mux_v
    port map (
            O => \N__21842\,
            I => \N__21839\
        );

    \I__5010\ : Sp12to4
    port map (
            O => \N__21839\,
            I => \N__21836\
        );

    \I__5009\ : Span12Mux_h
    port map (
            O => \N__21836\,
            I => \N__21833\
        );

    \I__5008\ : Span12Mux_v
    port map (
            O => \N__21833\,
            I => \N__21830\
        );

    \I__5007\ : Odrv12
    port map (
            O => \N__21830\,
            I => \line_buffer.n562\
        );

    \I__5006\ : InMux
    port map (
            O => \N__21827\,
            I => \N__21824\
        );

    \I__5005\ : LocalMux
    port map (
            O => \N__21824\,
            I => \N__21821\
        );

    \I__5004\ : Odrv12
    port map (
            O => \N__21821\,
            I => \line_buffer.n3543\
        );

    \I__5003\ : InMux
    port map (
            O => \N__21818\,
            I => \N__21815\
        );

    \I__5002\ : LocalMux
    port map (
            O => \N__21815\,
            I => \N__21812\
        );

    \I__5001\ : Span4Mux_v
    port map (
            O => \N__21812\,
            I => \N__21809\
        );

    \I__5000\ : Odrv4
    port map (
            O => \N__21809\,
            I => \line_buffer.n3656\
        );

    \I__4999\ : InMux
    port map (
            O => \N__21806\,
            I => \N__21803\
        );

    \I__4998\ : LocalMux
    port map (
            O => \N__21803\,
            I => \N__21800\
        );

    \I__4997\ : Span4Mux_v
    port map (
            O => \N__21800\,
            I => \N__21797\
        );

    \I__4996\ : Sp12to4
    port map (
            O => \N__21797\,
            I => \N__21794\
        );

    \I__4995\ : Odrv12
    port map (
            O => \N__21794\,
            I => \line_buffer.n599\
        );

    \I__4994\ : InMux
    port map (
            O => \N__21791\,
            I => \N__21788\
        );

    \I__4993\ : LocalMux
    port map (
            O => \N__21788\,
            I => \N__21785\
        );

    \I__4992\ : Span12Mux_v
    port map (
            O => \N__21785\,
            I => \N__21782\
        );

    \I__4991\ : Odrv12
    port map (
            O => \N__21782\,
            I => \line_buffer.n591\
        );

    \I__4990\ : InMux
    port map (
            O => \N__21779\,
            I => \N__21776\
        );

    \I__4989\ : LocalMux
    port map (
            O => \N__21776\,
            I => \line_buffer.n3626\
        );

    \I__4988\ : InMux
    port map (
            O => \N__21773\,
            I => \N__21770\
        );

    \I__4987\ : LocalMux
    port map (
            O => \N__21770\,
            I => \N__21767\
        );

    \I__4986\ : Odrv12
    port map (
            O => \N__21767\,
            I => \TX_DATA_2\
        );

    \I__4985\ : IoInMux
    port map (
            O => \N__21764\,
            I => \N__21761\
        );

    \I__4984\ : LocalMux
    port map (
            O => \N__21761\,
            I => \N__21757\
        );

    \I__4983\ : IoInMux
    port map (
            O => \N__21760\,
            I => \N__21754\
        );

    \I__4982\ : Span4Mux_s3_v
    port map (
            O => \N__21757\,
            I => \N__21751\
        );

    \I__4981\ : LocalMux
    port map (
            O => \N__21754\,
            I => \N__21748\
        );

    \I__4980\ : Span4Mux_v
    port map (
            O => \N__21751\,
            I => \N__21744\
        );

    \I__4979\ : IoSpan4Mux
    port map (
            O => \N__21748\,
            I => \N__21741\
        );

    \I__4978\ : IoInMux
    port map (
            O => \N__21747\,
            I => \N__21738\
        );

    \I__4977\ : Span4Mux_v
    port map (
            O => \N__21744\,
            I => \N__21733\
        );

    \I__4976\ : Span4Mux_s3_h
    port map (
            O => \N__21741\,
            I => \N__21733\
        );

    \I__4975\ : LocalMux
    port map (
            O => \N__21738\,
            I => \N__21730\
        );

    \I__4974\ : Span4Mux_h
    port map (
            O => \N__21733\,
            I => \N__21727\
        );

    \I__4973\ : Span4Mux_s3_v
    port map (
            O => \N__21730\,
            I => \N__21724\
        );

    \I__4972\ : Span4Mux_h
    port map (
            O => \N__21727\,
            I => \N__21721\
        );

    \I__4971\ : Span4Mux_v
    port map (
            O => \N__21724\,
            I => \N__21718\
        );

    \I__4970\ : Span4Mux_h
    port map (
            O => \N__21721\,
            I => \N__21713\
        );

    \I__4969\ : Span4Mux_v
    port map (
            O => \N__21718\,
            I => \N__21713\
        );

    \I__4968\ : Odrv4
    port map (
            O => \N__21713\,
            I => n1819
        );

    \I__4967\ : InMux
    port map (
            O => \N__21710\,
            I => \N__21707\
        );

    \I__4966\ : LocalMux
    port map (
            O => \N__21707\,
            I => \line_buffer.n3537\
        );

    \I__4965\ : InMux
    port map (
            O => \N__21704\,
            I => \N__21701\
        );

    \I__4964\ : LocalMux
    port map (
            O => \N__21701\,
            I => \N__21698\
        );

    \I__4963\ : Span12Mux_v
    port map (
            O => \N__21698\,
            I => \N__21695\
        );

    \I__4962\ : Odrv12
    port map (
            O => \N__21695\,
            I => \line_buffer.n3536\
        );

    \I__4961\ : InMux
    port map (
            O => \N__21692\,
            I => \N__21689\
        );

    \I__4960\ : LocalMux
    port map (
            O => \N__21689\,
            I => \line_buffer.n3614\
        );

    \I__4959\ : InMux
    port map (
            O => \N__21686\,
            I => \N__21683\
        );

    \I__4958\ : LocalMux
    port map (
            O => \N__21683\,
            I => \N__21680\
        );

    \I__4957\ : Span12Mux_s10_v
    port map (
            O => \N__21680\,
            I => \N__21677\
        );

    \I__4956\ : Odrv12
    port map (
            O => \N__21677\,
            I => \line_buffer.n469\
        );

    \I__4955\ : InMux
    port map (
            O => \N__21674\,
            I => \N__21671\
        );

    \I__4954\ : LocalMux
    port map (
            O => \N__21671\,
            I => \N__21668\
        );

    \I__4953\ : Span4Mux_v
    port map (
            O => \N__21668\,
            I => \N__21665\
        );

    \I__4952\ : Span4Mux_h
    port map (
            O => \N__21665\,
            I => \N__21662\
        );

    \I__4951\ : Span4Mux_h
    port map (
            O => \N__21662\,
            I => \N__21659\
        );

    \I__4950\ : Odrv4
    port map (
            O => \N__21659\,
            I => \line_buffer.n461\
        );

    \I__4949\ : InMux
    port map (
            O => \N__21656\,
            I => \N__21653\
        );

    \I__4948\ : LocalMux
    port map (
            O => \N__21653\,
            I => \N__21650\
        );

    \I__4947\ : Span12Mux_v
    port map (
            O => \N__21650\,
            I => \N__21647\
        );

    \I__4946\ : Odrv12
    port map (
            O => \N__21647\,
            I => \line_buffer.n3569\
        );

    \I__4945\ : IoInMux
    port map (
            O => \N__21644\,
            I => \N__21641\
        );

    \I__4944\ : LocalMux
    port map (
            O => \N__21641\,
            I => \N__21638\
        );

    \I__4943\ : IoSpan4Mux
    port map (
            O => \N__21638\,
            I => \N__21635\
        );

    \I__4942\ : Span4Mux_s3_h
    port map (
            O => \N__21635\,
            I => \N__21632\
        );

    \I__4941\ : Span4Mux_h
    port map (
            O => \N__21632\,
            I => \N__21629\
        );

    \I__4940\ : Span4Mux_h
    port map (
            O => \N__21629\,
            I => \N__21625\
        );

    \I__4939\ : InMux
    port map (
            O => \N__21628\,
            I => \N__21622\
        );

    \I__4938\ : Span4Mux_h
    port map (
            O => \N__21625\,
            I => \N__21617\
        );

    \I__4937\ : LocalMux
    port map (
            O => \N__21622\,
            I => \N__21617\
        );

    \I__4936\ : Span4Mux_h
    port map (
            O => \N__21617\,
            I => \N__21614\
        );

    \I__4935\ : Sp12to4
    port map (
            O => \N__21614\,
            I => \N__21611\
        );

    \I__4934\ : Odrv12
    port map (
            O => \N__21611\,
            I => \DEBUG_c_2_c\
        );

    \I__4933\ : InMux
    port map (
            O => \N__21608\,
            I => \N__21605\
        );

    \I__4932\ : LocalMux
    port map (
            O => \N__21605\,
            I => \tvp_hs_buffer.BUFFER_0_0\
        );

    \I__4931\ : InMux
    port map (
            O => \N__21602\,
            I => \N__21599\
        );

    \I__4930\ : LocalMux
    port map (
            O => \N__21599\,
            I => \N__21596\
        );

    \I__4929\ : Span4Mux_v
    port map (
            O => \N__21596\,
            I => \N__21593\
        );

    \I__4928\ : Sp12to4
    port map (
            O => \N__21593\,
            I => \N__21590\
        );

    \I__4927\ : Odrv12
    port map (
            O => \N__21590\,
            I => \line_buffer.n598\
        );

    \I__4926\ : InMux
    port map (
            O => \N__21587\,
            I => \N__21584\
        );

    \I__4925\ : LocalMux
    port map (
            O => \N__21584\,
            I => \N__21581\
        );

    \I__4924\ : Span4Mux_v
    port map (
            O => \N__21581\,
            I => \N__21578\
        );

    \I__4923\ : Sp12to4
    port map (
            O => \N__21578\,
            I => \N__21575\
        );

    \I__4922\ : Span12Mux_h
    port map (
            O => \N__21575\,
            I => \N__21572\
        );

    \I__4921\ : Span12Mux_v
    port map (
            O => \N__21572\,
            I => \N__21569\
        );

    \I__4920\ : Odrv12
    port map (
            O => \N__21569\,
            I => \line_buffer.n590\
        );

    \I__4919\ : InMux
    port map (
            O => \N__21566\,
            I => \N__21563\
        );

    \I__4918\ : LocalMux
    port map (
            O => \N__21563\,
            I => \line_buffer.n3573\
        );

    \I__4917\ : InMux
    port map (
            O => \N__21560\,
            I => \N__21557\
        );

    \I__4916\ : LocalMux
    port map (
            O => \N__21557\,
            I => \line_buffer.n3659\
        );

    \I__4915\ : InMux
    port map (
            O => \N__21554\,
            I => \N__21551\
        );

    \I__4914\ : LocalMux
    port map (
            O => \N__21551\,
            I => \N__21548\
        );

    \I__4913\ : Span4Mux_v
    port map (
            O => \N__21548\,
            I => \N__21545\
        );

    \I__4912\ : Span4Mux_v
    port map (
            O => \N__21545\,
            I => \N__21542\
        );

    \I__4911\ : Sp12to4
    port map (
            O => \N__21542\,
            I => \N__21539\
        );

    \I__4910\ : Odrv12
    port map (
            O => \N__21539\,
            I => \line_buffer.n564\
        );

    \I__4909\ : InMux
    port map (
            O => \N__21536\,
            I => \N__21533\
        );

    \I__4908\ : LocalMux
    port map (
            O => \N__21533\,
            I => \N__21530\
        );

    \I__4907\ : Span4Mux_v
    port map (
            O => \N__21530\,
            I => \N__21527\
        );

    \I__4906\ : Span4Mux_h
    port map (
            O => \N__21527\,
            I => \N__21524\
        );

    \I__4905\ : Odrv4
    port map (
            O => \N__21524\,
            I => \line_buffer.n556\
        );

    \I__4904\ : InMux
    port map (
            O => \N__21521\,
            I => \N__21518\
        );

    \I__4903\ : LocalMux
    port map (
            O => \N__21518\,
            I => \N__21515\
        );

    \I__4902\ : Span4Mux_v
    port map (
            O => \N__21515\,
            I => \N__21512\
        );

    \I__4901\ : Span4Mux_h
    port map (
            O => \N__21512\,
            I => \N__21509\
        );

    \I__4900\ : Span4Mux_h
    port map (
            O => \N__21509\,
            I => \N__21506\
        );

    \I__4899\ : Odrv4
    port map (
            O => \N__21506\,
            I => \line_buffer.n534\
        );

    \I__4898\ : InMux
    port map (
            O => \N__21503\,
            I => \N__21500\
        );

    \I__4897\ : LocalMux
    port map (
            O => \N__21500\,
            I => \N__21497\
        );

    \I__4896\ : Odrv12
    port map (
            O => \N__21497\,
            I => \line_buffer.n526\
        );

    \I__4895\ : InMux
    port map (
            O => \N__21494\,
            I => \N__21491\
        );

    \I__4894\ : LocalMux
    port map (
            O => \N__21491\,
            I => \N__21488\
        );

    \I__4893\ : Odrv4
    port map (
            O => \N__21488\,
            I => \transmit_module.X_DELTA_PATTERN_6\
        );

    \I__4892\ : InMux
    port map (
            O => \N__21485\,
            I => \N__21482\
        );

    \I__4891\ : LocalMux
    port map (
            O => \N__21482\,
            I => \N__21479\
        );

    \I__4890\ : Odrv4
    port map (
            O => \N__21479\,
            I => \transmit_module.X_DELTA_PATTERN_5\
        );

    \I__4889\ : CEMux
    port map (
            O => \N__21476\,
            I => \N__21471\
        );

    \I__4888\ : CEMux
    port map (
            O => \N__21475\,
            I => \N__21468\
        );

    \I__4887\ : CEMux
    port map (
            O => \N__21474\,
            I => \N__21465\
        );

    \I__4886\ : LocalMux
    port map (
            O => \N__21471\,
            I => \N__21461\
        );

    \I__4885\ : LocalMux
    port map (
            O => \N__21468\,
            I => \N__21458\
        );

    \I__4884\ : LocalMux
    port map (
            O => \N__21465\,
            I => \N__21455\
        );

    \I__4883\ : CEMux
    port map (
            O => \N__21464\,
            I => \N__21452\
        );

    \I__4882\ : Span4Mux_v
    port map (
            O => \N__21461\,
            I => \N__21449\
        );

    \I__4881\ : Span4Mux_h
    port map (
            O => \N__21458\,
            I => \N__21446\
        );

    \I__4880\ : Span4Mux_h
    port map (
            O => \N__21455\,
            I => \N__21443\
        );

    \I__4879\ : LocalMux
    port map (
            O => \N__21452\,
            I => \N__21440\
        );

    \I__4878\ : Odrv4
    port map (
            O => \N__21449\,
            I => \transmit_module.n2087\
        );

    \I__4877\ : Odrv4
    port map (
            O => \N__21446\,
            I => \transmit_module.n2087\
        );

    \I__4876\ : Odrv4
    port map (
            O => \N__21443\,
            I => \transmit_module.n2087\
        );

    \I__4875\ : Odrv12
    port map (
            O => \N__21440\,
            I => \transmit_module.n2087\
        );

    \I__4874\ : CEMux
    port map (
            O => \N__21431\,
            I => \N__21423\
        );

    \I__4873\ : CEMux
    port map (
            O => \N__21430\,
            I => \N__21420\
        );

    \I__4872\ : CEMux
    port map (
            O => \N__21429\,
            I => \N__21417\
        );

    \I__4871\ : CEMux
    port map (
            O => \N__21428\,
            I => \N__21414\
        );

    \I__4870\ : CEMux
    port map (
            O => \N__21427\,
            I => \N__21411\
        );

    \I__4869\ : CEMux
    port map (
            O => \N__21426\,
            I => \N__21408\
        );

    \I__4868\ : LocalMux
    port map (
            O => \N__21423\,
            I => \N__21402\
        );

    \I__4867\ : LocalMux
    port map (
            O => \N__21420\,
            I => \N__21399\
        );

    \I__4866\ : LocalMux
    port map (
            O => \N__21417\,
            I => \N__21392\
        );

    \I__4865\ : LocalMux
    port map (
            O => \N__21414\,
            I => \N__21392\
        );

    \I__4864\ : LocalMux
    port map (
            O => \N__21411\,
            I => \N__21392\
        );

    \I__4863\ : LocalMux
    port map (
            O => \N__21408\,
            I => \N__21389\
        );

    \I__4862\ : CEMux
    port map (
            O => \N__21407\,
            I => \N__21386\
        );

    \I__4861\ : CEMux
    port map (
            O => \N__21406\,
            I => \N__21383\
        );

    \I__4860\ : CEMux
    port map (
            O => \N__21405\,
            I => \N__21378\
        );

    \I__4859\ : Span4Mux_v
    port map (
            O => \N__21402\,
            I => \N__21373\
        );

    \I__4858\ : Span4Mux_v
    port map (
            O => \N__21399\,
            I => \N__21373\
        );

    \I__4857\ : Span4Mux_v
    port map (
            O => \N__21392\,
            I => \N__21366\
        );

    \I__4856\ : Span4Mux_h
    port map (
            O => \N__21389\,
            I => \N__21366\
        );

    \I__4855\ : LocalMux
    port map (
            O => \N__21386\,
            I => \N__21366\
        );

    \I__4854\ : LocalMux
    port map (
            O => \N__21383\,
            I => \N__21363\
        );

    \I__4853\ : CEMux
    port map (
            O => \N__21382\,
            I => \N__21359\
        );

    \I__4852\ : CEMux
    port map (
            O => \N__21381\,
            I => \N__21356\
        );

    \I__4851\ : LocalMux
    port map (
            O => \N__21378\,
            I => \N__21351\
        );

    \I__4850\ : Span4Mux_h
    port map (
            O => \N__21373\,
            I => \N__21344\
        );

    \I__4849\ : Span4Mux_h
    port map (
            O => \N__21366\,
            I => \N__21344\
        );

    \I__4848\ : Span4Mux_v
    port map (
            O => \N__21363\,
            I => \N__21344\
        );

    \I__4847\ : SRMux
    port map (
            O => \N__21362\,
            I => \N__21341\
        );

    \I__4846\ : LocalMux
    port map (
            O => \N__21359\,
            I => \N__21338\
        );

    \I__4845\ : LocalMux
    port map (
            O => \N__21356\,
            I => \N__21335\
        );

    \I__4844\ : SRMux
    port map (
            O => \N__21355\,
            I => \N__21332\
        );

    \I__4843\ : SRMux
    port map (
            O => \N__21354\,
            I => \N__21328\
        );

    \I__4842\ : Span4Mux_v
    port map (
            O => \N__21351\,
            I => \N__21322\
        );

    \I__4841\ : Span4Mux_h
    port map (
            O => \N__21344\,
            I => \N__21322\
        );

    \I__4840\ : LocalMux
    port map (
            O => \N__21341\,
            I => \N__21319\
        );

    \I__4839\ : Span4Mux_h
    port map (
            O => \N__21338\,
            I => \N__21312\
        );

    \I__4838\ : Span4Mux_v
    port map (
            O => \N__21335\,
            I => \N__21312\
        );

    \I__4837\ : LocalMux
    port map (
            O => \N__21332\,
            I => \N__21312\
        );

    \I__4836\ : CEMux
    port map (
            O => \N__21331\,
            I => \N__21309\
        );

    \I__4835\ : LocalMux
    port map (
            O => \N__21328\,
            I => \N__21306\
        );

    \I__4834\ : SRMux
    port map (
            O => \N__21327\,
            I => \N__21303\
        );

    \I__4833\ : Span4Mux_h
    port map (
            O => \N__21322\,
            I => \N__21300\
        );

    \I__4832\ : Span4Mux_h
    port map (
            O => \N__21319\,
            I => \N__21297\
        );

    \I__4831\ : Span4Mux_h
    port map (
            O => \N__21312\,
            I => \N__21294\
        );

    \I__4830\ : LocalMux
    port map (
            O => \N__21309\,
            I => \N__21287\
        );

    \I__4829\ : Sp12to4
    port map (
            O => \N__21306\,
            I => \N__21287\
        );

    \I__4828\ : LocalMux
    port map (
            O => \N__21303\,
            I => \N__21287\
        );

    \I__4827\ : Odrv4
    port map (
            O => \N__21300\,
            I => \transmit_module.n3682\
        );

    \I__4826\ : Odrv4
    port map (
            O => \N__21297\,
            I => \transmit_module.n3682\
        );

    \I__4825\ : Odrv4
    port map (
            O => \N__21294\,
            I => \transmit_module.n3682\
        );

    \I__4824\ : Odrv12
    port map (
            O => \N__21287\,
            I => \transmit_module.n3682\
        );

    \I__4823\ : InMux
    port map (
            O => \N__21278\,
            I => \N__21275\
        );

    \I__4822\ : LocalMux
    port map (
            O => \N__21275\,
            I => \N__21272\
        );

    \I__4821\ : Span4Mux_h
    port map (
            O => \N__21272\,
            I => \N__21269\
        );

    \I__4820\ : Sp12to4
    port map (
            O => \N__21269\,
            I => \N__21266\
        );

    \I__4819\ : Span12Mux_v
    port map (
            O => \N__21266\,
            I => \N__21263\
        );

    \I__4818\ : Odrv12
    port map (
            O => \N__21263\,
            I => \line_buffer.n533\
        );

    \I__4817\ : CascadeMux
    port map (
            O => \N__21260\,
            I => \N__21257\
        );

    \I__4816\ : InMux
    port map (
            O => \N__21257\,
            I => \N__21254\
        );

    \I__4815\ : LocalMux
    port map (
            O => \N__21254\,
            I => \N__21251\
        );

    \I__4814\ : Span4Mux_v
    port map (
            O => \N__21251\,
            I => \N__21248\
        );

    \I__4813\ : Span4Mux_h
    port map (
            O => \N__21248\,
            I => \N__21245\
        );

    \I__4812\ : Odrv4
    port map (
            O => \N__21245\,
            I => \line_buffer.n525\
        );

    \I__4811\ : InMux
    port map (
            O => \N__21242\,
            I => \N__21239\
        );

    \I__4810\ : LocalMux
    port map (
            O => \N__21239\,
            I => \line_buffer.n3653\
        );

    \I__4809\ : InMux
    port map (
            O => \N__21236\,
            I => \N__21233\
        );

    \I__4808\ : LocalMux
    port map (
            O => \N__21233\,
            I => \N__21230\
        );

    \I__4807\ : Span12Mux_v
    port map (
            O => \N__21230\,
            I => \N__21227\
        );

    \I__4806\ : Odrv12
    port map (
            O => \N__21227\,
            I => \line_buffer.n468\
        );

    \I__4805\ : CascadeMux
    port map (
            O => \N__21224\,
            I => \N__21221\
        );

    \I__4804\ : InMux
    port map (
            O => \N__21221\,
            I => \N__21218\
        );

    \I__4803\ : LocalMux
    port map (
            O => \N__21218\,
            I => \N__21215\
        );

    \I__4802\ : Span12Mux_v
    port map (
            O => \N__21215\,
            I => \N__21212\
        );

    \I__4801\ : Odrv12
    port map (
            O => \N__21212\,
            I => \line_buffer.n460\
        );

    \I__4800\ : InMux
    port map (
            O => \N__21209\,
            I => \N__21206\
        );

    \I__4799\ : LocalMux
    port map (
            O => \N__21206\,
            I => \line_buffer.n3635\
        );

    \I__4798\ : InMux
    port map (
            O => \N__21203\,
            I => \N__21200\
        );

    \I__4797\ : LocalMux
    port map (
            O => \N__21200\,
            I => \N__21197\
        );

    \I__4796\ : Span4Mux_v
    port map (
            O => \N__21197\,
            I => \N__21194\
        );

    \I__4795\ : Span4Mux_h
    port map (
            O => \N__21194\,
            I => \N__21191\
        );

    \I__4794\ : Span4Mux_h
    port map (
            O => \N__21191\,
            I => \N__21188\
        );

    \I__4793\ : Odrv4
    port map (
            O => \N__21188\,
            I => \line_buffer.n566\
        );

    \I__4792\ : InMux
    port map (
            O => \N__21185\,
            I => \N__21182\
        );

    \I__4791\ : LocalMux
    port map (
            O => \N__21182\,
            I => \N__21179\
        );

    \I__4790\ : Odrv12
    port map (
            O => \N__21179\,
            I => \line_buffer.n558\
        );

    \I__4789\ : InMux
    port map (
            O => \N__21176\,
            I => \N__21173\
        );

    \I__4788\ : LocalMux
    port map (
            O => \N__21173\,
            I => \N__21170\
        );

    \I__4787\ : Odrv12
    port map (
            O => \N__21170\,
            I => \line_buffer.n557\
        );

    \I__4786\ : InMux
    port map (
            O => \N__21167\,
            I => \N__21164\
        );

    \I__4785\ : LocalMux
    port map (
            O => \N__21164\,
            I => \N__21161\
        );

    \I__4784\ : Span4Mux_v
    port map (
            O => \N__21161\,
            I => \N__21158\
        );

    \I__4783\ : Span4Mux_h
    port map (
            O => \N__21158\,
            I => \N__21155\
        );

    \I__4782\ : Span4Mux_h
    port map (
            O => \N__21155\,
            I => \N__21152\
        );

    \I__4781\ : Odrv4
    port map (
            O => \N__21152\,
            I => \line_buffer.n565\
        );

    \I__4780\ : InMux
    port map (
            O => \N__21149\,
            I => \N__21146\
        );

    \I__4779\ : LocalMux
    port map (
            O => \N__21146\,
            I => \line_buffer.n3632\
        );

    \I__4778\ : InMux
    port map (
            O => \N__21143\,
            I => \N__21140\
        );

    \I__4777\ : LocalMux
    port map (
            O => \N__21140\,
            I => \N__21137\
        );

    \I__4776\ : Span4Mux_v
    port map (
            O => \N__21137\,
            I => \N__21134\
        );

    \I__4775\ : Odrv4
    port map (
            O => \N__21134\,
            I => \line_buffer.n3572\
        );

    \I__4774\ : CascadeMux
    port map (
            O => \N__21131\,
            I => \line_buffer.n3602_cascade_\
        );

    \I__4773\ : InMux
    port map (
            O => \N__21128\,
            I => \N__21125\
        );

    \I__4772\ : LocalMux
    port map (
            O => \N__21125\,
            I => \line_buffer.n3570\
        );

    \I__4771\ : InMux
    port map (
            O => \N__21122\,
            I => \N__21119\
        );

    \I__4770\ : LocalMux
    port map (
            O => \N__21119\,
            I => \N__21116\
        );

    \I__4769\ : Span4Mux_h
    port map (
            O => \N__21116\,
            I => \N__21113\
        );

    \I__4768\ : Span4Mux_h
    port map (
            O => \N__21113\,
            I => \N__21110\
        );

    \I__4767\ : Odrv4
    port map (
            O => \N__21110\,
            I => \line_buffer.n472\
        );

    \I__4766\ : CascadeMux
    port map (
            O => \N__21107\,
            I => \N__21104\
        );

    \I__4765\ : InMux
    port map (
            O => \N__21104\,
            I => \N__21101\
        );

    \I__4764\ : LocalMux
    port map (
            O => \N__21101\,
            I => \N__21098\
        );

    \I__4763\ : Span4Mux_v
    port map (
            O => \N__21098\,
            I => \N__21095\
        );

    \I__4762\ : Sp12to4
    port map (
            O => \N__21095\,
            I => \N__21092\
        );

    \I__4761\ : Span12Mux_h
    port map (
            O => \N__21092\,
            I => \N__21089\
        );

    \I__4760\ : Odrv12
    port map (
            O => \N__21089\,
            I => \line_buffer.n464\
        );

    \I__4759\ : CascadeMux
    port map (
            O => \N__21086\,
            I => \line_buffer.n3593_cascade_\
        );

    \I__4758\ : InMux
    port map (
            O => \N__21083\,
            I => \N__21080\
        );

    \I__4757\ : LocalMux
    port map (
            O => \N__21080\,
            I => \N__21077\
        );

    \I__4756\ : Odrv4
    port map (
            O => \N__21077\,
            I => \line_buffer.n3629\
        );

    \I__4755\ : InMux
    port map (
            O => \N__21074\,
            I => \N__21071\
        );

    \I__4754\ : LocalMux
    port map (
            O => \N__21071\,
            I => \TX_DATA_3\
        );

    \I__4753\ : InMux
    port map (
            O => \N__21068\,
            I => \N__21065\
        );

    \I__4752\ : LocalMux
    port map (
            O => \N__21065\,
            I => \N__21062\
        );

    \I__4751\ : Span4Mux_v
    port map (
            O => \N__21062\,
            I => \N__21059\
        );

    \I__4750\ : Sp12to4
    port map (
            O => \N__21059\,
            I => \N__21056\
        );

    \I__4749\ : Odrv12
    port map (
            O => \N__21056\,
            I => \line_buffer.n471\
        );

    \I__4748\ : InMux
    port map (
            O => \N__21053\,
            I => \N__21050\
        );

    \I__4747\ : LocalMux
    port map (
            O => \N__21050\,
            I => \N__21047\
        );

    \I__4746\ : Span4Mux_h
    port map (
            O => \N__21047\,
            I => \N__21044\
        );

    \I__4745\ : Span4Mux_v
    port map (
            O => \N__21044\,
            I => \N__21041\
        );

    \I__4744\ : Span4Mux_h
    port map (
            O => \N__21041\,
            I => \N__21038\
        );

    \I__4743\ : Odrv4
    port map (
            O => \N__21038\,
            I => \line_buffer.n463\
        );

    \I__4742\ : InMux
    port map (
            O => \N__21035\,
            I => \N__21032\
        );

    \I__4741\ : LocalMux
    port map (
            O => \N__21032\,
            I => \N__21029\
        );

    \I__4740\ : Span4Mux_v
    port map (
            O => \N__21029\,
            I => \N__21026\
        );

    \I__4739\ : Span4Mux_v
    port map (
            O => \N__21026\,
            I => \N__21023\
        );

    \I__4738\ : Odrv4
    port map (
            O => \N__21023\,
            I => \line_buffer.n3552\
        );

    \I__4737\ : CascadeMux
    port map (
            O => \N__21020\,
            I => \line_buffer.n3551_cascade_\
        );

    \I__4736\ : InMux
    port map (
            O => \N__21017\,
            I => \N__21014\
        );

    \I__4735\ : LocalMux
    port map (
            O => \N__21014\,
            I => \N__21011\
        );

    \I__4734\ : Span4Mux_v
    port map (
            O => \N__21011\,
            I => \N__21008\
        );

    \I__4733\ : Span4Mux_h
    port map (
            O => \N__21008\,
            I => \N__21005\
        );

    \I__4732\ : Span4Mux_h
    port map (
            O => \N__21005\,
            I => \N__21002\
        );

    \I__4731\ : Span4Mux_v
    port map (
            O => \N__21002\,
            I => \N__20999\
        );

    \I__4730\ : Odrv4
    port map (
            O => \N__20999\,
            I => \line_buffer.n600\
        );

    \I__4729\ : InMux
    port map (
            O => \N__20996\,
            I => \N__20993\
        );

    \I__4728\ : LocalMux
    port map (
            O => \N__20993\,
            I => \N__20990\
        );

    \I__4727\ : Span4Mux_v
    port map (
            O => \N__20990\,
            I => \N__20987\
        );

    \I__4726\ : Span4Mux_h
    port map (
            O => \N__20987\,
            I => \N__20984\
        );

    \I__4725\ : Span4Mux_h
    port map (
            O => \N__20984\,
            I => \N__20981\
        );

    \I__4724\ : Odrv4
    port map (
            O => \N__20981\,
            I => \line_buffer.n592\
        );

    \I__4723\ : InMux
    port map (
            O => \N__20978\,
            I => \N__20975\
        );

    \I__4722\ : LocalMux
    port map (
            O => \N__20975\,
            I => \N__20972\
        );

    \I__4721\ : Odrv4
    port map (
            O => \N__20972\,
            I => \TX_DATA_4\
        );

    \I__4720\ : IoInMux
    port map (
            O => \N__20969\,
            I => \N__20966\
        );

    \I__4719\ : LocalMux
    port map (
            O => \N__20966\,
            I => \N__20961\
        );

    \I__4718\ : IoInMux
    port map (
            O => \N__20965\,
            I => \N__20958\
        );

    \I__4717\ : IoInMux
    port map (
            O => \N__20964\,
            I => \N__20955\
        );

    \I__4716\ : IoSpan4Mux
    port map (
            O => \N__20961\,
            I => \N__20952\
        );

    \I__4715\ : LocalMux
    port map (
            O => \N__20958\,
            I => \N__20949\
        );

    \I__4714\ : LocalMux
    port map (
            O => \N__20955\,
            I => \N__20946\
        );

    \I__4713\ : Span4Mux_s0_v
    port map (
            O => \N__20952\,
            I => \N__20943\
        );

    \I__4712\ : IoSpan4Mux
    port map (
            O => \N__20949\,
            I => \N__20940\
        );

    \I__4711\ : IoSpan4Mux
    port map (
            O => \N__20946\,
            I => \N__20937\
        );

    \I__4710\ : Span4Mux_v
    port map (
            O => \N__20943\,
            I => \N__20934\
        );

    \I__4709\ : Span4Mux_s3_h
    port map (
            O => \N__20940\,
            I => \N__20931\
        );

    \I__4708\ : Span4Mux_s2_v
    port map (
            O => \N__20937\,
            I => \N__20928\
        );

    \I__4707\ : Span4Mux_v
    port map (
            O => \N__20934\,
            I => \N__20923\
        );

    \I__4706\ : Span4Mux_h
    port map (
            O => \N__20931\,
            I => \N__20923\
        );

    \I__4705\ : Sp12to4
    port map (
            O => \N__20928\,
            I => \N__20920\
        );

    \I__4704\ : Span4Mux_h
    port map (
            O => \N__20923\,
            I => \N__20917\
        );

    \I__4703\ : Span12Mux_s8_v
    port map (
            O => \N__20920\,
            I => \N__20914\
        );

    \I__4702\ : Span4Mux_h
    port map (
            O => \N__20917\,
            I => \N__20911\
        );

    \I__4701\ : Odrv12
    port map (
            O => \N__20914\,
            I => n1817
        );

    \I__4700\ : Odrv4
    port map (
            O => \N__20911\,
            I => n1817
        );

    \I__4699\ : InMux
    port map (
            O => \N__20906\,
            I => \N__20903\
        );

    \I__4698\ : LocalMux
    port map (
            O => \N__20903\,
            I => \N__20900\
        );

    \I__4697\ : Span12Mux_s10_v
    port map (
            O => \N__20900\,
            I => \N__20897\
        );

    \I__4696\ : Odrv12
    port map (
            O => \N__20897\,
            I => \TX_DATA_1\
        );

    \I__4695\ : IoInMux
    port map (
            O => \N__20894\,
            I => \N__20891\
        );

    \I__4694\ : LocalMux
    port map (
            O => \N__20891\,
            I => \N__20887\
        );

    \I__4693\ : IoInMux
    port map (
            O => \N__20890\,
            I => \N__20884\
        );

    \I__4692\ : IoSpan4Mux
    port map (
            O => \N__20887\,
            I => \N__20879\
        );

    \I__4691\ : LocalMux
    port map (
            O => \N__20884\,
            I => \N__20879\
        );

    \I__4690\ : IoSpan4Mux
    port map (
            O => \N__20879\,
            I => \N__20876\
        );

    \I__4689\ : Span4Mux_s2_h
    port map (
            O => \N__20876\,
            I => \N__20872\
        );

    \I__4688\ : IoInMux
    port map (
            O => \N__20875\,
            I => \N__20869\
        );

    \I__4687\ : Span4Mux_h
    port map (
            O => \N__20872\,
            I => \N__20866\
        );

    \I__4686\ : LocalMux
    port map (
            O => \N__20869\,
            I => \N__20863\
        );

    \I__4685\ : Span4Mux_h
    port map (
            O => \N__20866\,
            I => \N__20860\
        );

    \I__4684\ : Span4Mux_s3_v
    port map (
            O => \N__20863\,
            I => \N__20857\
        );

    \I__4683\ : Span4Mux_h
    port map (
            O => \N__20860\,
            I => \N__20852\
        );

    \I__4682\ : Span4Mux_v
    port map (
            O => \N__20857\,
            I => \N__20852\
        );

    \I__4681\ : Odrv4
    port map (
            O => \N__20852\,
            I => n1820
        );

    \I__4680\ : InMux
    port map (
            O => \N__20849\,
            I => \N__20846\
        );

    \I__4679\ : LocalMux
    port map (
            O => \N__20846\,
            I => \N__20843\
        );

    \I__4678\ : Odrv4
    port map (
            O => \N__20843\,
            I => \tvp_hs_buffer.BUFFER_1_0\
        );

    \I__4677\ : InMux
    port map (
            O => \N__20840\,
            I => \N__20837\
        );

    \I__4676\ : LocalMux
    port map (
            O => \N__20837\,
            I => \N__20834\
        );

    \I__4675\ : Span4Mux_v
    port map (
            O => \N__20834\,
            I => \N__20831\
        );

    \I__4674\ : Span4Mux_h
    port map (
            O => \N__20831\,
            I => \N__20828\
        );

    \I__4673\ : Span4Mux_h
    port map (
            O => \N__20828\,
            I => \N__20825\
        );

    \I__4672\ : Odrv4
    port map (
            O => \N__20825\,
            I => \line_buffer.n536\
        );

    \I__4671\ : InMux
    port map (
            O => \N__20822\,
            I => \N__20819\
        );

    \I__4670\ : LocalMux
    port map (
            O => \N__20819\,
            I => \N__20816\
        );

    \I__4669\ : Span12Mux_v
    port map (
            O => \N__20816\,
            I => \N__20813\
        );

    \I__4668\ : Odrv12
    port map (
            O => \N__20813\,
            I => \line_buffer.n528\
        );

    \I__4667\ : InMux
    port map (
            O => \N__20810\,
            I => \N__20807\
        );

    \I__4666\ : LocalMux
    port map (
            O => \N__20807\,
            I => \N__20801\
        );

    \I__4665\ : InMux
    port map (
            O => \N__20806\,
            I => \N__20798\
        );

    \I__4664\ : InMux
    port map (
            O => \N__20805\,
            I => \N__20795\
        );

    \I__4663\ : InMux
    port map (
            O => \N__20804\,
            I => \N__20792\
        );

    \I__4662\ : Odrv12
    port map (
            O => \N__20801\,
            I => \transmit_module.TX_ADDR_4\
        );

    \I__4661\ : LocalMux
    port map (
            O => \N__20798\,
            I => \transmit_module.TX_ADDR_4\
        );

    \I__4660\ : LocalMux
    port map (
            O => \N__20795\,
            I => \transmit_module.TX_ADDR_4\
        );

    \I__4659\ : LocalMux
    port map (
            O => \N__20792\,
            I => \transmit_module.TX_ADDR_4\
        );

    \I__4658\ : InMux
    port map (
            O => \N__20783\,
            I => \N__20780\
        );

    \I__4657\ : LocalMux
    port map (
            O => \N__20780\,
            I => \N__20777\
        );

    \I__4656\ : Odrv4
    port map (
            O => \N__20777\,
            I => \transmit_module.ADDR_Y_COMPONENT_4\
        );

    \I__4655\ : CEMux
    port map (
            O => \N__20774\,
            I => \N__20768\
        );

    \I__4654\ : CEMux
    port map (
            O => \N__20773\,
            I => \N__20765\
        );

    \I__4653\ : CEMux
    port map (
            O => \N__20772\,
            I => \N__20761\
        );

    \I__4652\ : CEMux
    port map (
            O => \N__20771\,
            I => \N__20758\
        );

    \I__4651\ : LocalMux
    port map (
            O => \N__20768\,
            I => \N__20752\
        );

    \I__4650\ : LocalMux
    port map (
            O => \N__20765\,
            I => \N__20752\
        );

    \I__4649\ : CEMux
    port map (
            O => \N__20764\,
            I => \N__20749\
        );

    \I__4648\ : LocalMux
    port map (
            O => \N__20761\,
            I => \N__20745\
        );

    \I__4647\ : LocalMux
    port map (
            O => \N__20758\,
            I => \N__20742\
        );

    \I__4646\ : CEMux
    port map (
            O => \N__20757\,
            I => \N__20739\
        );

    \I__4645\ : Span4Mux_h
    port map (
            O => \N__20752\,
            I => \N__20735\
        );

    \I__4644\ : LocalMux
    port map (
            O => \N__20749\,
            I => \N__20732\
        );

    \I__4643\ : CEMux
    port map (
            O => \N__20748\,
            I => \N__20729\
        );

    \I__4642\ : Span4Mux_v
    port map (
            O => \N__20745\,
            I => \N__20724\
        );

    \I__4641\ : Span4Mux_h
    port map (
            O => \N__20742\,
            I => \N__20724\
        );

    \I__4640\ : LocalMux
    port map (
            O => \N__20739\,
            I => \N__20721\
        );

    \I__4639\ : CEMux
    port map (
            O => \N__20738\,
            I => \N__20718\
        );

    \I__4638\ : Span4Mux_v
    port map (
            O => \N__20735\,
            I => \N__20713\
        );

    \I__4637\ : Span4Mux_h
    port map (
            O => \N__20732\,
            I => \N__20713\
        );

    \I__4636\ : LocalMux
    port map (
            O => \N__20729\,
            I => \N__20710\
        );

    \I__4635\ : Span4Mux_h
    port map (
            O => \N__20724\,
            I => \N__20707\
        );

    \I__4634\ : Span4Mux_h
    port map (
            O => \N__20721\,
            I => \N__20704\
        );

    \I__4633\ : LocalMux
    port map (
            O => \N__20718\,
            I => \N__20701\
        );

    \I__4632\ : Odrv4
    port map (
            O => \N__20713\,
            I => \transmit_module.n2313\
        );

    \I__4631\ : Odrv12
    port map (
            O => \N__20710\,
            I => \transmit_module.n2313\
        );

    \I__4630\ : Odrv4
    port map (
            O => \N__20707\,
            I => \transmit_module.n2313\
        );

    \I__4629\ : Odrv4
    port map (
            O => \N__20704\,
            I => \transmit_module.n2313\
        );

    \I__4628\ : Odrv4
    port map (
            O => \N__20701\,
            I => \transmit_module.n2313\
        );

    \I__4627\ : InMux
    port map (
            O => \N__20690\,
            I => \N__20687\
        );

    \I__4626\ : LocalMux
    port map (
            O => \N__20687\,
            I => \transmit_module.ADDR_Y_COMPONENT_2\
        );

    \I__4625\ : InMux
    port map (
            O => \N__20684\,
            I => \N__20679\
        );

    \I__4624\ : InMux
    port map (
            O => \N__20683\,
            I => \N__20673\
        );

    \I__4623\ : InMux
    port map (
            O => \N__20682\,
            I => \N__20668\
        );

    \I__4622\ : LocalMux
    port map (
            O => \N__20679\,
            I => \N__20665\
        );

    \I__4621\ : InMux
    port map (
            O => \N__20678\,
            I => \N__20662\
        );

    \I__4620\ : InMux
    port map (
            O => \N__20677\,
            I => \N__20656\
        );

    \I__4619\ : InMux
    port map (
            O => \N__20676\,
            I => \N__20656\
        );

    \I__4618\ : LocalMux
    port map (
            O => \N__20673\,
            I => \N__20652\
        );

    \I__4617\ : InMux
    port map (
            O => \N__20672\,
            I => \N__20649\
        );

    \I__4616\ : InMux
    port map (
            O => \N__20671\,
            I => \N__20644\
        );

    \I__4615\ : LocalMux
    port map (
            O => \N__20668\,
            I => \N__20641\
        );

    \I__4614\ : Span4Mux_h
    port map (
            O => \N__20665\,
            I => \N__20636\
        );

    \I__4613\ : LocalMux
    port map (
            O => \N__20662\,
            I => \N__20636\
        );

    \I__4612\ : InMux
    port map (
            O => \N__20661\,
            I => \N__20633\
        );

    \I__4611\ : LocalMux
    port map (
            O => \N__20656\,
            I => \N__20630\
        );

    \I__4610\ : InMux
    port map (
            O => \N__20655\,
            I => \N__20627\
        );

    \I__4609\ : Span4Mux_h
    port map (
            O => \N__20652\,
            I => \N__20620\
        );

    \I__4608\ : LocalMux
    port map (
            O => \N__20649\,
            I => \N__20620\
        );

    \I__4607\ : InMux
    port map (
            O => \N__20648\,
            I => \N__20615\
        );

    \I__4606\ : InMux
    port map (
            O => \N__20647\,
            I => \N__20615\
        );

    \I__4605\ : LocalMux
    port map (
            O => \N__20644\,
            I => \N__20612\
        );

    \I__4604\ : Span4Mux_v
    port map (
            O => \N__20641\,
            I => \N__20605\
        );

    \I__4603\ : Span4Mux_v
    port map (
            O => \N__20636\,
            I => \N__20605\
        );

    \I__4602\ : LocalMux
    port map (
            O => \N__20633\,
            I => \N__20605\
        );

    \I__4601\ : Span4Mux_v
    port map (
            O => \N__20630\,
            I => \N__20600\
        );

    \I__4600\ : LocalMux
    port map (
            O => \N__20627\,
            I => \N__20600\
        );

    \I__4599\ : InMux
    port map (
            O => \N__20626\,
            I => \N__20597\
        );

    \I__4598\ : InMux
    port map (
            O => \N__20625\,
            I => \N__20594\
        );

    \I__4597\ : Odrv4
    port map (
            O => \N__20620\,
            I => \transmit_module.Y_DELTA_PATTERN_0\
        );

    \I__4596\ : LocalMux
    port map (
            O => \N__20615\,
            I => \transmit_module.Y_DELTA_PATTERN_0\
        );

    \I__4595\ : Odrv4
    port map (
            O => \N__20612\,
            I => \transmit_module.Y_DELTA_PATTERN_0\
        );

    \I__4594\ : Odrv4
    port map (
            O => \N__20605\,
            I => \transmit_module.Y_DELTA_PATTERN_0\
        );

    \I__4593\ : Odrv4
    port map (
            O => \N__20600\,
            I => \transmit_module.Y_DELTA_PATTERN_0\
        );

    \I__4592\ : LocalMux
    port map (
            O => \N__20597\,
            I => \transmit_module.Y_DELTA_PATTERN_0\
        );

    \I__4591\ : LocalMux
    port map (
            O => \N__20594\,
            I => \transmit_module.Y_DELTA_PATTERN_0\
        );

    \I__4590\ : InMux
    port map (
            O => \N__20579\,
            I => \N__20574\
        );

    \I__4589\ : InMux
    port map (
            O => \N__20578\,
            I => \N__20570\
        );

    \I__4588\ : InMux
    port map (
            O => \N__20577\,
            I => \N__20567\
        );

    \I__4587\ : LocalMux
    port map (
            O => \N__20574\,
            I => \N__20564\
        );

    \I__4586\ : InMux
    port map (
            O => \N__20573\,
            I => \N__20561\
        );

    \I__4585\ : LocalMux
    port map (
            O => \N__20570\,
            I => \transmit_module.TX_ADDR_2\
        );

    \I__4584\ : LocalMux
    port map (
            O => \N__20567\,
            I => \transmit_module.TX_ADDR_2\
        );

    \I__4583\ : Odrv4
    port map (
            O => \N__20564\,
            I => \transmit_module.TX_ADDR_2\
        );

    \I__4582\ : LocalMux
    port map (
            O => \N__20561\,
            I => \transmit_module.TX_ADDR_2\
        );

    \I__4581\ : InMux
    port map (
            O => \N__20552\,
            I => \N__20549\
        );

    \I__4580\ : LocalMux
    port map (
            O => \N__20549\,
            I => \N__20545\
        );

    \I__4579\ : InMux
    port map (
            O => \N__20548\,
            I => \N__20542\
        );

    \I__4578\ : Odrv4
    port map (
            O => \N__20545\,
            I => \transmit_module.n114\
        );

    \I__4577\ : LocalMux
    port map (
            O => \N__20542\,
            I => \transmit_module.n114\
        );

    \I__4576\ : InMux
    port map (
            O => \N__20537\,
            I => \N__20534\
        );

    \I__4575\ : LocalMux
    port map (
            O => \N__20534\,
            I => \N__20531\
        );

    \I__4574\ : Odrv4
    port map (
            O => \N__20531\,
            I => \transmit_module.n145\
        );

    \I__4573\ : CascadeMux
    port map (
            O => \N__20528\,
            I => \N__20524\
        );

    \I__4572\ : CascadeMux
    port map (
            O => \N__20527\,
            I => \N__20521\
        );

    \I__4571\ : CascadeBuf
    port map (
            O => \N__20524\,
            I => \N__20518\
        );

    \I__4570\ : CascadeBuf
    port map (
            O => \N__20521\,
            I => \N__20515\
        );

    \I__4569\ : CascadeMux
    port map (
            O => \N__20518\,
            I => \N__20512\
        );

    \I__4568\ : CascadeMux
    port map (
            O => \N__20515\,
            I => \N__20509\
        );

    \I__4567\ : CascadeBuf
    port map (
            O => \N__20512\,
            I => \N__20506\
        );

    \I__4566\ : CascadeBuf
    port map (
            O => \N__20509\,
            I => \N__20503\
        );

    \I__4565\ : CascadeMux
    port map (
            O => \N__20506\,
            I => \N__20500\
        );

    \I__4564\ : CascadeMux
    port map (
            O => \N__20503\,
            I => \N__20497\
        );

    \I__4563\ : CascadeBuf
    port map (
            O => \N__20500\,
            I => \N__20494\
        );

    \I__4562\ : CascadeBuf
    port map (
            O => \N__20497\,
            I => \N__20491\
        );

    \I__4561\ : CascadeMux
    port map (
            O => \N__20494\,
            I => \N__20488\
        );

    \I__4560\ : CascadeMux
    port map (
            O => \N__20491\,
            I => \N__20485\
        );

    \I__4559\ : CascadeBuf
    port map (
            O => \N__20488\,
            I => \N__20482\
        );

    \I__4558\ : CascadeBuf
    port map (
            O => \N__20485\,
            I => \N__20479\
        );

    \I__4557\ : CascadeMux
    port map (
            O => \N__20482\,
            I => \N__20476\
        );

    \I__4556\ : CascadeMux
    port map (
            O => \N__20479\,
            I => \N__20473\
        );

    \I__4555\ : CascadeBuf
    port map (
            O => \N__20476\,
            I => \N__20470\
        );

    \I__4554\ : CascadeBuf
    port map (
            O => \N__20473\,
            I => \N__20467\
        );

    \I__4553\ : CascadeMux
    port map (
            O => \N__20470\,
            I => \N__20464\
        );

    \I__4552\ : CascadeMux
    port map (
            O => \N__20467\,
            I => \N__20461\
        );

    \I__4551\ : CascadeBuf
    port map (
            O => \N__20464\,
            I => \N__20458\
        );

    \I__4550\ : CascadeBuf
    port map (
            O => \N__20461\,
            I => \N__20455\
        );

    \I__4549\ : CascadeMux
    port map (
            O => \N__20458\,
            I => \N__20452\
        );

    \I__4548\ : CascadeMux
    port map (
            O => \N__20455\,
            I => \N__20449\
        );

    \I__4547\ : CascadeBuf
    port map (
            O => \N__20452\,
            I => \N__20446\
        );

    \I__4546\ : CascadeBuf
    port map (
            O => \N__20449\,
            I => \N__20443\
        );

    \I__4545\ : CascadeMux
    port map (
            O => \N__20446\,
            I => \N__20440\
        );

    \I__4544\ : CascadeMux
    port map (
            O => \N__20443\,
            I => \N__20437\
        );

    \I__4543\ : CascadeBuf
    port map (
            O => \N__20440\,
            I => \N__20434\
        );

    \I__4542\ : CascadeBuf
    port map (
            O => \N__20437\,
            I => \N__20431\
        );

    \I__4541\ : CascadeMux
    port map (
            O => \N__20434\,
            I => \N__20428\
        );

    \I__4540\ : CascadeMux
    port map (
            O => \N__20431\,
            I => \N__20425\
        );

    \I__4539\ : CascadeBuf
    port map (
            O => \N__20428\,
            I => \N__20422\
        );

    \I__4538\ : CascadeBuf
    port map (
            O => \N__20425\,
            I => \N__20419\
        );

    \I__4537\ : CascadeMux
    port map (
            O => \N__20422\,
            I => \N__20416\
        );

    \I__4536\ : CascadeMux
    port map (
            O => \N__20419\,
            I => \N__20413\
        );

    \I__4535\ : CascadeBuf
    port map (
            O => \N__20416\,
            I => \N__20410\
        );

    \I__4534\ : CascadeBuf
    port map (
            O => \N__20413\,
            I => \N__20407\
        );

    \I__4533\ : CascadeMux
    port map (
            O => \N__20410\,
            I => \N__20404\
        );

    \I__4532\ : CascadeMux
    port map (
            O => \N__20407\,
            I => \N__20401\
        );

    \I__4531\ : CascadeBuf
    port map (
            O => \N__20404\,
            I => \N__20398\
        );

    \I__4530\ : CascadeBuf
    port map (
            O => \N__20401\,
            I => \N__20395\
        );

    \I__4529\ : CascadeMux
    port map (
            O => \N__20398\,
            I => \N__20392\
        );

    \I__4528\ : CascadeMux
    port map (
            O => \N__20395\,
            I => \N__20389\
        );

    \I__4527\ : CascadeBuf
    port map (
            O => \N__20392\,
            I => \N__20386\
        );

    \I__4526\ : CascadeBuf
    port map (
            O => \N__20389\,
            I => \N__20383\
        );

    \I__4525\ : CascadeMux
    port map (
            O => \N__20386\,
            I => \N__20380\
        );

    \I__4524\ : CascadeMux
    port map (
            O => \N__20383\,
            I => \N__20377\
        );

    \I__4523\ : CascadeBuf
    port map (
            O => \N__20380\,
            I => \N__20374\
        );

    \I__4522\ : CascadeBuf
    port map (
            O => \N__20377\,
            I => \N__20371\
        );

    \I__4521\ : CascadeMux
    port map (
            O => \N__20374\,
            I => \N__20368\
        );

    \I__4520\ : CascadeMux
    port map (
            O => \N__20371\,
            I => \N__20365\
        );

    \I__4519\ : CascadeBuf
    port map (
            O => \N__20368\,
            I => \N__20362\
        );

    \I__4518\ : CascadeBuf
    port map (
            O => \N__20365\,
            I => \N__20359\
        );

    \I__4517\ : CascadeMux
    port map (
            O => \N__20362\,
            I => \N__20356\
        );

    \I__4516\ : CascadeMux
    port map (
            O => \N__20359\,
            I => \N__20353\
        );

    \I__4515\ : CascadeBuf
    port map (
            O => \N__20356\,
            I => \N__20350\
        );

    \I__4514\ : CascadeBuf
    port map (
            O => \N__20353\,
            I => \N__20347\
        );

    \I__4513\ : CascadeMux
    port map (
            O => \N__20350\,
            I => \N__20344\
        );

    \I__4512\ : CascadeMux
    port map (
            O => \N__20347\,
            I => \N__20341\
        );

    \I__4511\ : InMux
    port map (
            O => \N__20344\,
            I => \N__20338\
        );

    \I__4510\ : InMux
    port map (
            O => \N__20341\,
            I => \N__20335\
        );

    \I__4509\ : LocalMux
    port map (
            O => \N__20338\,
            I => \N__20332\
        );

    \I__4508\ : LocalMux
    port map (
            O => \N__20335\,
            I => \N__20329\
        );

    \I__4507\ : Span4Mux_h
    port map (
            O => \N__20332\,
            I => \N__20326\
        );

    \I__4506\ : Span4Mux_v
    port map (
            O => \N__20329\,
            I => \N__20323\
        );

    \I__4505\ : Span4Mux_h
    port map (
            O => \N__20326\,
            I => \N__20320\
        );

    \I__4504\ : Sp12to4
    port map (
            O => \N__20323\,
            I => \N__20317\
        );

    \I__4503\ : Sp12to4
    port map (
            O => \N__20320\,
            I => \N__20314\
        );

    \I__4502\ : Span12Mux_h
    port map (
            O => \N__20317\,
            I => \N__20309\
        );

    \I__4501\ : Span12Mux_s5_v
    port map (
            O => \N__20314\,
            I => \N__20309\
        );

    \I__4500\ : Odrv12
    port map (
            O => \N__20309\,
            I => n26
        );

    \I__4499\ : InMux
    port map (
            O => \N__20306\,
            I => \N__20303\
        );

    \I__4498\ : LocalMux
    port map (
            O => \N__20303\,
            I => \N__20300\
        );

    \I__4497\ : Span4Mux_v
    port map (
            O => \N__20300\,
            I => \N__20297\
        );

    \I__4496\ : Span4Mux_h
    port map (
            O => \N__20297\,
            I => \N__20294\
        );

    \I__4495\ : Sp12to4
    port map (
            O => \N__20294\,
            I => \N__20291\
        );

    \I__4494\ : Span12Mux_v
    port map (
            O => \N__20291\,
            I => \N__20288\
        );

    \I__4493\ : Odrv12
    port map (
            O => \N__20288\,
            I => \line_buffer.n535\
        );

    \I__4492\ : CascadeMux
    port map (
            O => \N__20285\,
            I => \N__20282\
        );

    \I__4491\ : InMux
    port map (
            O => \N__20282\,
            I => \N__20279\
        );

    \I__4490\ : LocalMux
    port map (
            O => \N__20279\,
            I => \N__20276\
        );

    \I__4489\ : Span4Mux_h
    port map (
            O => \N__20276\,
            I => \N__20273\
        );

    \I__4488\ : Sp12to4
    port map (
            O => \N__20273\,
            I => \N__20270\
        );

    \I__4487\ : Span12Mux_v
    port map (
            O => \N__20270\,
            I => \N__20267\
        );

    \I__4486\ : Odrv12
    port map (
            O => \N__20267\,
            I => \line_buffer.n527\
        );

    \I__4485\ : InMux
    port map (
            O => \N__20264\,
            I => \N__20248\
        );

    \I__4484\ : InMux
    port map (
            O => \N__20263\,
            I => \N__20243\
        );

    \I__4483\ : InMux
    port map (
            O => \N__20262\,
            I => \N__20243\
        );

    \I__4482\ : InMux
    port map (
            O => \N__20261\,
            I => \N__20240\
        );

    \I__4481\ : CascadeMux
    port map (
            O => \N__20260\,
            I => \N__20237\
        );

    \I__4480\ : InMux
    port map (
            O => \N__20259\,
            I => \N__20233\
        );

    \I__4479\ : InMux
    port map (
            O => \N__20258\,
            I => \N__20230\
        );

    \I__4478\ : InMux
    port map (
            O => \N__20257\,
            I => \N__20227\
        );

    \I__4477\ : InMux
    port map (
            O => \N__20256\,
            I => \N__20223\
        );

    \I__4476\ : InMux
    port map (
            O => \N__20255\,
            I => \N__20220\
        );

    \I__4475\ : InMux
    port map (
            O => \N__20254\,
            I => \N__20217\
        );

    \I__4474\ : InMux
    port map (
            O => \N__20253\,
            I => \N__20214\
        );

    \I__4473\ : InMux
    port map (
            O => \N__20252\,
            I => \N__20209\
        );

    \I__4472\ : InMux
    port map (
            O => \N__20251\,
            I => \N__20209\
        );

    \I__4471\ : LocalMux
    port map (
            O => \N__20248\,
            I => \N__20206\
        );

    \I__4470\ : LocalMux
    port map (
            O => \N__20243\,
            I => \N__20201\
        );

    \I__4469\ : LocalMux
    port map (
            O => \N__20240\,
            I => \N__20201\
        );

    \I__4468\ : InMux
    port map (
            O => \N__20237\,
            I => \N__20196\
        );

    \I__4467\ : InMux
    port map (
            O => \N__20236\,
            I => \N__20196\
        );

    \I__4466\ : LocalMux
    port map (
            O => \N__20233\,
            I => \N__20190\
        );

    \I__4465\ : LocalMux
    port map (
            O => \N__20230\,
            I => \N__20185\
        );

    \I__4464\ : LocalMux
    port map (
            O => \N__20227\,
            I => \N__20185\
        );

    \I__4463\ : InMux
    port map (
            O => \N__20226\,
            I => \N__20182\
        );

    \I__4462\ : LocalMux
    port map (
            O => \N__20223\,
            I => \N__20172\
        );

    \I__4461\ : LocalMux
    port map (
            O => \N__20220\,
            I => \N__20172\
        );

    \I__4460\ : LocalMux
    port map (
            O => \N__20217\,
            I => \N__20172\
        );

    \I__4459\ : LocalMux
    port map (
            O => \N__20214\,
            I => \N__20167\
        );

    \I__4458\ : LocalMux
    port map (
            O => \N__20209\,
            I => \N__20167\
        );

    \I__4457\ : Span4Mux_h
    port map (
            O => \N__20206\,
            I => \N__20164\
        );

    \I__4456\ : Span4Mux_v
    port map (
            O => \N__20201\,
            I => \N__20156\
        );

    \I__4455\ : LocalMux
    port map (
            O => \N__20196\,
            I => \N__20156\
        );

    \I__4454\ : InMux
    port map (
            O => \N__20195\,
            I => \N__20153\
        );

    \I__4453\ : InMux
    port map (
            O => \N__20194\,
            I => \N__20150\
        );

    \I__4452\ : InMux
    port map (
            O => \N__20193\,
            I => \N__20147\
        );

    \I__4451\ : Span4Mux_v
    port map (
            O => \N__20190\,
            I => \N__20144\
        );

    \I__4450\ : Span4Mux_v
    port map (
            O => \N__20185\,
            I => \N__20141\
        );

    \I__4449\ : LocalMux
    port map (
            O => \N__20182\,
            I => \N__20138\
        );

    \I__4448\ : InMux
    port map (
            O => \N__20181\,
            I => \N__20135\
        );

    \I__4447\ : InMux
    port map (
            O => \N__20180\,
            I => \N__20130\
        );

    \I__4446\ : InMux
    port map (
            O => \N__20179\,
            I => \N__20130\
        );

    \I__4445\ : Span4Mux_v
    port map (
            O => \N__20172\,
            I => \N__20122\
        );

    \I__4444\ : Span4Mux_v
    port map (
            O => \N__20167\,
            I => \N__20122\
        );

    \I__4443\ : Span4Mux_v
    port map (
            O => \N__20164\,
            I => \N__20119\
        );

    \I__4442\ : InMux
    port map (
            O => \N__20163\,
            I => \N__20112\
        );

    \I__4441\ : InMux
    port map (
            O => \N__20162\,
            I => \N__20112\
        );

    \I__4440\ : InMux
    port map (
            O => \N__20161\,
            I => \N__20112\
        );

    \I__4439\ : Span4Mux_v
    port map (
            O => \N__20156\,
            I => \N__20109\
        );

    \I__4438\ : LocalMux
    port map (
            O => \N__20153\,
            I => \N__20104\
        );

    \I__4437\ : LocalMux
    port map (
            O => \N__20150\,
            I => \N__20104\
        );

    \I__4436\ : LocalMux
    port map (
            O => \N__20147\,
            I => \N__20091\
        );

    \I__4435\ : Span4Mux_h
    port map (
            O => \N__20144\,
            I => \N__20091\
        );

    \I__4434\ : Span4Mux_h
    port map (
            O => \N__20141\,
            I => \N__20091\
        );

    \I__4433\ : Span4Mux_v
    port map (
            O => \N__20138\,
            I => \N__20091\
        );

    \I__4432\ : LocalMux
    port map (
            O => \N__20135\,
            I => \N__20091\
        );

    \I__4431\ : LocalMux
    port map (
            O => \N__20130\,
            I => \N__20091\
        );

    \I__4430\ : InMux
    port map (
            O => \N__20129\,
            I => \N__20084\
        );

    \I__4429\ : InMux
    port map (
            O => \N__20128\,
            I => \N__20084\
        );

    \I__4428\ : InMux
    port map (
            O => \N__20127\,
            I => \N__20084\
        );

    \I__4427\ : Odrv4
    port map (
            O => \N__20122\,
            I => \transmit_module.n3678\
        );

    \I__4426\ : Odrv4
    port map (
            O => \N__20119\,
            I => \transmit_module.n3678\
        );

    \I__4425\ : LocalMux
    port map (
            O => \N__20112\,
            I => \transmit_module.n3678\
        );

    \I__4424\ : Odrv4
    port map (
            O => \N__20109\,
            I => \transmit_module.n3678\
        );

    \I__4423\ : Odrv12
    port map (
            O => \N__20104\,
            I => \transmit_module.n3678\
        );

    \I__4422\ : Odrv4
    port map (
            O => \N__20091\,
            I => \transmit_module.n3678\
        );

    \I__4421\ : LocalMux
    port map (
            O => \N__20084\,
            I => \transmit_module.n3678\
        );

    \I__4420\ : SRMux
    port map (
            O => \N__20069\,
            I => \N__20062\
        );

    \I__4419\ : SRMux
    port map (
            O => \N__20068\,
            I => \N__20051\
        );

    \I__4418\ : SRMux
    port map (
            O => \N__20067\,
            I => \N__20046\
        );

    \I__4417\ : CascadeMux
    port map (
            O => \N__20066\,
            I => \N__20038\
        );

    \I__4416\ : SRMux
    port map (
            O => \N__20065\,
            I => \N__20029\
        );

    \I__4415\ : LocalMux
    port map (
            O => \N__20062\,
            I => \N__20026\
        );

    \I__4414\ : SRMux
    port map (
            O => \N__20061\,
            I => \N__20023\
        );

    \I__4413\ : SRMux
    port map (
            O => \N__20060\,
            I => \N__20020\
        );

    \I__4412\ : CascadeMux
    port map (
            O => \N__20059\,
            I => \N__20014\
        );

    \I__4411\ : SRMux
    port map (
            O => \N__20058\,
            I => \N__20008\
        );

    \I__4410\ : SRMux
    port map (
            O => \N__20057\,
            I => \N__20003\
        );

    \I__4409\ : SRMux
    port map (
            O => \N__20056\,
            I => \N__19998\
        );

    \I__4408\ : SRMux
    port map (
            O => \N__20055\,
            I => \N__19991\
        );

    \I__4407\ : SRMux
    port map (
            O => \N__20054\,
            I => \N__19988\
        );

    \I__4406\ : LocalMux
    port map (
            O => \N__20051\,
            I => \N__19985\
        );

    \I__4405\ : SRMux
    port map (
            O => \N__20050\,
            I => \N__19982\
        );

    \I__4404\ : SRMux
    port map (
            O => \N__20049\,
            I => \N__19978\
        );

    \I__4403\ : LocalMux
    port map (
            O => \N__20046\,
            I => \N__19975\
        );

    \I__4402\ : SRMux
    port map (
            O => \N__20045\,
            I => \N__19972\
        );

    \I__4401\ : SRMux
    port map (
            O => \N__20044\,
            I => \N__19968\
        );

    \I__4400\ : SRMux
    port map (
            O => \N__20043\,
            I => \N__19965\
        );

    \I__4399\ : SRMux
    port map (
            O => \N__20042\,
            I => \N__19960\
        );

    \I__4398\ : SRMux
    port map (
            O => \N__20041\,
            I => \N__19957\
        );

    \I__4397\ : InMux
    port map (
            O => \N__20038\,
            I => \N__19952\
        );

    \I__4396\ : InMux
    port map (
            O => \N__20037\,
            I => \N__19952\
        );

    \I__4395\ : SRMux
    port map (
            O => \N__20036\,
            I => \N__19948\
        );

    \I__4394\ : CascadeMux
    port map (
            O => \N__20035\,
            I => \N__19945\
        );

    \I__4393\ : CascadeMux
    port map (
            O => \N__20034\,
            I => \N__19942\
        );

    \I__4392\ : CascadeMux
    port map (
            O => \N__20033\,
            I => \N__19939\
        );

    \I__4391\ : SRMux
    port map (
            O => \N__20032\,
            I => \N__19936\
        );

    \I__4390\ : LocalMux
    port map (
            O => \N__20029\,
            I => \N__19932\
        );

    \I__4389\ : Span4Mux_v
    port map (
            O => \N__20026\,
            I => \N__19925\
        );

    \I__4388\ : LocalMux
    port map (
            O => \N__20023\,
            I => \N__19925\
        );

    \I__4387\ : LocalMux
    port map (
            O => \N__20020\,
            I => \N__19925\
        );

    \I__4386\ : SRMux
    port map (
            O => \N__20019\,
            I => \N__19922\
        );

    \I__4385\ : SRMux
    port map (
            O => \N__20018\,
            I => \N__19919\
        );

    \I__4384\ : SRMux
    port map (
            O => \N__20017\,
            I => \N__19916\
        );

    \I__4383\ : InMux
    port map (
            O => \N__20014\,
            I => \N__19913\
        );

    \I__4382\ : CascadeMux
    port map (
            O => \N__20013\,
            I => \N__19907\
        );

    \I__4381\ : SRMux
    port map (
            O => \N__20012\,
            I => \N__19904\
        );

    \I__4380\ : SRMux
    port map (
            O => \N__20011\,
            I => \N__19901\
        );

    \I__4379\ : LocalMux
    port map (
            O => \N__20008\,
            I => \N__19898\
        );

    \I__4378\ : SRMux
    port map (
            O => \N__20007\,
            I => \N__19895\
        );

    \I__4377\ : SRMux
    port map (
            O => \N__20006\,
            I => \N__19892\
        );

    \I__4376\ : LocalMux
    port map (
            O => \N__20003\,
            I => \N__19889\
        );

    \I__4375\ : SRMux
    port map (
            O => \N__20002\,
            I => \N__19886\
        );

    \I__4374\ : SRMux
    port map (
            O => \N__20001\,
            I => \N__19883\
        );

    \I__4373\ : LocalMux
    port map (
            O => \N__19998\,
            I => \N__19880\
        );

    \I__4372\ : SRMux
    port map (
            O => \N__19997\,
            I => \N__19877\
        );

    \I__4371\ : IoInMux
    port map (
            O => \N__19996\,
            I => \N__19870\
        );

    \I__4370\ : CascadeMux
    port map (
            O => \N__19995\,
            I => \N__19867\
        );

    \I__4369\ : SRMux
    port map (
            O => \N__19994\,
            I => \N__19863\
        );

    \I__4368\ : LocalMux
    port map (
            O => \N__19991\,
            I => \N__19860\
        );

    \I__4367\ : LocalMux
    port map (
            O => \N__19988\,
            I => \N__19857\
        );

    \I__4366\ : Span4Mux_v
    port map (
            O => \N__19985\,
            I => \N__19852\
        );

    \I__4365\ : LocalMux
    port map (
            O => \N__19982\,
            I => \N__19852\
        );

    \I__4364\ : SRMux
    port map (
            O => \N__19981\,
            I => \N__19849\
        );

    \I__4363\ : LocalMux
    port map (
            O => \N__19978\,
            I => \N__19842\
        );

    \I__4362\ : Span4Mux_v
    port map (
            O => \N__19975\,
            I => \N__19842\
        );

    \I__4361\ : LocalMux
    port map (
            O => \N__19972\,
            I => \N__19842\
        );

    \I__4360\ : SRMux
    port map (
            O => \N__19971\,
            I => \N__19839\
        );

    \I__4359\ : LocalMux
    port map (
            O => \N__19968\,
            I => \N__19831\
        );

    \I__4358\ : LocalMux
    port map (
            O => \N__19965\,
            I => \N__19831\
        );

    \I__4357\ : SRMux
    port map (
            O => \N__19964\,
            I => \N__19828\
        );

    \I__4356\ : SRMux
    port map (
            O => \N__19963\,
            I => \N__19825\
        );

    \I__4355\ : LocalMux
    port map (
            O => \N__19960\,
            I => \N__19818\
        );

    \I__4354\ : LocalMux
    port map (
            O => \N__19957\,
            I => \N__19818\
        );

    \I__4353\ : LocalMux
    port map (
            O => \N__19952\,
            I => \N__19818\
        );

    \I__4352\ : CascadeMux
    port map (
            O => \N__19951\,
            I => \N__19815\
        );

    \I__4351\ : LocalMux
    port map (
            O => \N__19948\,
            I => \N__19812\
        );

    \I__4350\ : InMux
    port map (
            O => \N__19945\,
            I => \N__19807\
        );

    \I__4349\ : InMux
    port map (
            O => \N__19942\,
            I => \N__19807\
        );

    \I__4348\ : InMux
    port map (
            O => \N__19939\,
            I => \N__19804\
        );

    \I__4347\ : LocalMux
    port map (
            O => \N__19936\,
            I => \N__19801\
        );

    \I__4346\ : SRMux
    port map (
            O => \N__19935\,
            I => \N__19798\
        );

    \I__4345\ : Span4Mux_h
    port map (
            O => \N__19932\,
            I => \N__19791\
        );

    \I__4344\ : Span4Mux_h
    port map (
            O => \N__19925\,
            I => \N__19791\
        );

    \I__4343\ : LocalMux
    port map (
            O => \N__19922\,
            I => \N__19791\
        );

    \I__4342\ : LocalMux
    port map (
            O => \N__19919\,
            I => \N__19786\
        );

    \I__4341\ : LocalMux
    port map (
            O => \N__19916\,
            I => \N__19786\
        );

    \I__4340\ : LocalMux
    port map (
            O => \N__19913\,
            I => \N__19783\
        );

    \I__4339\ : SRMux
    port map (
            O => \N__19912\,
            I => \N__19780\
        );

    \I__4338\ : SRMux
    port map (
            O => \N__19911\,
            I => \N__19777\
        );

    \I__4337\ : InMux
    port map (
            O => \N__19910\,
            I => \N__19772\
        );

    \I__4336\ : InMux
    port map (
            O => \N__19907\,
            I => \N__19772\
        );

    \I__4335\ : LocalMux
    port map (
            O => \N__19904\,
            I => \N__19769\
        );

    \I__4334\ : LocalMux
    port map (
            O => \N__19901\,
            I => \N__19766\
        );

    \I__4333\ : Span4Mux_v
    port map (
            O => \N__19898\,
            I => \N__19763\
        );

    \I__4332\ : LocalMux
    port map (
            O => \N__19895\,
            I => \N__19758\
        );

    \I__4331\ : LocalMux
    port map (
            O => \N__19892\,
            I => \N__19758\
        );

    \I__4330\ : Span4Mux_h
    port map (
            O => \N__19889\,
            I => \N__19751\
        );

    \I__4329\ : LocalMux
    port map (
            O => \N__19886\,
            I => \N__19751\
        );

    \I__4328\ : LocalMux
    port map (
            O => \N__19883\,
            I => \N__19751\
        );

    \I__4327\ : Span4Mux_h
    port map (
            O => \N__19880\,
            I => \N__19746\
        );

    \I__4326\ : LocalMux
    port map (
            O => \N__19877\,
            I => \N__19746\
        );

    \I__4325\ : SRMux
    port map (
            O => \N__19876\,
            I => \N__19743\
        );

    \I__4324\ : CascadeMux
    port map (
            O => \N__19875\,
            I => \N__19740\
        );

    \I__4323\ : InMux
    port map (
            O => \N__19874\,
            I => \N__19734\
        );

    \I__4322\ : InMux
    port map (
            O => \N__19873\,
            I => \N__19734\
        );

    \I__4321\ : LocalMux
    port map (
            O => \N__19870\,
            I => \N__19731\
        );

    \I__4320\ : InMux
    port map (
            O => \N__19867\,
            I => \N__19728\
        );

    \I__4319\ : CascadeMux
    port map (
            O => \N__19866\,
            I => \N__19724\
        );

    \I__4318\ : LocalMux
    port map (
            O => \N__19863\,
            I => \N__19718\
        );

    \I__4317\ : Span4Mux_v
    port map (
            O => \N__19860\,
            I => \N__19709\
        );

    \I__4316\ : Span4Mux_h
    port map (
            O => \N__19857\,
            I => \N__19709\
        );

    \I__4315\ : Span4Mux_v
    port map (
            O => \N__19852\,
            I => \N__19709\
        );

    \I__4314\ : LocalMux
    port map (
            O => \N__19849\,
            I => \N__19709\
        );

    \I__4313\ : Span4Mux_v
    port map (
            O => \N__19842\,
            I => \N__19704\
        );

    \I__4312\ : LocalMux
    port map (
            O => \N__19839\,
            I => \N__19704\
        );

    \I__4311\ : CascadeMux
    port map (
            O => \N__19838\,
            I => \N__19701\
        );

    \I__4310\ : CascadeMux
    port map (
            O => \N__19837\,
            I => \N__19698\
        );

    \I__4309\ : CascadeMux
    port map (
            O => \N__19836\,
            I => \N__19695\
        );

    \I__4308\ : Span4Mux_h
    port map (
            O => \N__19831\,
            I => \N__19685\
        );

    \I__4307\ : LocalMux
    port map (
            O => \N__19828\,
            I => \N__19685\
        );

    \I__4306\ : LocalMux
    port map (
            O => \N__19825\,
            I => \N__19685\
        );

    \I__4305\ : Span4Mux_v
    port map (
            O => \N__19818\,
            I => \N__19682\
        );

    \I__4304\ : InMux
    port map (
            O => \N__19815\,
            I => \N__19679\
        );

    \I__4303\ : Span4Mux_v
    port map (
            O => \N__19812\,
            I => \N__19674\
        );

    \I__4302\ : LocalMux
    port map (
            O => \N__19807\,
            I => \N__19674\
        );

    \I__4301\ : LocalMux
    port map (
            O => \N__19804\,
            I => \N__19671\
        );

    \I__4300\ : Span4Mux_v
    port map (
            O => \N__19801\,
            I => \N__19660\
        );

    \I__4299\ : LocalMux
    port map (
            O => \N__19798\,
            I => \N__19660\
        );

    \I__4298\ : Span4Mux_h
    port map (
            O => \N__19791\,
            I => \N__19660\
        );

    \I__4297\ : Span4Mux_v
    port map (
            O => \N__19786\,
            I => \N__19660\
        );

    \I__4296\ : Span4Mux_h
    port map (
            O => \N__19783\,
            I => \N__19660\
        );

    \I__4295\ : LocalMux
    port map (
            O => \N__19780\,
            I => \N__19653\
        );

    \I__4294\ : LocalMux
    port map (
            O => \N__19777\,
            I => \N__19653\
        );

    \I__4293\ : LocalMux
    port map (
            O => \N__19772\,
            I => \N__19653\
        );

    \I__4292\ : Span4Mux_h
    port map (
            O => \N__19769\,
            I => \N__19638\
        );

    \I__4291\ : Span4Mux_v
    port map (
            O => \N__19766\,
            I => \N__19638\
        );

    \I__4290\ : Span4Mux_v
    port map (
            O => \N__19763\,
            I => \N__19638\
        );

    \I__4289\ : Span4Mux_h
    port map (
            O => \N__19758\,
            I => \N__19638\
        );

    \I__4288\ : Span4Mux_v
    port map (
            O => \N__19751\,
            I => \N__19638\
        );

    \I__4287\ : Span4Mux_v
    port map (
            O => \N__19746\,
            I => \N__19638\
        );

    \I__4286\ : LocalMux
    port map (
            O => \N__19743\,
            I => \N__19638\
        );

    \I__4285\ : InMux
    port map (
            O => \N__19740\,
            I => \N__19633\
        );

    \I__4284\ : InMux
    port map (
            O => \N__19739\,
            I => \N__19633\
        );

    \I__4283\ : LocalMux
    port map (
            O => \N__19734\,
            I => \N__19630\
        );

    \I__4282\ : Span12Mux_s0_h
    port map (
            O => \N__19731\,
            I => \N__19627\
        );

    \I__4281\ : LocalMux
    port map (
            O => \N__19728\,
            I => \N__19624\
        );

    \I__4280\ : InMux
    port map (
            O => \N__19727\,
            I => \N__19621\
        );

    \I__4279\ : InMux
    port map (
            O => \N__19724\,
            I => \N__19616\
        );

    \I__4278\ : InMux
    port map (
            O => \N__19723\,
            I => \N__19616\
        );

    \I__4277\ : CascadeMux
    port map (
            O => \N__19722\,
            I => \N__19613\
        );

    \I__4276\ : CascadeMux
    port map (
            O => \N__19721\,
            I => \N__19609\
        );

    \I__4275\ : Span4Mux_v
    port map (
            O => \N__19718\,
            I => \N__19604\
        );

    \I__4274\ : Span4Mux_v
    port map (
            O => \N__19709\,
            I => \N__19599\
        );

    \I__4273\ : Span4Mux_h
    port map (
            O => \N__19704\,
            I => \N__19599\
        );

    \I__4272\ : InMux
    port map (
            O => \N__19701\,
            I => \N__19596\
        );

    \I__4271\ : InMux
    port map (
            O => \N__19698\,
            I => \N__19593\
        );

    \I__4270\ : InMux
    port map (
            O => \N__19695\,
            I => \N__19586\
        );

    \I__4269\ : InMux
    port map (
            O => \N__19694\,
            I => \N__19586\
        );

    \I__4268\ : InMux
    port map (
            O => \N__19693\,
            I => \N__19586\
        );

    \I__4267\ : InMux
    port map (
            O => \N__19692\,
            I => \N__19583\
        );

    \I__4266\ : Span4Mux_v
    port map (
            O => \N__19685\,
            I => \N__19568\
        );

    \I__4265\ : Span4Mux_h
    port map (
            O => \N__19682\,
            I => \N__19568\
        );

    \I__4264\ : LocalMux
    port map (
            O => \N__19679\,
            I => \N__19568\
        );

    \I__4263\ : Span4Mux_h
    port map (
            O => \N__19674\,
            I => \N__19568\
        );

    \I__4262\ : Span4Mux_v
    port map (
            O => \N__19671\,
            I => \N__19568\
        );

    \I__4261\ : Span4Mux_v
    port map (
            O => \N__19660\,
            I => \N__19568\
        );

    \I__4260\ : Span4Mux_v
    port map (
            O => \N__19653\,
            I => \N__19568\
        );

    \I__4259\ : Span4Mux_h
    port map (
            O => \N__19638\,
            I => \N__19561\
        );

    \I__4258\ : LocalMux
    port map (
            O => \N__19633\,
            I => \N__19561\
        );

    \I__4257\ : Span4Mux_v
    port map (
            O => \N__19630\,
            I => \N__19561\
        );

    \I__4256\ : Span12Mux_h
    port map (
            O => \N__19627\,
            I => \N__19552\
        );

    \I__4255\ : Sp12to4
    port map (
            O => \N__19624\,
            I => \N__19552\
        );

    \I__4254\ : LocalMux
    port map (
            O => \N__19621\,
            I => \N__19552\
        );

    \I__4253\ : LocalMux
    port map (
            O => \N__19616\,
            I => \N__19552\
        );

    \I__4252\ : InMux
    port map (
            O => \N__19613\,
            I => \N__19547\
        );

    \I__4251\ : InMux
    port map (
            O => \N__19612\,
            I => \N__19547\
        );

    \I__4250\ : InMux
    port map (
            O => \N__19609\,
            I => \N__19540\
        );

    \I__4249\ : InMux
    port map (
            O => \N__19608\,
            I => \N__19540\
        );

    \I__4248\ : InMux
    port map (
            O => \N__19607\,
            I => \N__19540\
        );

    \I__4247\ : Odrv4
    port map (
            O => \N__19604\,
            I => \ADV_VSYNC_c\
        );

    \I__4246\ : Odrv4
    port map (
            O => \N__19599\,
            I => \ADV_VSYNC_c\
        );

    \I__4245\ : LocalMux
    port map (
            O => \N__19596\,
            I => \ADV_VSYNC_c\
        );

    \I__4244\ : LocalMux
    port map (
            O => \N__19593\,
            I => \ADV_VSYNC_c\
        );

    \I__4243\ : LocalMux
    port map (
            O => \N__19586\,
            I => \ADV_VSYNC_c\
        );

    \I__4242\ : LocalMux
    port map (
            O => \N__19583\,
            I => \ADV_VSYNC_c\
        );

    \I__4241\ : Odrv4
    port map (
            O => \N__19568\,
            I => \ADV_VSYNC_c\
        );

    \I__4240\ : Odrv4
    port map (
            O => \N__19561\,
            I => \ADV_VSYNC_c\
        );

    \I__4239\ : Odrv12
    port map (
            O => \N__19552\,
            I => \ADV_VSYNC_c\
        );

    \I__4238\ : LocalMux
    port map (
            O => \N__19547\,
            I => \ADV_VSYNC_c\
        );

    \I__4237\ : LocalMux
    port map (
            O => \N__19540\,
            I => \ADV_VSYNC_c\
        );

    \I__4236\ : InMux
    port map (
            O => \N__19517\,
            I => \N__19513\
        );

    \I__4235\ : CascadeMux
    port map (
            O => \N__19516\,
            I => \N__19510\
        );

    \I__4234\ : LocalMux
    port map (
            O => \N__19513\,
            I => \N__19507\
        );

    \I__4233\ : InMux
    port map (
            O => \N__19510\,
            I => \N__19504\
        );

    \I__4232\ : Odrv12
    port map (
            O => \N__19507\,
            I => \transmit_module.n113\
        );

    \I__4231\ : LocalMux
    port map (
            O => \N__19504\,
            I => \transmit_module.n113\
        );

    \I__4230\ : InMux
    port map (
            O => \N__19499\,
            I => \N__19496\
        );

    \I__4229\ : LocalMux
    port map (
            O => \N__19496\,
            I => \N__19492\
        );

    \I__4228\ : InMux
    port map (
            O => \N__19495\,
            I => \N__19489\
        );

    \I__4227\ : Span4Mux_v
    port map (
            O => \N__19492\,
            I => \N__19486\
        );

    \I__4226\ : LocalMux
    port map (
            O => \N__19489\,
            I => \transmit_module.n144\
        );

    \I__4225\ : Odrv4
    port map (
            O => \N__19486\,
            I => \transmit_module.n144\
        );

    \I__4224\ : CascadeMux
    port map (
            O => \N__19481\,
            I => \N__19477\
        );

    \I__4223\ : CascadeMux
    port map (
            O => \N__19480\,
            I => \N__19474\
        );

    \I__4222\ : CascadeBuf
    port map (
            O => \N__19477\,
            I => \N__19471\
        );

    \I__4221\ : CascadeBuf
    port map (
            O => \N__19474\,
            I => \N__19468\
        );

    \I__4220\ : CascadeMux
    port map (
            O => \N__19471\,
            I => \N__19465\
        );

    \I__4219\ : CascadeMux
    port map (
            O => \N__19468\,
            I => \N__19462\
        );

    \I__4218\ : CascadeBuf
    port map (
            O => \N__19465\,
            I => \N__19459\
        );

    \I__4217\ : CascadeBuf
    port map (
            O => \N__19462\,
            I => \N__19456\
        );

    \I__4216\ : CascadeMux
    port map (
            O => \N__19459\,
            I => \N__19453\
        );

    \I__4215\ : CascadeMux
    port map (
            O => \N__19456\,
            I => \N__19450\
        );

    \I__4214\ : CascadeBuf
    port map (
            O => \N__19453\,
            I => \N__19447\
        );

    \I__4213\ : CascadeBuf
    port map (
            O => \N__19450\,
            I => \N__19444\
        );

    \I__4212\ : CascadeMux
    port map (
            O => \N__19447\,
            I => \N__19441\
        );

    \I__4211\ : CascadeMux
    port map (
            O => \N__19444\,
            I => \N__19438\
        );

    \I__4210\ : CascadeBuf
    port map (
            O => \N__19441\,
            I => \N__19435\
        );

    \I__4209\ : CascadeBuf
    port map (
            O => \N__19438\,
            I => \N__19432\
        );

    \I__4208\ : CascadeMux
    port map (
            O => \N__19435\,
            I => \N__19429\
        );

    \I__4207\ : CascadeMux
    port map (
            O => \N__19432\,
            I => \N__19426\
        );

    \I__4206\ : CascadeBuf
    port map (
            O => \N__19429\,
            I => \N__19423\
        );

    \I__4205\ : CascadeBuf
    port map (
            O => \N__19426\,
            I => \N__19420\
        );

    \I__4204\ : CascadeMux
    port map (
            O => \N__19423\,
            I => \N__19417\
        );

    \I__4203\ : CascadeMux
    port map (
            O => \N__19420\,
            I => \N__19414\
        );

    \I__4202\ : CascadeBuf
    port map (
            O => \N__19417\,
            I => \N__19411\
        );

    \I__4201\ : CascadeBuf
    port map (
            O => \N__19414\,
            I => \N__19408\
        );

    \I__4200\ : CascadeMux
    port map (
            O => \N__19411\,
            I => \N__19405\
        );

    \I__4199\ : CascadeMux
    port map (
            O => \N__19408\,
            I => \N__19402\
        );

    \I__4198\ : CascadeBuf
    port map (
            O => \N__19405\,
            I => \N__19399\
        );

    \I__4197\ : CascadeBuf
    port map (
            O => \N__19402\,
            I => \N__19396\
        );

    \I__4196\ : CascadeMux
    port map (
            O => \N__19399\,
            I => \N__19393\
        );

    \I__4195\ : CascadeMux
    port map (
            O => \N__19396\,
            I => \N__19390\
        );

    \I__4194\ : CascadeBuf
    port map (
            O => \N__19393\,
            I => \N__19387\
        );

    \I__4193\ : CascadeBuf
    port map (
            O => \N__19390\,
            I => \N__19384\
        );

    \I__4192\ : CascadeMux
    port map (
            O => \N__19387\,
            I => \N__19381\
        );

    \I__4191\ : CascadeMux
    port map (
            O => \N__19384\,
            I => \N__19378\
        );

    \I__4190\ : CascadeBuf
    port map (
            O => \N__19381\,
            I => \N__19375\
        );

    \I__4189\ : CascadeBuf
    port map (
            O => \N__19378\,
            I => \N__19372\
        );

    \I__4188\ : CascadeMux
    port map (
            O => \N__19375\,
            I => \N__19369\
        );

    \I__4187\ : CascadeMux
    port map (
            O => \N__19372\,
            I => \N__19366\
        );

    \I__4186\ : CascadeBuf
    port map (
            O => \N__19369\,
            I => \N__19363\
        );

    \I__4185\ : CascadeBuf
    port map (
            O => \N__19366\,
            I => \N__19360\
        );

    \I__4184\ : CascadeMux
    port map (
            O => \N__19363\,
            I => \N__19357\
        );

    \I__4183\ : CascadeMux
    port map (
            O => \N__19360\,
            I => \N__19354\
        );

    \I__4182\ : CascadeBuf
    port map (
            O => \N__19357\,
            I => \N__19351\
        );

    \I__4181\ : CascadeBuf
    port map (
            O => \N__19354\,
            I => \N__19348\
        );

    \I__4180\ : CascadeMux
    port map (
            O => \N__19351\,
            I => \N__19345\
        );

    \I__4179\ : CascadeMux
    port map (
            O => \N__19348\,
            I => \N__19342\
        );

    \I__4178\ : CascadeBuf
    port map (
            O => \N__19345\,
            I => \N__19339\
        );

    \I__4177\ : CascadeBuf
    port map (
            O => \N__19342\,
            I => \N__19336\
        );

    \I__4176\ : CascadeMux
    port map (
            O => \N__19339\,
            I => \N__19333\
        );

    \I__4175\ : CascadeMux
    port map (
            O => \N__19336\,
            I => \N__19330\
        );

    \I__4174\ : CascadeBuf
    port map (
            O => \N__19333\,
            I => \N__19327\
        );

    \I__4173\ : CascadeBuf
    port map (
            O => \N__19330\,
            I => \N__19324\
        );

    \I__4172\ : CascadeMux
    port map (
            O => \N__19327\,
            I => \N__19321\
        );

    \I__4171\ : CascadeMux
    port map (
            O => \N__19324\,
            I => \N__19318\
        );

    \I__4170\ : CascadeBuf
    port map (
            O => \N__19321\,
            I => \N__19315\
        );

    \I__4169\ : CascadeBuf
    port map (
            O => \N__19318\,
            I => \N__19312\
        );

    \I__4168\ : CascadeMux
    port map (
            O => \N__19315\,
            I => \N__19309\
        );

    \I__4167\ : CascadeMux
    port map (
            O => \N__19312\,
            I => \N__19306\
        );

    \I__4166\ : CascadeBuf
    port map (
            O => \N__19309\,
            I => \N__19303\
        );

    \I__4165\ : CascadeBuf
    port map (
            O => \N__19306\,
            I => \N__19300\
        );

    \I__4164\ : CascadeMux
    port map (
            O => \N__19303\,
            I => \N__19297\
        );

    \I__4163\ : CascadeMux
    port map (
            O => \N__19300\,
            I => \N__19294\
        );

    \I__4162\ : InMux
    port map (
            O => \N__19297\,
            I => \N__19291\
        );

    \I__4161\ : InMux
    port map (
            O => \N__19294\,
            I => \N__19288\
        );

    \I__4160\ : LocalMux
    port map (
            O => \N__19291\,
            I => \N__19285\
        );

    \I__4159\ : LocalMux
    port map (
            O => \N__19288\,
            I => \N__19282\
        );

    \I__4158\ : Span12Mux_s11_h
    port map (
            O => \N__19285\,
            I => \N__19279\
        );

    \I__4157\ : Sp12to4
    port map (
            O => \N__19282\,
            I => \N__19276\
        );

    \I__4156\ : Span12Mux_v
    port map (
            O => \N__19279\,
            I => \N__19271\
        );

    \I__4155\ : Span12Mux_v
    port map (
            O => \N__19276\,
            I => \N__19271\
        );

    \I__4154\ : Odrv12
    port map (
            O => \N__19271\,
            I => n25
        );

    \I__4153\ : IoInMux
    port map (
            O => \N__19268\,
            I => \N__19265\
        );

    \I__4152\ : LocalMux
    port map (
            O => \N__19265\,
            I => \N__19260\
        );

    \I__4151\ : IoInMux
    port map (
            O => \N__19264\,
            I => \N__19257\
        );

    \I__4150\ : IoInMux
    port map (
            O => \N__19263\,
            I => \N__19254\
        );

    \I__4149\ : IoSpan4Mux
    port map (
            O => \N__19260\,
            I => \N__19251\
        );

    \I__4148\ : LocalMux
    port map (
            O => \N__19257\,
            I => \N__19248\
        );

    \I__4147\ : LocalMux
    port map (
            O => \N__19254\,
            I => \N__19245\
        );

    \I__4146\ : Span4Mux_s2_v
    port map (
            O => \N__19251\,
            I => \N__19242\
        );

    \I__4145\ : IoSpan4Mux
    port map (
            O => \N__19248\,
            I => \N__19239\
        );

    \I__4144\ : Span4Mux_s3_h
    port map (
            O => \N__19245\,
            I => \N__19236\
        );

    \I__4143\ : Sp12to4
    port map (
            O => \N__19242\,
            I => \N__19233\
        );

    \I__4142\ : Span4Mux_s1_v
    port map (
            O => \N__19239\,
            I => \N__19230\
        );

    \I__4141\ : Span4Mux_h
    port map (
            O => \N__19236\,
            I => \N__19227\
        );

    \I__4140\ : Span12Mux_v
    port map (
            O => \N__19233\,
            I => \N__19224\
        );

    \I__4139\ : Sp12to4
    port map (
            O => \N__19230\,
            I => \N__19221\
        );

    \I__4138\ : Span4Mux_h
    port map (
            O => \N__19227\,
            I => \N__19218\
        );

    \I__4137\ : Span12Mux_h
    port map (
            O => \N__19224\,
            I => \N__19213\
        );

    \I__4136\ : Span12Mux_h
    port map (
            O => \N__19221\,
            I => \N__19213\
        );

    \I__4135\ : Span4Mux_h
    port map (
            O => \N__19218\,
            I => \N__19210\
        );

    \I__4134\ : Odrv12
    port map (
            O => \N__19213\,
            I => n1818
        );

    \I__4133\ : Odrv4
    port map (
            O => \N__19210\,
            I => n1818
        );

    \I__4132\ : InMux
    port map (
            O => \N__19205\,
            I => \N__19202\
        );

    \I__4131\ : LocalMux
    port map (
            O => \N__19202\,
            I => \N__19199\
        );

    \I__4130\ : Sp12to4
    port map (
            O => \N__19199\,
            I => \N__19196\
        );

    \I__4129\ : Odrv12
    port map (
            O => \N__19196\,
            I => \line_buffer.n470\
        );

    \I__4128\ : CascadeMux
    port map (
            O => \N__19193\,
            I => \N__19190\
        );

    \I__4127\ : InMux
    port map (
            O => \N__19190\,
            I => \N__19187\
        );

    \I__4126\ : LocalMux
    port map (
            O => \N__19187\,
            I => \N__19184\
        );

    \I__4125\ : Span4Mux_v
    port map (
            O => \N__19184\,
            I => \N__19181\
        );

    \I__4124\ : Sp12to4
    port map (
            O => \N__19181\,
            I => \N__19178\
        );

    \I__4123\ : Span12Mux_h
    port map (
            O => \N__19178\,
            I => \N__19175\
        );

    \I__4122\ : Odrv12
    port map (
            O => \N__19175\,
            I => \line_buffer.n462\
        );

    \I__4121\ : InMux
    port map (
            O => \N__19172\,
            I => \N__19169\
        );

    \I__4120\ : LocalMux
    port map (
            O => \N__19169\,
            I => \N__19166\
        );

    \I__4119\ : Odrv12
    port map (
            O => \N__19166\,
            I => \line_buffer.n3590\
        );

    \I__4118\ : SRMux
    port map (
            O => \N__19163\,
            I => \N__19160\
        );

    \I__4117\ : LocalMux
    port map (
            O => \N__19160\,
            I => \receive_module.rx_counter.n2550\
        );

    \I__4116\ : InMux
    port map (
            O => \N__19157\,
            I => \N__19154\
        );

    \I__4115\ : LocalMux
    port map (
            O => \N__19154\,
            I => \N__19151\
        );

    \I__4114\ : Odrv4
    port map (
            O => \N__19151\,
            I => \tvp_video_buffer.BUFFER_1_6\
        );

    \I__4113\ : InMux
    port map (
            O => \N__19148\,
            I => \N__19143\
        );

    \I__4112\ : InMux
    port map (
            O => \N__19147\,
            I => \N__19140\
        );

    \I__4111\ : InMux
    port map (
            O => \N__19146\,
            I => \N__19137\
        );

    \I__4110\ : LocalMux
    port map (
            O => \N__19143\,
            I => \N__19130\
        );

    \I__4109\ : LocalMux
    port map (
            O => \N__19140\,
            I => \N__19130\
        );

    \I__4108\ : LocalMux
    port map (
            O => \N__19137\,
            I => \N__19127\
        );

    \I__4107\ : InMux
    port map (
            O => \N__19136\,
            I => \N__19124\
        );

    \I__4106\ : InMux
    port map (
            O => \N__19135\,
            I => \N__19121\
        );

    \I__4105\ : Span4Mux_v
    port map (
            O => \N__19130\,
            I => \N__19112\
        );

    \I__4104\ : Span4Mux_h
    port map (
            O => \N__19127\,
            I => \N__19112\
        );

    \I__4103\ : LocalMux
    port map (
            O => \N__19124\,
            I => \N__19112\
        );

    \I__4102\ : LocalMux
    port map (
            O => \N__19121\,
            I => \N__19108\
        );

    \I__4101\ : InMux
    port map (
            O => \N__19120\,
            I => \N__19105\
        );

    \I__4100\ : InMux
    port map (
            O => \N__19119\,
            I => \N__19102\
        );

    \I__4099\ : Span4Mux_v
    port map (
            O => \N__19112\,
            I => \N__19099\
        );

    \I__4098\ : InMux
    port map (
            O => \N__19111\,
            I => \N__19096\
        );

    \I__4097\ : Span4Mux_v
    port map (
            O => \N__19108\,
            I => \N__19093\
        );

    \I__4096\ : LocalMux
    port map (
            O => \N__19105\,
            I => \N__19090\
        );

    \I__4095\ : LocalMux
    port map (
            O => \N__19102\,
            I => \N__19087\
        );

    \I__4094\ : Span4Mux_v
    port map (
            O => \N__19099\,
            I => \N__19082\
        );

    \I__4093\ : LocalMux
    port map (
            O => \N__19096\,
            I => \N__19082\
        );

    \I__4092\ : Sp12to4
    port map (
            O => \N__19093\,
            I => \N__19078\
        );

    \I__4091\ : Span4Mux_s2_v
    port map (
            O => \N__19090\,
            I => \N__19073\
        );

    \I__4090\ : Span4Mux_v
    port map (
            O => \N__19087\,
            I => \N__19073\
        );

    \I__4089\ : Span4Mux_v
    port map (
            O => \N__19082\,
            I => \N__19070\
        );

    \I__4088\ : InMux
    port map (
            O => \N__19081\,
            I => \N__19067\
        );

    \I__4087\ : Span12Mux_h
    port map (
            O => \N__19078\,
            I => \N__19064\
        );

    \I__4086\ : Sp12to4
    port map (
            O => \N__19073\,
            I => \N__19061\
        );

    \I__4085\ : Span4Mux_h
    port map (
            O => \N__19070\,
            I => \N__19056\
        );

    \I__4084\ : LocalMux
    port map (
            O => \N__19067\,
            I => \N__19056\
        );

    \I__4083\ : Span12Mux_v
    port map (
            O => \N__19064\,
            I => \N__19051\
        );

    \I__4082\ : Span12Mux_h
    port map (
            O => \N__19061\,
            I => \N__19051\
        );

    \I__4081\ : Span4Mux_h
    port map (
            O => \N__19056\,
            I => \N__19048\
        );

    \I__4080\ : Odrv12
    port map (
            O => \N__19051\,
            I => \RX_DATA_6\
        );

    \I__4079\ : Odrv4
    port map (
            O => \N__19048\,
            I => \RX_DATA_6\
        );

    \I__4078\ : InMux
    port map (
            O => \N__19043\,
            I => \N__19040\
        );

    \I__4077\ : LocalMux
    port map (
            O => \N__19040\,
            I => \N__19037\
        );

    \I__4076\ : Span4Mux_v
    port map (
            O => \N__19037\,
            I => \N__19031\
        );

    \I__4075\ : InMux
    port map (
            O => \N__19036\,
            I => \N__19028\
        );

    \I__4074\ : InMux
    port map (
            O => \N__19035\,
            I => \N__19025\
        );

    \I__4073\ : InMux
    port map (
            O => \N__19034\,
            I => \N__19022\
        );

    \I__4072\ : Span4Mux_v
    port map (
            O => \N__19031\,
            I => \N__19016\
        );

    \I__4071\ : LocalMux
    port map (
            O => \N__19028\,
            I => \N__19016\
        );

    \I__4070\ : LocalMux
    port map (
            O => \N__19025\,
            I => \N__19013\
        );

    \I__4069\ : LocalMux
    port map (
            O => \N__19022\,
            I => \N__19010\
        );

    \I__4068\ : InMux
    port map (
            O => \N__19021\,
            I => \N__19007\
        );

    \I__4067\ : Span4Mux_v
    port map (
            O => \N__19016\,
            I => \N__19003\
        );

    \I__4066\ : Sp12to4
    port map (
            O => \N__19013\,
            I => \N__18998\
        );

    \I__4065\ : Span4Mux_h
    port map (
            O => \N__19010\,
            I => \N__18995\
        );

    \I__4064\ : LocalMux
    port map (
            O => \N__19007\,
            I => \N__18992\
        );

    \I__4063\ : InMux
    port map (
            O => \N__19006\,
            I => \N__18989\
        );

    \I__4062\ : Span4Mux_v
    port map (
            O => \N__19003\,
            I => \N__18986\
        );

    \I__4061\ : InMux
    port map (
            O => \N__19002\,
            I => \N__18983\
        );

    \I__4060\ : InMux
    port map (
            O => \N__19001\,
            I => \N__18980\
        );

    \I__4059\ : Span12Mux_s9_v
    port map (
            O => \N__18998\,
            I => \N__18977\
        );

    \I__4058\ : Span4Mux_h
    port map (
            O => \N__18995\,
            I => \N__18974\
        );

    \I__4057\ : Span4Mux_h
    port map (
            O => \N__18992\,
            I => \N__18971\
        );

    \I__4056\ : LocalMux
    port map (
            O => \N__18989\,
            I => \N__18968\
        );

    \I__4055\ : Sp12to4
    port map (
            O => \N__18986\,
            I => \N__18963\
        );

    \I__4054\ : LocalMux
    port map (
            O => \N__18983\,
            I => \N__18963\
        );

    \I__4053\ : LocalMux
    port map (
            O => \N__18980\,
            I => \N__18960\
        );

    \I__4052\ : Span12Mux_v
    port map (
            O => \N__18977\,
            I => \N__18956\
        );

    \I__4051\ : Span4Mux_h
    port map (
            O => \N__18974\,
            I => \N__18951\
        );

    \I__4050\ : Span4Mux_h
    port map (
            O => \N__18971\,
            I => \N__18951\
        );

    \I__4049\ : Span12Mux_h
    port map (
            O => \N__18968\,
            I => \N__18944\
        );

    \I__4048\ : Span12Mux_h
    port map (
            O => \N__18963\,
            I => \N__18944\
        );

    \I__4047\ : Span12Mux_h
    port map (
            O => \N__18960\,
            I => \N__18944\
        );

    \I__4046\ : InMux
    port map (
            O => \N__18959\,
            I => \N__18941\
        );

    \I__4045\ : Odrv12
    port map (
            O => \N__18956\,
            I => \RX_DATA_4\
        );

    \I__4044\ : Odrv4
    port map (
            O => \N__18951\,
            I => \RX_DATA_4\
        );

    \I__4043\ : Odrv12
    port map (
            O => \N__18944\,
            I => \RX_DATA_4\
        );

    \I__4042\ : LocalMux
    port map (
            O => \N__18941\,
            I => \RX_DATA_4\
        );

    \I__4041\ : CascadeMux
    port map (
            O => \N__18932\,
            I => \receive_module.sync_wd.n6_cascade_\
        );

    \I__4040\ : CascadeMux
    port map (
            O => \N__18929\,
            I => \receive_module.sync_wd.n4_cascade_\
        );

    \I__4039\ : InMux
    port map (
            O => \N__18926\,
            I => \N__18920\
        );

    \I__4038\ : InMux
    port map (
            O => \N__18925\,
            I => \N__18920\
        );

    \I__4037\ : LocalMux
    port map (
            O => \N__18920\,
            I => \N__18915\
        );

    \I__4036\ : InMux
    port map (
            O => \N__18919\,
            I => \N__18912\
        );

    \I__4035\ : InMux
    port map (
            O => \N__18918\,
            I => \N__18909\
        );

    \I__4034\ : Span4Mux_s2_v
    port map (
            O => \N__18915\,
            I => \N__18901\
        );

    \I__4033\ : LocalMux
    port map (
            O => \N__18912\,
            I => \N__18901\
        );

    \I__4032\ : LocalMux
    port map (
            O => \N__18909\,
            I => \N__18901\
        );

    \I__4031\ : InMux
    port map (
            O => \N__18908\,
            I => \N__18898\
        );

    \I__4030\ : Span4Mux_v
    port map (
            O => \N__18901\,
            I => \N__18887\
        );

    \I__4029\ : LocalMux
    port map (
            O => \N__18898\,
            I => \N__18887\
        );

    \I__4028\ : InMux
    port map (
            O => \N__18897\,
            I => \N__18880\
        );

    \I__4027\ : InMux
    port map (
            O => \N__18896\,
            I => \N__18880\
        );

    \I__4026\ : InMux
    port map (
            O => \N__18895\,
            I => \N__18880\
        );

    \I__4025\ : InMux
    port map (
            O => \N__18894\,
            I => \N__18873\
        );

    \I__4024\ : InMux
    port map (
            O => \N__18893\,
            I => \N__18873\
        );

    \I__4023\ : InMux
    port map (
            O => \N__18892\,
            I => \N__18873\
        );

    \I__4022\ : Span4Mux_v
    port map (
            O => \N__18887\,
            I => \N__18863\
        );

    \I__4021\ : LocalMux
    port map (
            O => \N__18880\,
            I => \N__18863\
        );

    \I__4020\ : LocalMux
    port map (
            O => \N__18873\,
            I => \N__18863\
        );

    \I__4019\ : InMux
    port map (
            O => \N__18872\,
            I => \N__18855\
        );

    \I__4018\ : InMux
    port map (
            O => \N__18871\,
            I => \N__18855\
        );

    \I__4017\ : InMux
    port map (
            O => \N__18870\,
            I => \N__18855\
        );

    \I__4016\ : Span4Mux_v
    port map (
            O => \N__18863\,
            I => \N__18851\
        );

    \I__4015\ : InMux
    port map (
            O => \N__18862\,
            I => \N__18848\
        );

    \I__4014\ : LocalMux
    port map (
            O => \N__18855\,
            I => \N__18845\
        );

    \I__4013\ : InMux
    port map (
            O => \N__18854\,
            I => \N__18840\
        );

    \I__4012\ : Span4Mux_v
    port map (
            O => \N__18851\,
            I => \N__18835\
        );

    \I__4011\ : LocalMux
    port map (
            O => \N__18848\,
            I => \N__18835\
        );

    \I__4010\ : Span4Mux_h
    port map (
            O => \N__18845\,
            I => \N__18832\
        );

    \I__4009\ : InMux
    port map (
            O => \N__18844\,
            I => \N__18827\
        );

    \I__4008\ : InMux
    port map (
            O => \N__18843\,
            I => \N__18827\
        );

    \I__4007\ : LocalMux
    port map (
            O => \N__18840\,
            I => \TVP_VSYNC_buff\
        );

    \I__4006\ : Odrv4
    port map (
            O => \N__18835\,
            I => \TVP_VSYNC_buff\
        );

    \I__4005\ : Odrv4
    port map (
            O => \N__18832\,
            I => \TVP_VSYNC_buff\
        );

    \I__4004\ : LocalMux
    port map (
            O => \N__18827\,
            I => \TVP_VSYNC_buff\
        );

    \I__4003\ : IoInMux
    port map (
            O => \N__18818\,
            I => \N__18815\
        );

    \I__4002\ : LocalMux
    port map (
            O => \N__18815\,
            I => \N__18812\
        );

    \I__4001\ : Span4Mux_s3_h
    port map (
            O => \N__18812\,
            I => \N__18809\
        );

    \I__4000\ : Sp12to4
    port map (
            O => \N__18809\,
            I => \N__18806\
        );

    \I__3999\ : Span12Mux_v
    port map (
            O => \N__18806\,
            I => \N__18802\
        );

    \I__3998\ : InMux
    port map (
            O => \N__18805\,
            I => \N__18799\
        );

    \I__3997\ : Span12Mux_h
    port map (
            O => \N__18802\,
            I => \N__18793\
        );

    \I__3996\ : LocalMux
    port map (
            O => \N__18799\,
            I => \N__18793\
        );

    \I__3995\ : InMux
    port map (
            O => \N__18798\,
            I => \N__18790\
        );

    \I__3994\ : Odrv12
    port map (
            O => \N__18793\,
            I => \DEBUG_c_0\
        );

    \I__3993\ : LocalMux
    port map (
            O => \N__18790\,
            I => \DEBUG_c_0\
        );

    \I__3992\ : CascadeMux
    port map (
            O => \N__18785\,
            I => \N__18781\
        );

    \I__3991\ : CascadeMux
    port map (
            O => \N__18784\,
            I => \N__18778\
        );

    \I__3990\ : InMux
    port map (
            O => \N__18781\,
            I => \N__18772\
        );

    \I__3989\ : InMux
    port map (
            O => \N__18778\,
            I => \N__18772\
        );

    \I__3988\ : CascadeMux
    port map (
            O => \N__18777\,
            I => \N__18769\
        );

    \I__3987\ : LocalMux
    port map (
            O => \N__18772\,
            I => \N__18763\
        );

    \I__3986\ : InMux
    port map (
            O => \N__18769\,
            I => \N__18760\
        );

    \I__3985\ : CascadeMux
    port map (
            O => \N__18768\,
            I => \N__18757\
        );

    \I__3984\ : IoInMux
    port map (
            O => \N__18767\,
            I => \N__18750\
        );

    \I__3983\ : CascadeMux
    port map (
            O => \N__18766\,
            I => \N__18747\
        );

    \I__3982\ : Span4Mux_h
    port map (
            O => \N__18763\,
            I => \N__18744\
        );

    \I__3981\ : LocalMux
    port map (
            O => \N__18760\,
            I => \N__18741\
        );

    \I__3980\ : InMux
    port map (
            O => \N__18757\,
            I => \N__18738\
        );

    \I__3979\ : CascadeMux
    port map (
            O => \N__18756\,
            I => \N__18734\
        );

    \I__3978\ : CascadeMux
    port map (
            O => \N__18755\,
            I => \N__18730\
        );

    \I__3977\ : CascadeMux
    port map (
            O => \N__18754\,
            I => \N__18727\
        );

    \I__3976\ : CascadeMux
    port map (
            O => \N__18753\,
            I => \N__18724\
        );

    \I__3975\ : LocalMux
    port map (
            O => \N__18750\,
            I => \N__18721\
        );

    \I__3974\ : InMux
    port map (
            O => \N__18747\,
            I => \N__18718\
        );

    \I__3973\ : Span4Mux_v
    port map (
            O => \N__18744\,
            I => \N__18713\
        );

    \I__3972\ : Span4Mux_h
    port map (
            O => \N__18741\,
            I => \N__18713\
        );

    \I__3971\ : LocalMux
    port map (
            O => \N__18738\,
            I => \N__18710\
        );

    \I__3970\ : InMux
    port map (
            O => \N__18737\,
            I => \N__18697\
        );

    \I__3969\ : InMux
    port map (
            O => \N__18734\,
            I => \N__18697\
        );

    \I__3968\ : InMux
    port map (
            O => \N__18733\,
            I => \N__18697\
        );

    \I__3967\ : InMux
    port map (
            O => \N__18730\,
            I => \N__18697\
        );

    \I__3966\ : InMux
    port map (
            O => \N__18727\,
            I => \N__18697\
        );

    \I__3965\ : InMux
    port map (
            O => \N__18724\,
            I => \N__18697\
        );

    \I__3964\ : Span12Mux_s1_h
    port map (
            O => \N__18721\,
            I => \N__18694\
        );

    \I__3963\ : LocalMux
    port map (
            O => \N__18718\,
            I => \N__18691\
        );

    \I__3962\ : Span4Mux_v
    port map (
            O => \N__18713\,
            I => \N__18686\
        );

    \I__3961\ : Span4Mux_h
    port map (
            O => \N__18710\,
            I => \N__18686\
        );

    \I__3960\ : LocalMux
    port map (
            O => \N__18697\,
            I => \N__18683\
        );

    \I__3959\ : Span12Mux_h
    port map (
            O => \N__18694\,
            I => \N__18675\
        );

    \I__3958\ : Span12Mux_h
    port map (
            O => \N__18691\,
            I => \N__18675\
        );

    \I__3957\ : Span4Mux_v
    port map (
            O => \N__18686\,
            I => \N__18670\
        );

    \I__3956\ : Span4Mux_h
    port map (
            O => \N__18683\,
            I => \N__18670\
        );

    \I__3955\ : InMux
    port map (
            O => \N__18682\,
            I => \N__18666\
        );

    \I__3954\ : InMux
    port map (
            O => \N__18681\,
            I => \N__18654\
        );

    \I__3953\ : InMux
    port map (
            O => \N__18680\,
            I => \N__18654\
        );

    \I__3952\ : Span12Mux_v
    port map (
            O => \N__18675\,
            I => \N__18651\
        );

    \I__3951\ : Span4Mux_v
    port map (
            O => \N__18670\,
            I => \N__18648\
        );

    \I__3950\ : InMux
    port map (
            O => \N__18669\,
            I => \N__18645\
        );

    \I__3949\ : LocalMux
    port map (
            O => \N__18666\,
            I => \N__18642\
        );

    \I__3948\ : InMux
    port map (
            O => \N__18665\,
            I => \N__18635\
        );

    \I__3947\ : InMux
    port map (
            O => \N__18664\,
            I => \N__18635\
        );

    \I__3946\ : InMux
    port map (
            O => \N__18663\,
            I => \N__18635\
        );

    \I__3945\ : InMux
    port map (
            O => \N__18662\,
            I => \N__18632\
        );

    \I__3944\ : InMux
    port map (
            O => \N__18661\,
            I => \N__18627\
        );

    \I__3943\ : InMux
    port map (
            O => \N__18660\,
            I => \N__18627\
        );

    \I__3942\ : InMux
    port map (
            O => \N__18659\,
            I => \N__18624\
        );

    \I__3941\ : LocalMux
    port map (
            O => \N__18654\,
            I => \N__18621\
        );

    \I__3940\ : Odrv12
    port map (
            O => \N__18651\,
            I => \DEBUG_c_4\
        );

    \I__3939\ : Odrv4
    port map (
            O => \N__18648\,
            I => \DEBUG_c_4\
        );

    \I__3938\ : LocalMux
    port map (
            O => \N__18645\,
            I => \DEBUG_c_4\
        );

    \I__3937\ : Odrv4
    port map (
            O => \N__18642\,
            I => \DEBUG_c_4\
        );

    \I__3936\ : LocalMux
    port map (
            O => \N__18635\,
            I => \DEBUG_c_4\
        );

    \I__3935\ : LocalMux
    port map (
            O => \N__18632\,
            I => \DEBUG_c_4\
        );

    \I__3934\ : LocalMux
    port map (
            O => \N__18627\,
            I => \DEBUG_c_4\
        );

    \I__3933\ : LocalMux
    port map (
            O => \N__18624\,
            I => \DEBUG_c_4\
        );

    \I__3932\ : Odrv4
    port map (
            O => \N__18621\,
            I => \DEBUG_c_4\
        );

    \I__3931\ : InMux
    port map (
            O => \N__18602\,
            I => \N__18599\
        );

    \I__3930\ : LocalMux
    port map (
            O => \N__18599\,
            I => \receive_module.sync_wd.old_visible\
        );

    \I__3929\ : InMux
    port map (
            O => \N__18596\,
            I => \N__18593\
        );

    \I__3928\ : LocalMux
    port map (
            O => \N__18593\,
            I => \N__18588\
        );

    \I__3927\ : InMux
    port map (
            O => \N__18592\,
            I => \N__18585\
        );

    \I__3926\ : InMux
    port map (
            O => \N__18591\,
            I => \N__18582\
        );

    \I__3925\ : Span4Mux_v
    port map (
            O => \N__18588\,
            I => \N__18572\
        );

    \I__3924\ : LocalMux
    port map (
            O => \N__18585\,
            I => \N__18572\
        );

    \I__3923\ : LocalMux
    port map (
            O => \N__18582\,
            I => \N__18572\
        );

    \I__3922\ : InMux
    port map (
            O => \N__18581\,
            I => \N__18569\
        );

    \I__3921\ : InMux
    port map (
            O => \N__18580\,
            I => \N__18566\
        );

    \I__3920\ : InMux
    port map (
            O => \N__18579\,
            I => \N__18563\
        );

    \I__3919\ : Span4Mux_v
    port map (
            O => \N__18572\,
            I => \N__18558\
        );

    \I__3918\ : LocalMux
    port map (
            O => \N__18569\,
            I => \N__18558\
        );

    \I__3917\ : LocalMux
    port map (
            O => \N__18566\,
            I => \N__18553\
        );

    \I__3916\ : LocalMux
    port map (
            O => \N__18563\,
            I => \N__18550\
        );

    \I__3915\ : Span4Mux_v
    port map (
            O => \N__18558\,
            I => \N__18547\
        );

    \I__3914\ : InMux
    port map (
            O => \N__18557\,
            I => \N__18544\
        );

    \I__3913\ : InMux
    port map (
            O => \N__18556\,
            I => \N__18541\
        );

    \I__3912\ : Span12Mux_s10_h
    port map (
            O => \N__18553\,
            I => \N__18538\
        );

    \I__3911\ : Span12Mux_s10_h
    port map (
            O => \N__18550\,
            I => \N__18535\
        );

    \I__3910\ : Span4Mux_h
    port map (
            O => \N__18547\,
            I => \N__18532\
        );

    \I__3909\ : LocalMux
    port map (
            O => \N__18544\,
            I => \N__18529\
        );

    \I__3908\ : LocalMux
    port map (
            O => \N__18541\,
            I => \N__18526\
        );

    \I__3907\ : Span12Mux_v
    port map (
            O => \N__18538\,
            I => \N__18520\
        );

    \I__3906\ : Span12Mux_v
    port map (
            O => \N__18535\,
            I => \N__18520\
        );

    \I__3905\ : Span4Mux_v
    port map (
            O => \N__18532\,
            I => \N__18517\
        );

    \I__3904\ : Span12Mux_h
    port map (
            O => \N__18529\,
            I => \N__18512\
        );

    \I__3903\ : Span12Mux_h
    port map (
            O => \N__18526\,
            I => \N__18512\
        );

    \I__3902\ : InMux
    port map (
            O => \N__18525\,
            I => \N__18509\
        );

    \I__3901\ : Odrv12
    port map (
            O => \N__18520\,
            I => \RX_DATA_7\
        );

    \I__3900\ : Odrv4
    port map (
            O => \N__18517\,
            I => \RX_DATA_7\
        );

    \I__3899\ : Odrv12
    port map (
            O => \N__18512\,
            I => \RX_DATA_7\
        );

    \I__3898\ : LocalMux
    port map (
            O => \N__18509\,
            I => \RX_DATA_7\
        );

    \I__3897\ : InMux
    port map (
            O => \N__18500\,
            I => \N__18497\
        );

    \I__3896\ : LocalMux
    port map (
            O => \N__18497\,
            I => \N__18494\
        );

    \I__3895\ : Span4Mux_v
    port map (
            O => \N__18494\,
            I => \N__18491\
        );

    \I__3894\ : Span4Mux_h
    port map (
            O => \N__18491\,
            I => \N__18488\
        );

    \I__3893\ : Span4Mux_h
    port map (
            O => \N__18488\,
            I => \N__18485\
        );

    \I__3892\ : Odrv4
    port map (
            O => \N__18485\,
            I => \line_buffer.n569\
        );

    \I__3891\ : InMux
    port map (
            O => \N__18482\,
            I => \N__18479\
        );

    \I__3890\ : LocalMux
    port map (
            O => \N__18479\,
            I => \N__18476\
        );

    \I__3889\ : Span4Mux_v
    port map (
            O => \N__18476\,
            I => \N__18473\
        );

    \I__3888\ : Sp12to4
    port map (
            O => \N__18473\,
            I => \N__18470\
        );

    \I__3887\ : Odrv12
    port map (
            O => \N__18470\,
            I => \line_buffer.n561\
        );

    \I__3886\ : InMux
    port map (
            O => \N__18467\,
            I => \N__18464\
        );

    \I__3885\ : LocalMux
    port map (
            O => \N__18464\,
            I => \N__18461\
        );

    \I__3884\ : Span4Mux_v
    port map (
            O => \N__18461\,
            I => \N__18458\
        );

    \I__3883\ : Span4Mux_h
    port map (
            O => \N__18458\,
            I => \N__18455\
        );

    \I__3882\ : Span4Mux_h
    port map (
            O => \N__18455\,
            I => \N__18452\
        );

    \I__3881\ : Odrv4
    port map (
            O => \N__18452\,
            I => \line_buffer.n567\
        );

    \I__3880\ : InMux
    port map (
            O => \N__18449\,
            I => \N__18446\
        );

    \I__3879\ : LocalMux
    port map (
            O => \N__18446\,
            I => \N__18443\
        );

    \I__3878\ : Span12Mux_h
    port map (
            O => \N__18443\,
            I => \N__18440\
        );

    \I__3877\ : Odrv12
    port map (
            O => \N__18440\,
            I => \line_buffer.n559\
        );

    \I__3876\ : CascadeMux
    port map (
            O => \N__18437\,
            I => \receive_module.rx_counter.n3522_cascade_\
        );

    \I__3875\ : InMux
    port map (
            O => \N__18434\,
            I => \N__18431\
        );

    \I__3874\ : LocalMux
    port map (
            O => \N__18431\,
            I => \receive_module.rx_counter.n7_adj_619\
        );

    \I__3873\ : InMux
    port map (
            O => \N__18428\,
            I => \N__18424\
        );

    \I__3872\ : InMux
    port map (
            O => \N__18427\,
            I => \N__18421\
        );

    \I__3871\ : LocalMux
    port map (
            O => \N__18424\,
            I => \receive_module.rx_counter.n11\
        );

    \I__3870\ : LocalMux
    port map (
            O => \N__18421\,
            I => \receive_module.rx_counter.n11\
        );

    \I__3869\ : InMux
    port map (
            O => \N__18416\,
            I => \N__18412\
        );

    \I__3868\ : InMux
    port map (
            O => \N__18415\,
            I => \N__18409\
        );

    \I__3867\ : LocalMux
    port map (
            O => \N__18412\,
            I => \receive_module.rx_counter.FRAME_COUNTER_0\
        );

    \I__3866\ : LocalMux
    port map (
            O => \N__18409\,
            I => \receive_module.rx_counter.FRAME_COUNTER_0\
        );

    \I__3865\ : InMux
    port map (
            O => \N__18404\,
            I => \bfn_16_10_0_\
        );

    \I__3864\ : InMux
    port map (
            O => \N__18401\,
            I => \N__18397\
        );

    \I__3863\ : InMux
    port map (
            O => \N__18400\,
            I => \N__18394\
        );

    \I__3862\ : LocalMux
    port map (
            O => \N__18397\,
            I => \receive_module.rx_counter.FRAME_COUNTER_1\
        );

    \I__3861\ : LocalMux
    port map (
            O => \N__18394\,
            I => \receive_module.rx_counter.FRAME_COUNTER_1\
        );

    \I__3860\ : InMux
    port map (
            O => \N__18389\,
            I => \receive_module.rx_counter.n3205\
        );

    \I__3859\ : InMux
    port map (
            O => \N__18386\,
            I => \N__18382\
        );

    \I__3858\ : InMux
    port map (
            O => \N__18385\,
            I => \N__18379\
        );

    \I__3857\ : LocalMux
    port map (
            O => \N__18382\,
            I => \receive_module.rx_counter.FRAME_COUNTER_2\
        );

    \I__3856\ : LocalMux
    port map (
            O => \N__18379\,
            I => \receive_module.rx_counter.FRAME_COUNTER_2\
        );

    \I__3855\ : InMux
    port map (
            O => \N__18374\,
            I => \receive_module.rx_counter.n3206\
        );

    \I__3854\ : InMux
    port map (
            O => \N__18371\,
            I => \N__18367\
        );

    \I__3853\ : InMux
    port map (
            O => \N__18370\,
            I => \N__18364\
        );

    \I__3852\ : LocalMux
    port map (
            O => \N__18367\,
            I => \receive_module.rx_counter.FRAME_COUNTER_3\
        );

    \I__3851\ : LocalMux
    port map (
            O => \N__18364\,
            I => \receive_module.rx_counter.FRAME_COUNTER_3\
        );

    \I__3850\ : InMux
    port map (
            O => \N__18359\,
            I => \receive_module.rx_counter.n3207\
        );

    \I__3849\ : InMux
    port map (
            O => \N__18356\,
            I => \N__18352\
        );

    \I__3848\ : InMux
    port map (
            O => \N__18355\,
            I => \N__18349\
        );

    \I__3847\ : LocalMux
    port map (
            O => \N__18352\,
            I => \receive_module.rx_counter.FRAME_COUNTER_4\
        );

    \I__3846\ : LocalMux
    port map (
            O => \N__18349\,
            I => \receive_module.rx_counter.FRAME_COUNTER_4\
        );

    \I__3845\ : InMux
    port map (
            O => \N__18344\,
            I => \receive_module.rx_counter.n3208\
        );

    \I__3844\ : InMux
    port map (
            O => \N__18341\,
            I => \receive_module.rx_counter.n3209\
        );

    \I__3843\ : InMux
    port map (
            O => \N__18338\,
            I => \N__18334\
        );

    \I__3842\ : InMux
    port map (
            O => \N__18337\,
            I => \N__18331\
        );

    \I__3841\ : LocalMux
    port map (
            O => \N__18334\,
            I => \receive_module.rx_counter.FRAME_COUNTER_5\
        );

    \I__3840\ : LocalMux
    port map (
            O => \N__18331\,
            I => \receive_module.rx_counter.FRAME_COUNTER_5\
        );

    \I__3839\ : CEMux
    port map (
            O => \N__18326\,
            I => \N__18322\
        );

    \I__3838\ : CEMux
    port map (
            O => \N__18325\,
            I => \N__18319\
        );

    \I__3837\ : LocalMux
    port map (
            O => \N__18322\,
            I => \N__18316\
        );

    \I__3836\ : LocalMux
    port map (
            O => \N__18319\,
            I => \N__18313\
        );

    \I__3835\ : Span4Mux_v
    port map (
            O => \N__18316\,
            I => \N__18310\
        );

    \I__3834\ : Span4Mux_h
    port map (
            O => \N__18313\,
            I => \N__18307\
        );

    \I__3833\ : Odrv4
    port map (
            O => \N__18310\,
            I => \receive_module.rx_counter.n3675\
        );

    \I__3832\ : Odrv4
    port map (
            O => \N__18307\,
            I => \receive_module.rx_counter.n3675\
        );

    \I__3831\ : InMux
    port map (
            O => \N__18302\,
            I => \N__18299\
        );

    \I__3830\ : LocalMux
    port map (
            O => \N__18299\,
            I => \N__18296\
        );

    \I__3829\ : Span12Mux_s9_v
    port map (
            O => \N__18296\,
            I => \N__18293\
        );

    \I__3828\ : Span12Mux_v
    port map (
            O => \N__18293\,
            I => \N__18290\
        );

    \I__3827\ : Odrv12
    port map (
            O => \N__18290\,
            I => \receive_module.n137\
        );

    \I__3826\ : CascadeMux
    port map (
            O => \N__18287\,
            I => \N__18284\
        );

    \I__3825\ : CascadeBuf
    port map (
            O => \N__18284\,
            I => \N__18281\
        );

    \I__3824\ : CascadeMux
    port map (
            O => \N__18281\,
            I => \N__18277\
        );

    \I__3823\ : CascadeMux
    port map (
            O => \N__18280\,
            I => \N__18274\
        );

    \I__3822\ : CascadeBuf
    port map (
            O => \N__18277\,
            I => \N__18271\
        );

    \I__3821\ : CascadeBuf
    port map (
            O => \N__18274\,
            I => \N__18268\
        );

    \I__3820\ : CascadeMux
    port map (
            O => \N__18271\,
            I => \N__18265\
        );

    \I__3819\ : CascadeMux
    port map (
            O => \N__18268\,
            I => \N__18262\
        );

    \I__3818\ : CascadeBuf
    port map (
            O => \N__18265\,
            I => \N__18259\
        );

    \I__3817\ : CascadeBuf
    port map (
            O => \N__18262\,
            I => \N__18256\
        );

    \I__3816\ : CascadeMux
    port map (
            O => \N__18259\,
            I => \N__18253\
        );

    \I__3815\ : CascadeMux
    port map (
            O => \N__18256\,
            I => \N__18250\
        );

    \I__3814\ : CascadeBuf
    port map (
            O => \N__18253\,
            I => \N__18247\
        );

    \I__3813\ : CascadeBuf
    port map (
            O => \N__18250\,
            I => \N__18244\
        );

    \I__3812\ : CascadeMux
    port map (
            O => \N__18247\,
            I => \N__18241\
        );

    \I__3811\ : CascadeMux
    port map (
            O => \N__18244\,
            I => \N__18238\
        );

    \I__3810\ : CascadeBuf
    port map (
            O => \N__18241\,
            I => \N__18235\
        );

    \I__3809\ : CascadeBuf
    port map (
            O => \N__18238\,
            I => \N__18232\
        );

    \I__3808\ : CascadeMux
    port map (
            O => \N__18235\,
            I => \N__18229\
        );

    \I__3807\ : CascadeMux
    port map (
            O => \N__18232\,
            I => \N__18226\
        );

    \I__3806\ : CascadeBuf
    port map (
            O => \N__18229\,
            I => \N__18223\
        );

    \I__3805\ : CascadeBuf
    port map (
            O => \N__18226\,
            I => \N__18220\
        );

    \I__3804\ : CascadeMux
    port map (
            O => \N__18223\,
            I => \N__18217\
        );

    \I__3803\ : CascadeMux
    port map (
            O => \N__18220\,
            I => \N__18214\
        );

    \I__3802\ : CascadeBuf
    port map (
            O => \N__18217\,
            I => \N__18211\
        );

    \I__3801\ : CascadeBuf
    port map (
            O => \N__18214\,
            I => \N__18208\
        );

    \I__3800\ : CascadeMux
    port map (
            O => \N__18211\,
            I => \N__18205\
        );

    \I__3799\ : CascadeMux
    port map (
            O => \N__18208\,
            I => \N__18202\
        );

    \I__3798\ : CascadeBuf
    port map (
            O => \N__18205\,
            I => \N__18199\
        );

    \I__3797\ : CascadeBuf
    port map (
            O => \N__18202\,
            I => \N__18196\
        );

    \I__3796\ : CascadeMux
    port map (
            O => \N__18199\,
            I => \N__18193\
        );

    \I__3795\ : CascadeMux
    port map (
            O => \N__18196\,
            I => \N__18190\
        );

    \I__3794\ : CascadeBuf
    port map (
            O => \N__18193\,
            I => \N__18187\
        );

    \I__3793\ : CascadeBuf
    port map (
            O => \N__18190\,
            I => \N__18184\
        );

    \I__3792\ : CascadeMux
    port map (
            O => \N__18187\,
            I => \N__18181\
        );

    \I__3791\ : CascadeMux
    port map (
            O => \N__18184\,
            I => \N__18178\
        );

    \I__3790\ : CascadeBuf
    port map (
            O => \N__18181\,
            I => \N__18175\
        );

    \I__3789\ : CascadeBuf
    port map (
            O => \N__18178\,
            I => \N__18172\
        );

    \I__3788\ : CascadeMux
    port map (
            O => \N__18175\,
            I => \N__18169\
        );

    \I__3787\ : CascadeMux
    port map (
            O => \N__18172\,
            I => \N__18166\
        );

    \I__3786\ : CascadeBuf
    port map (
            O => \N__18169\,
            I => \N__18163\
        );

    \I__3785\ : CascadeBuf
    port map (
            O => \N__18166\,
            I => \N__18160\
        );

    \I__3784\ : CascadeMux
    port map (
            O => \N__18163\,
            I => \N__18157\
        );

    \I__3783\ : CascadeMux
    port map (
            O => \N__18160\,
            I => \N__18154\
        );

    \I__3782\ : CascadeBuf
    port map (
            O => \N__18157\,
            I => \N__18151\
        );

    \I__3781\ : CascadeBuf
    port map (
            O => \N__18154\,
            I => \N__18148\
        );

    \I__3780\ : CascadeMux
    port map (
            O => \N__18151\,
            I => \N__18145\
        );

    \I__3779\ : CascadeMux
    port map (
            O => \N__18148\,
            I => \N__18142\
        );

    \I__3778\ : CascadeBuf
    port map (
            O => \N__18145\,
            I => \N__18139\
        );

    \I__3777\ : CascadeBuf
    port map (
            O => \N__18142\,
            I => \N__18136\
        );

    \I__3776\ : CascadeMux
    port map (
            O => \N__18139\,
            I => \N__18133\
        );

    \I__3775\ : CascadeMux
    port map (
            O => \N__18136\,
            I => \N__18130\
        );

    \I__3774\ : CascadeBuf
    port map (
            O => \N__18133\,
            I => \N__18127\
        );

    \I__3773\ : CascadeBuf
    port map (
            O => \N__18130\,
            I => \N__18124\
        );

    \I__3772\ : CascadeMux
    port map (
            O => \N__18127\,
            I => \N__18121\
        );

    \I__3771\ : CascadeMux
    port map (
            O => \N__18124\,
            I => \N__18118\
        );

    \I__3770\ : CascadeBuf
    port map (
            O => \N__18121\,
            I => \N__18115\
        );

    \I__3769\ : CascadeBuf
    port map (
            O => \N__18118\,
            I => \N__18112\
        );

    \I__3768\ : CascadeMux
    port map (
            O => \N__18115\,
            I => \N__18109\
        );

    \I__3767\ : CascadeMux
    port map (
            O => \N__18112\,
            I => \N__18106\
        );

    \I__3766\ : InMux
    port map (
            O => \N__18109\,
            I => \N__18103\
        );

    \I__3765\ : CascadeBuf
    port map (
            O => \N__18106\,
            I => \N__18100\
        );

    \I__3764\ : LocalMux
    port map (
            O => \N__18103\,
            I => \N__18096\
        );

    \I__3763\ : CascadeMux
    port map (
            O => \N__18100\,
            I => \N__18093\
        );

    \I__3762\ : InMux
    port map (
            O => \N__18099\,
            I => \N__18090\
        );

    \I__3761\ : Span4Mux_h
    port map (
            O => \N__18096\,
            I => \N__18087\
        );

    \I__3760\ : InMux
    port map (
            O => \N__18093\,
            I => \N__18084\
        );

    \I__3759\ : LocalMux
    port map (
            O => \N__18090\,
            I => \N__18081\
        );

    \I__3758\ : Span4Mux_v
    port map (
            O => \N__18087\,
            I => \N__18077\
        );

    \I__3757\ : LocalMux
    port map (
            O => \N__18084\,
            I => \N__18074\
        );

    \I__3756\ : Span12Mux_v
    port map (
            O => \N__18081\,
            I => \N__18071\
        );

    \I__3755\ : InMux
    port map (
            O => \N__18080\,
            I => \N__18068\
        );

    \I__3754\ : Sp12to4
    port map (
            O => \N__18077\,
            I => \N__18063\
        );

    \I__3753\ : Span12Mux_s4_v
    port map (
            O => \N__18074\,
            I => \N__18063\
        );

    \I__3752\ : Odrv12
    port map (
            O => \N__18071\,
            I => \RX_ADDR_0\
        );

    \I__3751\ : LocalMux
    port map (
            O => \N__18068\,
            I => \RX_ADDR_0\
        );

    \I__3750\ : Odrv12
    port map (
            O => \N__18063\,
            I => \RX_ADDR_0\
        );

    \I__3749\ : InMux
    port map (
            O => \N__18056\,
            I => \N__18053\
        );

    \I__3748\ : LocalMux
    port map (
            O => \N__18053\,
            I => \N__18050\
        );

    \I__3747\ : Span12Mux_s10_v
    port map (
            O => \N__18050\,
            I => \N__18047\
        );

    \I__3746\ : Odrv12
    port map (
            O => \N__18047\,
            I => \receive_module.n134\
        );

    \I__3745\ : CascadeMux
    port map (
            O => \N__18044\,
            I => \N__18040\
        );

    \I__3744\ : CascadeMux
    port map (
            O => \N__18043\,
            I => \N__18037\
        );

    \I__3743\ : CascadeBuf
    port map (
            O => \N__18040\,
            I => \N__18034\
        );

    \I__3742\ : CascadeBuf
    port map (
            O => \N__18037\,
            I => \N__18031\
        );

    \I__3741\ : CascadeMux
    port map (
            O => \N__18034\,
            I => \N__18028\
        );

    \I__3740\ : CascadeMux
    port map (
            O => \N__18031\,
            I => \N__18025\
        );

    \I__3739\ : CascadeBuf
    port map (
            O => \N__18028\,
            I => \N__18022\
        );

    \I__3738\ : CascadeBuf
    port map (
            O => \N__18025\,
            I => \N__18019\
        );

    \I__3737\ : CascadeMux
    port map (
            O => \N__18022\,
            I => \N__18016\
        );

    \I__3736\ : CascadeMux
    port map (
            O => \N__18019\,
            I => \N__18013\
        );

    \I__3735\ : CascadeBuf
    port map (
            O => \N__18016\,
            I => \N__18010\
        );

    \I__3734\ : CascadeBuf
    port map (
            O => \N__18013\,
            I => \N__18007\
        );

    \I__3733\ : CascadeMux
    port map (
            O => \N__18010\,
            I => \N__18004\
        );

    \I__3732\ : CascadeMux
    port map (
            O => \N__18007\,
            I => \N__18001\
        );

    \I__3731\ : CascadeBuf
    port map (
            O => \N__18004\,
            I => \N__17998\
        );

    \I__3730\ : CascadeBuf
    port map (
            O => \N__18001\,
            I => \N__17995\
        );

    \I__3729\ : CascadeMux
    port map (
            O => \N__17998\,
            I => \N__17992\
        );

    \I__3728\ : CascadeMux
    port map (
            O => \N__17995\,
            I => \N__17989\
        );

    \I__3727\ : CascadeBuf
    port map (
            O => \N__17992\,
            I => \N__17986\
        );

    \I__3726\ : CascadeBuf
    port map (
            O => \N__17989\,
            I => \N__17983\
        );

    \I__3725\ : CascadeMux
    port map (
            O => \N__17986\,
            I => \N__17980\
        );

    \I__3724\ : CascadeMux
    port map (
            O => \N__17983\,
            I => \N__17977\
        );

    \I__3723\ : CascadeBuf
    port map (
            O => \N__17980\,
            I => \N__17974\
        );

    \I__3722\ : CascadeBuf
    port map (
            O => \N__17977\,
            I => \N__17971\
        );

    \I__3721\ : CascadeMux
    port map (
            O => \N__17974\,
            I => \N__17968\
        );

    \I__3720\ : CascadeMux
    port map (
            O => \N__17971\,
            I => \N__17965\
        );

    \I__3719\ : CascadeBuf
    port map (
            O => \N__17968\,
            I => \N__17962\
        );

    \I__3718\ : CascadeBuf
    port map (
            O => \N__17965\,
            I => \N__17959\
        );

    \I__3717\ : CascadeMux
    port map (
            O => \N__17962\,
            I => \N__17956\
        );

    \I__3716\ : CascadeMux
    port map (
            O => \N__17959\,
            I => \N__17953\
        );

    \I__3715\ : CascadeBuf
    port map (
            O => \N__17956\,
            I => \N__17950\
        );

    \I__3714\ : CascadeBuf
    port map (
            O => \N__17953\,
            I => \N__17947\
        );

    \I__3713\ : CascadeMux
    port map (
            O => \N__17950\,
            I => \N__17944\
        );

    \I__3712\ : CascadeMux
    port map (
            O => \N__17947\,
            I => \N__17941\
        );

    \I__3711\ : CascadeBuf
    port map (
            O => \N__17944\,
            I => \N__17938\
        );

    \I__3710\ : CascadeBuf
    port map (
            O => \N__17941\,
            I => \N__17935\
        );

    \I__3709\ : CascadeMux
    port map (
            O => \N__17938\,
            I => \N__17932\
        );

    \I__3708\ : CascadeMux
    port map (
            O => \N__17935\,
            I => \N__17929\
        );

    \I__3707\ : CascadeBuf
    port map (
            O => \N__17932\,
            I => \N__17926\
        );

    \I__3706\ : CascadeBuf
    port map (
            O => \N__17929\,
            I => \N__17923\
        );

    \I__3705\ : CascadeMux
    port map (
            O => \N__17926\,
            I => \N__17920\
        );

    \I__3704\ : CascadeMux
    port map (
            O => \N__17923\,
            I => \N__17917\
        );

    \I__3703\ : CascadeBuf
    port map (
            O => \N__17920\,
            I => \N__17914\
        );

    \I__3702\ : CascadeBuf
    port map (
            O => \N__17917\,
            I => \N__17911\
        );

    \I__3701\ : CascadeMux
    port map (
            O => \N__17914\,
            I => \N__17908\
        );

    \I__3700\ : CascadeMux
    port map (
            O => \N__17911\,
            I => \N__17905\
        );

    \I__3699\ : CascadeBuf
    port map (
            O => \N__17908\,
            I => \N__17902\
        );

    \I__3698\ : CascadeBuf
    port map (
            O => \N__17905\,
            I => \N__17899\
        );

    \I__3697\ : CascadeMux
    port map (
            O => \N__17902\,
            I => \N__17896\
        );

    \I__3696\ : CascadeMux
    port map (
            O => \N__17899\,
            I => \N__17893\
        );

    \I__3695\ : CascadeBuf
    port map (
            O => \N__17896\,
            I => \N__17890\
        );

    \I__3694\ : CascadeBuf
    port map (
            O => \N__17893\,
            I => \N__17887\
        );

    \I__3693\ : CascadeMux
    port map (
            O => \N__17890\,
            I => \N__17884\
        );

    \I__3692\ : CascadeMux
    port map (
            O => \N__17887\,
            I => \N__17881\
        );

    \I__3691\ : CascadeBuf
    port map (
            O => \N__17884\,
            I => \N__17878\
        );

    \I__3690\ : CascadeBuf
    port map (
            O => \N__17881\,
            I => \N__17875\
        );

    \I__3689\ : CascadeMux
    port map (
            O => \N__17878\,
            I => \N__17872\
        );

    \I__3688\ : CascadeMux
    port map (
            O => \N__17875\,
            I => \N__17869\
        );

    \I__3687\ : CascadeBuf
    port map (
            O => \N__17872\,
            I => \N__17866\
        );

    \I__3686\ : CascadeBuf
    port map (
            O => \N__17869\,
            I => \N__17863\
        );

    \I__3685\ : CascadeMux
    port map (
            O => \N__17866\,
            I => \N__17859\
        );

    \I__3684\ : CascadeMux
    port map (
            O => \N__17863\,
            I => \N__17856\
        );

    \I__3683\ : InMux
    port map (
            O => \N__17862\,
            I => \N__17853\
        );

    \I__3682\ : InMux
    port map (
            O => \N__17859\,
            I => \N__17850\
        );

    \I__3681\ : InMux
    port map (
            O => \N__17856\,
            I => \N__17847\
        );

    \I__3680\ : LocalMux
    port map (
            O => \N__17853\,
            I => \N__17843\
        );

    \I__3679\ : LocalMux
    port map (
            O => \N__17850\,
            I => \N__17840\
        );

    \I__3678\ : LocalMux
    port map (
            O => \N__17847\,
            I => \N__17837\
        );

    \I__3677\ : InMux
    port map (
            O => \N__17846\,
            I => \N__17834\
        );

    \I__3676\ : Span12Mux_v
    port map (
            O => \N__17843\,
            I => \N__17827\
        );

    \I__3675\ : Span12Mux_h
    port map (
            O => \N__17840\,
            I => \N__17827\
        );

    \I__3674\ : Span12Mux_h
    port map (
            O => \N__17837\,
            I => \N__17827\
        );

    \I__3673\ : LocalMux
    port map (
            O => \N__17834\,
            I => \RX_ADDR_3\
        );

    \I__3672\ : Odrv12
    port map (
            O => \N__17827\,
            I => \RX_ADDR_3\
        );

    \I__3671\ : InMux
    port map (
            O => \N__17822\,
            I => \N__17819\
        );

    \I__3670\ : LocalMux
    port map (
            O => \N__17819\,
            I => \N__17816\
        );

    \I__3669\ : Span12Mux_s10_v
    port map (
            O => \N__17816\,
            I => \N__17813\
        );

    \I__3668\ : Odrv12
    port map (
            O => \N__17813\,
            I => \receive_module.n127\
        );

    \I__3667\ : CascadeMux
    port map (
            O => \N__17810\,
            I => \N__17807\
        );

    \I__3666\ : CascadeBuf
    port map (
            O => \N__17807\,
            I => \N__17803\
        );

    \I__3665\ : CascadeMux
    port map (
            O => \N__17806\,
            I => \N__17800\
        );

    \I__3664\ : CascadeMux
    port map (
            O => \N__17803\,
            I => \N__17797\
        );

    \I__3663\ : CascadeBuf
    port map (
            O => \N__17800\,
            I => \N__17794\
        );

    \I__3662\ : CascadeBuf
    port map (
            O => \N__17797\,
            I => \N__17791\
        );

    \I__3661\ : CascadeMux
    port map (
            O => \N__17794\,
            I => \N__17788\
        );

    \I__3660\ : CascadeMux
    port map (
            O => \N__17791\,
            I => \N__17785\
        );

    \I__3659\ : CascadeBuf
    port map (
            O => \N__17788\,
            I => \N__17782\
        );

    \I__3658\ : CascadeBuf
    port map (
            O => \N__17785\,
            I => \N__17779\
        );

    \I__3657\ : CascadeMux
    port map (
            O => \N__17782\,
            I => \N__17776\
        );

    \I__3656\ : CascadeMux
    port map (
            O => \N__17779\,
            I => \N__17773\
        );

    \I__3655\ : CascadeBuf
    port map (
            O => \N__17776\,
            I => \N__17770\
        );

    \I__3654\ : CascadeBuf
    port map (
            O => \N__17773\,
            I => \N__17767\
        );

    \I__3653\ : CascadeMux
    port map (
            O => \N__17770\,
            I => \N__17764\
        );

    \I__3652\ : CascadeMux
    port map (
            O => \N__17767\,
            I => \N__17761\
        );

    \I__3651\ : CascadeBuf
    port map (
            O => \N__17764\,
            I => \N__17758\
        );

    \I__3650\ : CascadeBuf
    port map (
            O => \N__17761\,
            I => \N__17755\
        );

    \I__3649\ : CascadeMux
    port map (
            O => \N__17758\,
            I => \N__17752\
        );

    \I__3648\ : CascadeMux
    port map (
            O => \N__17755\,
            I => \N__17749\
        );

    \I__3647\ : CascadeBuf
    port map (
            O => \N__17752\,
            I => \N__17746\
        );

    \I__3646\ : CascadeBuf
    port map (
            O => \N__17749\,
            I => \N__17743\
        );

    \I__3645\ : CascadeMux
    port map (
            O => \N__17746\,
            I => \N__17740\
        );

    \I__3644\ : CascadeMux
    port map (
            O => \N__17743\,
            I => \N__17737\
        );

    \I__3643\ : CascadeBuf
    port map (
            O => \N__17740\,
            I => \N__17734\
        );

    \I__3642\ : CascadeBuf
    port map (
            O => \N__17737\,
            I => \N__17731\
        );

    \I__3641\ : CascadeMux
    port map (
            O => \N__17734\,
            I => \N__17728\
        );

    \I__3640\ : CascadeMux
    port map (
            O => \N__17731\,
            I => \N__17725\
        );

    \I__3639\ : CascadeBuf
    port map (
            O => \N__17728\,
            I => \N__17722\
        );

    \I__3638\ : CascadeBuf
    port map (
            O => \N__17725\,
            I => \N__17719\
        );

    \I__3637\ : CascadeMux
    port map (
            O => \N__17722\,
            I => \N__17716\
        );

    \I__3636\ : CascadeMux
    port map (
            O => \N__17719\,
            I => \N__17713\
        );

    \I__3635\ : CascadeBuf
    port map (
            O => \N__17716\,
            I => \N__17710\
        );

    \I__3634\ : CascadeBuf
    port map (
            O => \N__17713\,
            I => \N__17707\
        );

    \I__3633\ : CascadeMux
    port map (
            O => \N__17710\,
            I => \N__17704\
        );

    \I__3632\ : CascadeMux
    port map (
            O => \N__17707\,
            I => \N__17701\
        );

    \I__3631\ : CascadeBuf
    port map (
            O => \N__17704\,
            I => \N__17698\
        );

    \I__3630\ : CascadeBuf
    port map (
            O => \N__17701\,
            I => \N__17695\
        );

    \I__3629\ : CascadeMux
    port map (
            O => \N__17698\,
            I => \N__17692\
        );

    \I__3628\ : CascadeMux
    port map (
            O => \N__17695\,
            I => \N__17689\
        );

    \I__3627\ : CascadeBuf
    port map (
            O => \N__17692\,
            I => \N__17686\
        );

    \I__3626\ : CascadeBuf
    port map (
            O => \N__17689\,
            I => \N__17683\
        );

    \I__3625\ : CascadeMux
    port map (
            O => \N__17686\,
            I => \N__17680\
        );

    \I__3624\ : CascadeMux
    port map (
            O => \N__17683\,
            I => \N__17677\
        );

    \I__3623\ : CascadeBuf
    port map (
            O => \N__17680\,
            I => \N__17674\
        );

    \I__3622\ : CascadeBuf
    port map (
            O => \N__17677\,
            I => \N__17671\
        );

    \I__3621\ : CascadeMux
    port map (
            O => \N__17674\,
            I => \N__17668\
        );

    \I__3620\ : CascadeMux
    port map (
            O => \N__17671\,
            I => \N__17665\
        );

    \I__3619\ : CascadeBuf
    port map (
            O => \N__17668\,
            I => \N__17662\
        );

    \I__3618\ : CascadeBuf
    port map (
            O => \N__17665\,
            I => \N__17659\
        );

    \I__3617\ : CascadeMux
    port map (
            O => \N__17662\,
            I => \N__17656\
        );

    \I__3616\ : CascadeMux
    port map (
            O => \N__17659\,
            I => \N__17653\
        );

    \I__3615\ : CascadeBuf
    port map (
            O => \N__17656\,
            I => \N__17650\
        );

    \I__3614\ : CascadeBuf
    port map (
            O => \N__17653\,
            I => \N__17647\
        );

    \I__3613\ : CascadeMux
    port map (
            O => \N__17650\,
            I => \N__17644\
        );

    \I__3612\ : CascadeMux
    port map (
            O => \N__17647\,
            I => \N__17641\
        );

    \I__3611\ : CascadeBuf
    port map (
            O => \N__17644\,
            I => \N__17638\
        );

    \I__3610\ : CascadeBuf
    port map (
            O => \N__17641\,
            I => \N__17635\
        );

    \I__3609\ : CascadeMux
    port map (
            O => \N__17638\,
            I => \N__17632\
        );

    \I__3608\ : CascadeMux
    port map (
            O => \N__17635\,
            I => \N__17629\
        );

    \I__3607\ : CascadeBuf
    port map (
            O => \N__17632\,
            I => \N__17626\
        );

    \I__3606\ : InMux
    port map (
            O => \N__17629\,
            I => \N__17622\
        );

    \I__3605\ : CascadeMux
    port map (
            O => \N__17626\,
            I => \N__17619\
        );

    \I__3604\ : InMux
    port map (
            O => \N__17625\,
            I => \N__17616\
        );

    \I__3603\ : LocalMux
    port map (
            O => \N__17622\,
            I => \N__17613\
        );

    \I__3602\ : InMux
    port map (
            O => \N__17619\,
            I => \N__17610\
        );

    \I__3601\ : LocalMux
    port map (
            O => \N__17616\,
            I => \N__17607\
        );

    \I__3600\ : Span4Mux_s1_v
    port map (
            O => \N__17613\,
            I => \N__17604\
        );

    \I__3599\ : LocalMux
    port map (
            O => \N__17610\,
            I => \N__17601\
        );

    \I__3598\ : Span12Mux_v
    port map (
            O => \N__17607\,
            I => \N__17598\
        );

    \I__3597\ : Span4Mux_h
    port map (
            O => \N__17604\,
            I => \N__17594\
        );

    \I__3596\ : Span4Mux_s1_v
    port map (
            O => \N__17601\,
            I => \N__17591\
        );

    \I__3595\ : Span12Mux_v
    port map (
            O => \N__17598\,
            I => \N__17588\
        );

    \I__3594\ : InMux
    port map (
            O => \N__17597\,
            I => \N__17585\
        );

    \I__3593\ : Span4Mux_h
    port map (
            O => \N__17594\,
            I => \N__17582\
        );

    \I__3592\ : Span4Mux_h
    port map (
            O => \N__17591\,
            I => \N__17579\
        );

    \I__3591\ : Odrv12
    port map (
            O => \N__17588\,
            I => \RX_ADDR_10\
        );

    \I__3590\ : LocalMux
    port map (
            O => \N__17585\,
            I => \RX_ADDR_10\
        );

    \I__3589\ : Odrv4
    port map (
            O => \N__17582\,
            I => \RX_ADDR_10\
        );

    \I__3588\ : Odrv4
    port map (
            O => \N__17579\,
            I => \RX_ADDR_10\
        );

    \I__3587\ : SRMux
    port map (
            O => \N__17570\,
            I => \N__17567\
        );

    \I__3586\ : LocalMux
    port map (
            O => \N__17567\,
            I => \N__17562\
        );

    \I__3585\ : SRMux
    port map (
            O => \N__17566\,
            I => \N__17559\
        );

    \I__3584\ : SRMux
    port map (
            O => \N__17565\,
            I => \N__17556\
        );

    \I__3583\ : Span4Mux_v
    port map (
            O => \N__17562\,
            I => \N__17549\
        );

    \I__3582\ : LocalMux
    port map (
            O => \N__17559\,
            I => \N__17549\
        );

    \I__3581\ : LocalMux
    port map (
            O => \N__17556\,
            I => \N__17546\
        );

    \I__3580\ : SRMux
    port map (
            O => \N__17555\,
            I => \N__17543\
        );

    \I__3579\ : SRMux
    port map (
            O => \N__17554\,
            I => \N__17538\
        );

    \I__3578\ : Span4Mux_v
    port map (
            O => \N__17549\,
            I => \N__17531\
        );

    \I__3577\ : Span4Mux_v
    port map (
            O => \N__17546\,
            I => \N__17531\
        );

    \I__3576\ : LocalMux
    port map (
            O => \N__17543\,
            I => \N__17531\
        );

    \I__3575\ : SRMux
    port map (
            O => \N__17542\,
            I => \N__17528\
        );

    \I__3574\ : SRMux
    port map (
            O => \N__17541\,
            I => \N__17525\
        );

    \I__3573\ : LocalMux
    port map (
            O => \N__17538\,
            I => \N__17522\
        );

    \I__3572\ : Span4Mux_v
    port map (
            O => \N__17531\,
            I => \N__17517\
        );

    \I__3571\ : LocalMux
    port map (
            O => \N__17528\,
            I => \N__17517\
        );

    \I__3570\ : LocalMux
    port map (
            O => \N__17525\,
            I => \N__17514\
        );

    \I__3569\ : Span4Mux_h
    port map (
            O => \N__17522\,
            I => \N__17510\
        );

    \I__3568\ : Span4Mux_v
    port map (
            O => \N__17517\,
            I => \N__17505\
        );

    \I__3567\ : Span4Mux_h
    port map (
            O => \N__17514\,
            I => \N__17505\
        );

    \I__3566\ : SRMux
    port map (
            O => \N__17513\,
            I => \N__17502\
        );

    \I__3565\ : Odrv4
    port map (
            O => \N__17510\,
            I => \receive_module.n3677\
        );

    \I__3564\ : Odrv4
    port map (
            O => \N__17505\,
            I => \receive_module.n3677\
        );

    \I__3563\ : LocalMux
    port map (
            O => \N__17502\,
            I => \receive_module.n3677\
        );

    \I__3562\ : IoInMux
    port map (
            O => \N__17495\,
            I => \N__17492\
        );

    \I__3561\ : LocalMux
    port map (
            O => \N__17492\,
            I => \N__17489\
        );

    \I__3560\ : Span4Mux_s1_v
    port map (
            O => \N__17489\,
            I => \N__17486\
        );

    \I__3559\ : Span4Mux_v
    port map (
            O => \N__17486\,
            I => \N__17483\
        );

    \I__3558\ : Span4Mux_h
    port map (
            O => \N__17483\,
            I => \N__17480\
        );

    \I__3557\ : Odrv4
    port map (
            O => \N__17480\,
            I => \LED_c\
        );

    \I__3556\ : InMux
    port map (
            O => \N__17477\,
            I => \N__17474\
        );

    \I__3555\ : LocalMux
    port map (
            O => \N__17474\,
            I => \N__17470\
        );

    \I__3554\ : InMux
    port map (
            O => \N__17473\,
            I => \N__17467\
        );

    \I__3553\ : Odrv4
    port map (
            O => \N__17470\,
            I => \PULSE_1HZ\
        );

    \I__3552\ : LocalMux
    port map (
            O => \N__17467\,
            I => \PULSE_1HZ\
        );

    \I__3551\ : InMux
    port map (
            O => \N__17462\,
            I => \N__17456\
        );

    \I__3550\ : InMux
    port map (
            O => \N__17461\,
            I => \N__17456\
        );

    \I__3549\ : LocalMux
    port map (
            O => \N__17456\,
            I => \receive_module.rx_counter.old_VS\
        );

    \I__3548\ : InMux
    port map (
            O => \N__17453\,
            I => \N__17450\
        );

    \I__3547\ : LocalMux
    port map (
            O => \N__17450\,
            I => \N__17447\
        );

    \I__3546\ : Span4Mux_v
    port map (
            O => \N__17447\,
            I => \N__17444\
        );

    \I__3545\ : Span4Mux_v
    port map (
            O => \N__17444\,
            I => \N__17441\
        );

    \I__3544\ : Odrv4
    port map (
            O => \N__17441\,
            I => \receive_module.n133\
        );

    \I__3543\ : CascadeMux
    port map (
            O => \N__17438\,
            I => \N__17434\
        );

    \I__3542\ : CascadeMux
    port map (
            O => \N__17437\,
            I => \N__17431\
        );

    \I__3541\ : CascadeBuf
    port map (
            O => \N__17434\,
            I => \N__17428\
        );

    \I__3540\ : CascadeBuf
    port map (
            O => \N__17431\,
            I => \N__17425\
        );

    \I__3539\ : CascadeMux
    port map (
            O => \N__17428\,
            I => \N__17422\
        );

    \I__3538\ : CascadeMux
    port map (
            O => \N__17425\,
            I => \N__17419\
        );

    \I__3537\ : CascadeBuf
    port map (
            O => \N__17422\,
            I => \N__17416\
        );

    \I__3536\ : CascadeBuf
    port map (
            O => \N__17419\,
            I => \N__17413\
        );

    \I__3535\ : CascadeMux
    port map (
            O => \N__17416\,
            I => \N__17410\
        );

    \I__3534\ : CascadeMux
    port map (
            O => \N__17413\,
            I => \N__17407\
        );

    \I__3533\ : CascadeBuf
    port map (
            O => \N__17410\,
            I => \N__17404\
        );

    \I__3532\ : CascadeBuf
    port map (
            O => \N__17407\,
            I => \N__17401\
        );

    \I__3531\ : CascadeMux
    port map (
            O => \N__17404\,
            I => \N__17398\
        );

    \I__3530\ : CascadeMux
    port map (
            O => \N__17401\,
            I => \N__17395\
        );

    \I__3529\ : CascadeBuf
    port map (
            O => \N__17398\,
            I => \N__17392\
        );

    \I__3528\ : CascadeBuf
    port map (
            O => \N__17395\,
            I => \N__17389\
        );

    \I__3527\ : CascadeMux
    port map (
            O => \N__17392\,
            I => \N__17386\
        );

    \I__3526\ : CascadeMux
    port map (
            O => \N__17389\,
            I => \N__17383\
        );

    \I__3525\ : CascadeBuf
    port map (
            O => \N__17386\,
            I => \N__17380\
        );

    \I__3524\ : CascadeBuf
    port map (
            O => \N__17383\,
            I => \N__17377\
        );

    \I__3523\ : CascadeMux
    port map (
            O => \N__17380\,
            I => \N__17374\
        );

    \I__3522\ : CascadeMux
    port map (
            O => \N__17377\,
            I => \N__17371\
        );

    \I__3521\ : CascadeBuf
    port map (
            O => \N__17374\,
            I => \N__17368\
        );

    \I__3520\ : CascadeBuf
    port map (
            O => \N__17371\,
            I => \N__17365\
        );

    \I__3519\ : CascadeMux
    port map (
            O => \N__17368\,
            I => \N__17362\
        );

    \I__3518\ : CascadeMux
    port map (
            O => \N__17365\,
            I => \N__17359\
        );

    \I__3517\ : CascadeBuf
    port map (
            O => \N__17362\,
            I => \N__17356\
        );

    \I__3516\ : CascadeBuf
    port map (
            O => \N__17359\,
            I => \N__17353\
        );

    \I__3515\ : CascadeMux
    port map (
            O => \N__17356\,
            I => \N__17350\
        );

    \I__3514\ : CascadeMux
    port map (
            O => \N__17353\,
            I => \N__17347\
        );

    \I__3513\ : CascadeBuf
    port map (
            O => \N__17350\,
            I => \N__17344\
        );

    \I__3512\ : CascadeBuf
    port map (
            O => \N__17347\,
            I => \N__17341\
        );

    \I__3511\ : CascadeMux
    port map (
            O => \N__17344\,
            I => \N__17338\
        );

    \I__3510\ : CascadeMux
    port map (
            O => \N__17341\,
            I => \N__17335\
        );

    \I__3509\ : CascadeBuf
    port map (
            O => \N__17338\,
            I => \N__17332\
        );

    \I__3508\ : CascadeBuf
    port map (
            O => \N__17335\,
            I => \N__17329\
        );

    \I__3507\ : CascadeMux
    port map (
            O => \N__17332\,
            I => \N__17326\
        );

    \I__3506\ : CascadeMux
    port map (
            O => \N__17329\,
            I => \N__17323\
        );

    \I__3505\ : CascadeBuf
    port map (
            O => \N__17326\,
            I => \N__17320\
        );

    \I__3504\ : CascadeBuf
    port map (
            O => \N__17323\,
            I => \N__17317\
        );

    \I__3503\ : CascadeMux
    port map (
            O => \N__17320\,
            I => \N__17314\
        );

    \I__3502\ : CascadeMux
    port map (
            O => \N__17317\,
            I => \N__17311\
        );

    \I__3501\ : CascadeBuf
    port map (
            O => \N__17314\,
            I => \N__17308\
        );

    \I__3500\ : CascadeBuf
    port map (
            O => \N__17311\,
            I => \N__17305\
        );

    \I__3499\ : CascadeMux
    port map (
            O => \N__17308\,
            I => \N__17302\
        );

    \I__3498\ : CascadeMux
    port map (
            O => \N__17305\,
            I => \N__17299\
        );

    \I__3497\ : CascadeBuf
    port map (
            O => \N__17302\,
            I => \N__17296\
        );

    \I__3496\ : CascadeBuf
    port map (
            O => \N__17299\,
            I => \N__17293\
        );

    \I__3495\ : CascadeMux
    port map (
            O => \N__17296\,
            I => \N__17290\
        );

    \I__3494\ : CascadeMux
    port map (
            O => \N__17293\,
            I => \N__17287\
        );

    \I__3493\ : CascadeBuf
    port map (
            O => \N__17290\,
            I => \N__17284\
        );

    \I__3492\ : CascadeBuf
    port map (
            O => \N__17287\,
            I => \N__17281\
        );

    \I__3491\ : CascadeMux
    port map (
            O => \N__17284\,
            I => \N__17278\
        );

    \I__3490\ : CascadeMux
    port map (
            O => \N__17281\,
            I => \N__17275\
        );

    \I__3489\ : CascadeBuf
    port map (
            O => \N__17278\,
            I => \N__17272\
        );

    \I__3488\ : CascadeBuf
    port map (
            O => \N__17275\,
            I => \N__17269\
        );

    \I__3487\ : CascadeMux
    port map (
            O => \N__17272\,
            I => \N__17266\
        );

    \I__3486\ : CascadeMux
    port map (
            O => \N__17269\,
            I => \N__17263\
        );

    \I__3485\ : CascadeBuf
    port map (
            O => \N__17266\,
            I => \N__17260\
        );

    \I__3484\ : CascadeBuf
    port map (
            O => \N__17263\,
            I => \N__17257\
        );

    \I__3483\ : CascadeMux
    port map (
            O => \N__17260\,
            I => \N__17254\
        );

    \I__3482\ : CascadeMux
    port map (
            O => \N__17257\,
            I => \N__17251\
        );

    \I__3481\ : InMux
    port map (
            O => \N__17254\,
            I => \N__17248\
        );

    \I__3480\ : InMux
    port map (
            O => \N__17251\,
            I => \N__17245\
        );

    \I__3479\ : LocalMux
    port map (
            O => \N__17248\,
            I => \N__17241\
        );

    \I__3478\ : LocalMux
    port map (
            O => \N__17245\,
            I => \N__17238\
        );

    \I__3477\ : InMux
    port map (
            O => \N__17244\,
            I => \N__17235\
        );

    \I__3476\ : Span4Mux_s1_v
    port map (
            O => \N__17241\,
            I => \N__17232\
        );

    \I__3475\ : Span4Mux_s1_v
    port map (
            O => \N__17238\,
            I => \N__17229\
        );

    \I__3474\ : LocalMux
    port map (
            O => \N__17235\,
            I => \N__17226\
        );

    \I__3473\ : Sp12to4
    port map (
            O => \N__17232\,
            I => \N__17223\
        );

    \I__3472\ : Sp12to4
    port map (
            O => \N__17229\,
            I => \N__17220\
        );

    \I__3471\ : Span4Mux_h
    port map (
            O => \N__17226\,
            I => \N__17216\
        );

    \I__3470\ : Span12Mux_s6_h
    port map (
            O => \N__17223\,
            I => \N__17213\
        );

    \I__3469\ : Span12Mux_s5_h
    port map (
            O => \N__17220\,
            I => \N__17210\
        );

    \I__3468\ : InMux
    port map (
            O => \N__17219\,
            I => \N__17207\
        );

    \I__3467\ : Span4Mux_v
    port map (
            O => \N__17216\,
            I => \N__17204\
        );

    \I__3466\ : Span12Mux_v
    port map (
            O => \N__17213\,
            I => \N__17201\
        );

    \I__3465\ : Span12Mux_v
    port map (
            O => \N__17210\,
            I => \N__17198\
        );

    \I__3464\ : LocalMux
    port map (
            O => \N__17207\,
            I => \RX_ADDR_4\
        );

    \I__3463\ : Odrv4
    port map (
            O => \N__17204\,
            I => \RX_ADDR_4\
        );

    \I__3462\ : Odrv12
    port map (
            O => \N__17201\,
            I => \RX_ADDR_4\
        );

    \I__3461\ : Odrv12
    port map (
            O => \N__17198\,
            I => \RX_ADDR_4\
        );

    \I__3460\ : InMux
    port map (
            O => \N__17189\,
            I => \N__17186\
        );

    \I__3459\ : LocalMux
    port map (
            O => \N__17186\,
            I => \N__17183\
        );

    \I__3458\ : Span12Mux_v
    port map (
            O => \N__17183\,
            I => \N__17180\
        );

    \I__3457\ : Odrv12
    port map (
            O => \N__17180\,
            I => \receive_module.n132\
        );

    \I__3456\ : CascadeMux
    port map (
            O => \N__17177\,
            I => \N__17173\
        );

    \I__3455\ : CascadeMux
    port map (
            O => \N__17176\,
            I => \N__17170\
        );

    \I__3454\ : CascadeBuf
    port map (
            O => \N__17173\,
            I => \N__17167\
        );

    \I__3453\ : CascadeBuf
    port map (
            O => \N__17170\,
            I => \N__17164\
        );

    \I__3452\ : CascadeMux
    port map (
            O => \N__17167\,
            I => \N__17161\
        );

    \I__3451\ : CascadeMux
    port map (
            O => \N__17164\,
            I => \N__17158\
        );

    \I__3450\ : CascadeBuf
    port map (
            O => \N__17161\,
            I => \N__17155\
        );

    \I__3449\ : CascadeBuf
    port map (
            O => \N__17158\,
            I => \N__17152\
        );

    \I__3448\ : CascadeMux
    port map (
            O => \N__17155\,
            I => \N__17149\
        );

    \I__3447\ : CascadeMux
    port map (
            O => \N__17152\,
            I => \N__17146\
        );

    \I__3446\ : CascadeBuf
    port map (
            O => \N__17149\,
            I => \N__17143\
        );

    \I__3445\ : CascadeBuf
    port map (
            O => \N__17146\,
            I => \N__17140\
        );

    \I__3444\ : CascadeMux
    port map (
            O => \N__17143\,
            I => \N__17137\
        );

    \I__3443\ : CascadeMux
    port map (
            O => \N__17140\,
            I => \N__17134\
        );

    \I__3442\ : CascadeBuf
    port map (
            O => \N__17137\,
            I => \N__17131\
        );

    \I__3441\ : CascadeBuf
    port map (
            O => \N__17134\,
            I => \N__17128\
        );

    \I__3440\ : CascadeMux
    port map (
            O => \N__17131\,
            I => \N__17125\
        );

    \I__3439\ : CascadeMux
    port map (
            O => \N__17128\,
            I => \N__17122\
        );

    \I__3438\ : CascadeBuf
    port map (
            O => \N__17125\,
            I => \N__17119\
        );

    \I__3437\ : CascadeBuf
    port map (
            O => \N__17122\,
            I => \N__17116\
        );

    \I__3436\ : CascadeMux
    port map (
            O => \N__17119\,
            I => \N__17113\
        );

    \I__3435\ : CascadeMux
    port map (
            O => \N__17116\,
            I => \N__17110\
        );

    \I__3434\ : CascadeBuf
    port map (
            O => \N__17113\,
            I => \N__17107\
        );

    \I__3433\ : CascadeBuf
    port map (
            O => \N__17110\,
            I => \N__17104\
        );

    \I__3432\ : CascadeMux
    port map (
            O => \N__17107\,
            I => \N__17101\
        );

    \I__3431\ : CascadeMux
    port map (
            O => \N__17104\,
            I => \N__17098\
        );

    \I__3430\ : CascadeBuf
    port map (
            O => \N__17101\,
            I => \N__17095\
        );

    \I__3429\ : CascadeBuf
    port map (
            O => \N__17098\,
            I => \N__17092\
        );

    \I__3428\ : CascadeMux
    port map (
            O => \N__17095\,
            I => \N__17089\
        );

    \I__3427\ : CascadeMux
    port map (
            O => \N__17092\,
            I => \N__17086\
        );

    \I__3426\ : CascadeBuf
    port map (
            O => \N__17089\,
            I => \N__17083\
        );

    \I__3425\ : CascadeBuf
    port map (
            O => \N__17086\,
            I => \N__17080\
        );

    \I__3424\ : CascadeMux
    port map (
            O => \N__17083\,
            I => \N__17077\
        );

    \I__3423\ : CascadeMux
    port map (
            O => \N__17080\,
            I => \N__17074\
        );

    \I__3422\ : CascadeBuf
    port map (
            O => \N__17077\,
            I => \N__17071\
        );

    \I__3421\ : CascadeBuf
    port map (
            O => \N__17074\,
            I => \N__17068\
        );

    \I__3420\ : CascadeMux
    port map (
            O => \N__17071\,
            I => \N__17065\
        );

    \I__3419\ : CascadeMux
    port map (
            O => \N__17068\,
            I => \N__17062\
        );

    \I__3418\ : CascadeBuf
    port map (
            O => \N__17065\,
            I => \N__17059\
        );

    \I__3417\ : CascadeBuf
    port map (
            O => \N__17062\,
            I => \N__17056\
        );

    \I__3416\ : CascadeMux
    port map (
            O => \N__17059\,
            I => \N__17053\
        );

    \I__3415\ : CascadeMux
    port map (
            O => \N__17056\,
            I => \N__17050\
        );

    \I__3414\ : CascadeBuf
    port map (
            O => \N__17053\,
            I => \N__17047\
        );

    \I__3413\ : CascadeBuf
    port map (
            O => \N__17050\,
            I => \N__17044\
        );

    \I__3412\ : CascadeMux
    port map (
            O => \N__17047\,
            I => \N__17041\
        );

    \I__3411\ : CascadeMux
    port map (
            O => \N__17044\,
            I => \N__17038\
        );

    \I__3410\ : CascadeBuf
    port map (
            O => \N__17041\,
            I => \N__17035\
        );

    \I__3409\ : CascadeBuf
    port map (
            O => \N__17038\,
            I => \N__17032\
        );

    \I__3408\ : CascadeMux
    port map (
            O => \N__17035\,
            I => \N__17029\
        );

    \I__3407\ : CascadeMux
    port map (
            O => \N__17032\,
            I => \N__17026\
        );

    \I__3406\ : CascadeBuf
    port map (
            O => \N__17029\,
            I => \N__17023\
        );

    \I__3405\ : CascadeBuf
    port map (
            O => \N__17026\,
            I => \N__17020\
        );

    \I__3404\ : CascadeMux
    port map (
            O => \N__17023\,
            I => \N__17017\
        );

    \I__3403\ : CascadeMux
    port map (
            O => \N__17020\,
            I => \N__17014\
        );

    \I__3402\ : CascadeBuf
    port map (
            O => \N__17017\,
            I => \N__17011\
        );

    \I__3401\ : CascadeBuf
    port map (
            O => \N__17014\,
            I => \N__17008\
        );

    \I__3400\ : CascadeMux
    port map (
            O => \N__17011\,
            I => \N__17005\
        );

    \I__3399\ : CascadeMux
    port map (
            O => \N__17008\,
            I => \N__17002\
        );

    \I__3398\ : CascadeBuf
    port map (
            O => \N__17005\,
            I => \N__16999\
        );

    \I__3397\ : CascadeBuf
    port map (
            O => \N__17002\,
            I => \N__16996\
        );

    \I__3396\ : CascadeMux
    port map (
            O => \N__16999\,
            I => \N__16993\
        );

    \I__3395\ : CascadeMux
    port map (
            O => \N__16996\,
            I => \N__16989\
        );

    \I__3394\ : InMux
    port map (
            O => \N__16993\,
            I => \N__16986\
        );

    \I__3393\ : InMux
    port map (
            O => \N__16992\,
            I => \N__16983\
        );

    \I__3392\ : InMux
    port map (
            O => \N__16989\,
            I => \N__16980\
        );

    \I__3391\ : LocalMux
    port map (
            O => \N__16986\,
            I => \N__16977\
        );

    \I__3390\ : LocalMux
    port map (
            O => \N__16983\,
            I => \N__16973\
        );

    \I__3389\ : LocalMux
    port map (
            O => \N__16980\,
            I => \N__16970\
        );

    \I__3388\ : Span4Mux_h
    port map (
            O => \N__16977\,
            I => \N__16967\
        );

    \I__3387\ : CascadeMux
    port map (
            O => \N__16976\,
            I => \N__16964\
        );

    \I__3386\ : Span4Mux_h
    port map (
            O => \N__16973\,
            I => \N__16961\
        );

    \I__3385\ : Sp12to4
    port map (
            O => \N__16970\,
            I => \N__16958\
        );

    \I__3384\ : Sp12to4
    port map (
            O => \N__16967\,
            I => \N__16955\
        );

    \I__3383\ : InMux
    port map (
            O => \N__16964\,
            I => \N__16952\
        );

    \I__3382\ : Span4Mux_v
    port map (
            O => \N__16961\,
            I => \N__16949\
        );

    \I__3381\ : Span12Mux_v
    port map (
            O => \N__16958\,
            I => \N__16946\
        );

    \I__3380\ : Span12Mux_v
    port map (
            O => \N__16955\,
            I => \N__16943\
        );

    \I__3379\ : LocalMux
    port map (
            O => \N__16952\,
            I => \RX_ADDR_5\
        );

    \I__3378\ : Odrv4
    port map (
            O => \N__16949\,
            I => \RX_ADDR_5\
        );

    \I__3377\ : Odrv12
    port map (
            O => \N__16946\,
            I => \RX_ADDR_5\
        );

    \I__3376\ : Odrv12
    port map (
            O => \N__16943\,
            I => \RX_ADDR_5\
        );

    \I__3375\ : InMux
    port map (
            O => \N__16934\,
            I => \N__16931\
        );

    \I__3374\ : LocalMux
    port map (
            O => \N__16931\,
            I => \N__16928\
        );

    \I__3373\ : Span4Mux_v
    port map (
            O => \N__16928\,
            I => \N__16925\
        );

    \I__3372\ : Span4Mux_v
    port map (
            O => \N__16925\,
            I => \N__16922\
        );

    \I__3371\ : Odrv4
    port map (
            O => \N__16922\,
            I => \receive_module.n131\
        );

    \I__3370\ : CascadeMux
    port map (
            O => \N__16919\,
            I => \N__16915\
        );

    \I__3369\ : CascadeMux
    port map (
            O => \N__16918\,
            I => \N__16912\
        );

    \I__3368\ : CascadeBuf
    port map (
            O => \N__16915\,
            I => \N__16909\
        );

    \I__3367\ : CascadeBuf
    port map (
            O => \N__16912\,
            I => \N__16906\
        );

    \I__3366\ : CascadeMux
    port map (
            O => \N__16909\,
            I => \N__16903\
        );

    \I__3365\ : CascadeMux
    port map (
            O => \N__16906\,
            I => \N__16900\
        );

    \I__3364\ : CascadeBuf
    port map (
            O => \N__16903\,
            I => \N__16897\
        );

    \I__3363\ : CascadeBuf
    port map (
            O => \N__16900\,
            I => \N__16894\
        );

    \I__3362\ : CascadeMux
    port map (
            O => \N__16897\,
            I => \N__16891\
        );

    \I__3361\ : CascadeMux
    port map (
            O => \N__16894\,
            I => \N__16888\
        );

    \I__3360\ : CascadeBuf
    port map (
            O => \N__16891\,
            I => \N__16885\
        );

    \I__3359\ : CascadeBuf
    port map (
            O => \N__16888\,
            I => \N__16882\
        );

    \I__3358\ : CascadeMux
    port map (
            O => \N__16885\,
            I => \N__16879\
        );

    \I__3357\ : CascadeMux
    port map (
            O => \N__16882\,
            I => \N__16876\
        );

    \I__3356\ : CascadeBuf
    port map (
            O => \N__16879\,
            I => \N__16873\
        );

    \I__3355\ : CascadeBuf
    port map (
            O => \N__16876\,
            I => \N__16870\
        );

    \I__3354\ : CascadeMux
    port map (
            O => \N__16873\,
            I => \N__16867\
        );

    \I__3353\ : CascadeMux
    port map (
            O => \N__16870\,
            I => \N__16864\
        );

    \I__3352\ : CascadeBuf
    port map (
            O => \N__16867\,
            I => \N__16861\
        );

    \I__3351\ : CascadeBuf
    port map (
            O => \N__16864\,
            I => \N__16858\
        );

    \I__3350\ : CascadeMux
    port map (
            O => \N__16861\,
            I => \N__16855\
        );

    \I__3349\ : CascadeMux
    port map (
            O => \N__16858\,
            I => \N__16852\
        );

    \I__3348\ : CascadeBuf
    port map (
            O => \N__16855\,
            I => \N__16849\
        );

    \I__3347\ : CascadeBuf
    port map (
            O => \N__16852\,
            I => \N__16846\
        );

    \I__3346\ : CascadeMux
    port map (
            O => \N__16849\,
            I => \N__16843\
        );

    \I__3345\ : CascadeMux
    port map (
            O => \N__16846\,
            I => \N__16840\
        );

    \I__3344\ : CascadeBuf
    port map (
            O => \N__16843\,
            I => \N__16837\
        );

    \I__3343\ : CascadeBuf
    port map (
            O => \N__16840\,
            I => \N__16834\
        );

    \I__3342\ : CascadeMux
    port map (
            O => \N__16837\,
            I => \N__16831\
        );

    \I__3341\ : CascadeMux
    port map (
            O => \N__16834\,
            I => \N__16828\
        );

    \I__3340\ : CascadeBuf
    port map (
            O => \N__16831\,
            I => \N__16825\
        );

    \I__3339\ : CascadeBuf
    port map (
            O => \N__16828\,
            I => \N__16822\
        );

    \I__3338\ : CascadeMux
    port map (
            O => \N__16825\,
            I => \N__16819\
        );

    \I__3337\ : CascadeMux
    port map (
            O => \N__16822\,
            I => \N__16816\
        );

    \I__3336\ : CascadeBuf
    port map (
            O => \N__16819\,
            I => \N__16813\
        );

    \I__3335\ : CascadeBuf
    port map (
            O => \N__16816\,
            I => \N__16810\
        );

    \I__3334\ : CascadeMux
    port map (
            O => \N__16813\,
            I => \N__16807\
        );

    \I__3333\ : CascadeMux
    port map (
            O => \N__16810\,
            I => \N__16804\
        );

    \I__3332\ : CascadeBuf
    port map (
            O => \N__16807\,
            I => \N__16801\
        );

    \I__3331\ : CascadeBuf
    port map (
            O => \N__16804\,
            I => \N__16798\
        );

    \I__3330\ : CascadeMux
    port map (
            O => \N__16801\,
            I => \N__16795\
        );

    \I__3329\ : CascadeMux
    port map (
            O => \N__16798\,
            I => \N__16792\
        );

    \I__3328\ : CascadeBuf
    port map (
            O => \N__16795\,
            I => \N__16789\
        );

    \I__3327\ : CascadeBuf
    port map (
            O => \N__16792\,
            I => \N__16786\
        );

    \I__3326\ : CascadeMux
    port map (
            O => \N__16789\,
            I => \N__16783\
        );

    \I__3325\ : CascadeMux
    port map (
            O => \N__16786\,
            I => \N__16780\
        );

    \I__3324\ : CascadeBuf
    port map (
            O => \N__16783\,
            I => \N__16777\
        );

    \I__3323\ : CascadeBuf
    port map (
            O => \N__16780\,
            I => \N__16774\
        );

    \I__3322\ : CascadeMux
    port map (
            O => \N__16777\,
            I => \N__16771\
        );

    \I__3321\ : CascadeMux
    port map (
            O => \N__16774\,
            I => \N__16768\
        );

    \I__3320\ : CascadeBuf
    port map (
            O => \N__16771\,
            I => \N__16765\
        );

    \I__3319\ : CascadeBuf
    port map (
            O => \N__16768\,
            I => \N__16762\
        );

    \I__3318\ : CascadeMux
    port map (
            O => \N__16765\,
            I => \N__16759\
        );

    \I__3317\ : CascadeMux
    port map (
            O => \N__16762\,
            I => \N__16756\
        );

    \I__3316\ : CascadeBuf
    port map (
            O => \N__16759\,
            I => \N__16753\
        );

    \I__3315\ : CascadeBuf
    port map (
            O => \N__16756\,
            I => \N__16750\
        );

    \I__3314\ : CascadeMux
    port map (
            O => \N__16753\,
            I => \N__16747\
        );

    \I__3313\ : CascadeMux
    port map (
            O => \N__16750\,
            I => \N__16744\
        );

    \I__3312\ : CascadeBuf
    port map (
            O => \N__16747\,
            I => \N__16741\
        );

    \I__3311\ : CascadeBuf
    port map (
            O => \N__16744\,
            I => \N__16738\
        );

    \I__3310\ : CascadeMux
    port map (
            O => \N__16741\,
            I => \N__16735\
        );

    \I__3309\ : CascadeMux
    port map (
            O => \N__16738\,
            I => \N__16732\
        );

    \I__3308\ : InMux
    port map (
            O => \N__16735\,
            I => \N__16729\
        );

    \I__3307\ : InMux
    port map (
            O => \N__16732\,
            I => \N__16726\
        );

    \I__3306\ : LocalMux
    port map (
            O => \N__16729\,
            I => \N__16722\
        );

    \I__3305\ : LocalMux
    port map (
            O => \N__16726\,
            I => \N__16719\
        );

    \I__3304\ : InMux
    port map (
            O => \N__16725\,
            I => \N__16716\
        );

    \I__3303\ : Span4Mux_s3_v
    port map (
            O => \N__16722\,
            I => \N__16713\
        );

    \I__3302\ : Span4Mux_s1_v
    port map (
            O => \N__16719\,
            I => \N__16710\
        );

    \I__3301\ : LocalMux
    port map (
            O => \N__16716\,
            I => \N__16707\
        );

    \I__3300\ : Span4Mux_v
    port map (
            O => \N__16713\,
            I => \N__16704\
        );

    \I__3299\ : Span4Mux_h
    port map (
            O => \N__16710\,
            I => \N__16701\
        );

    \I__3298\ : Span4Mux_v
    port map (
            O => \N__16707\,
            I => \N__16697\
        );

    \I__3297\ : Sp12to4
    port map (
            O => \N__16704\,
            I => \N__16694\
        );

    \I__3296\ : Sp12to4
    port map (
            O => \N__16701\,
            I => \N__16691\
        );

    \I__3295\ : InMux
    port map (
            O => \N__16700\,
            I => \N__16688\
        );

    \I__3294\ : Sp12to4
    port map (
            O => \N__16697\,
            I => \N__16683\
        );

    \I__3293\ : Span12Mux_h
    port map (
            O => \N__16694\,
            I => \N__16683\
        );

    \I__3292\ : Span12Mux_v
    port map (
            O => \N__16691\,
            I => \N__16680\
        );

    \I__3291\ : LocalMux
    port map (
            O => \N__16688\,
            I => \RX_ADDR_6\
        );

    \I__3290\ : Odrv12
    port map (
            O => \N__16683\,
            I => \RX_ADDR_6\
        );

    \I__3289\ : Odrv12
    port map (
            O => \N__16680\,
            I => \RX_ADDR_6\
        );

    \I__3288\ : InMux
    port map (
            O => \N__16673\,
            I => \N__16670\
        );

    \I__3287\ : LocalMux
    port map (
            O => \N__16670\,
            I => \N__16667\
        );

    \I__3286\ : Span4Mux_v
    port map (
            O => \N__16667\,
            I => \N__16664\
        );

    \I__3285\ : Span4Mux_v
    port map (
            O => \N__16664\,
            I => \N__16661\
        );

    \I__3284\ : Odrv4
    port map (
            O => \N__16661\,
            I => \receive_module.n130\
        );

    \I__3283\ : CascadeMux
    port map (
            O => \N__16658\,
            I => \N__16654\
        );

    \I__3282\ : CascadeMux
    port map (
            O => \N__16657\,
            I => \N__16651\
        );

    \I__3281\ : CascadeBuf
    port map (
            O => \N__16654\,
            I => \N__16648\
        );

    \I__3280\ : CascadeBuf
    port map (
            O => \N__16651\,
            I => \N__16645\
        );

    \I__3279\ : CascadeMux
    port map (
            O => \N__16648\,
            I => \N__16642\
        );

    \I__3278\ : CascadeMux
    port map (
            O => \N__16645\,
            I => \N__16639\
        );

    \I__3277\ : CascadeBuf
    port map (
            O => \N__16642\,
            I => \N__16636\
        );

    \I__3276\ : CascadeBuf
    port map (
            O => \N__16639\,
            I => \N__16633\
        );

    \I__3275\ : CascadeMux
    port map (
            O => \N__16636\,
            I => \N__16630\
        );

    \I__3274\ : CascadeMux
    port map (
            O => \N__16633\,
            I => \N__16627\
        );

    \I__3273\ : CascadeBuf
    port map (
            O => \N__16630\,
            I => \N__16624\
        );

    \I__3272\ : CascadeBuf
    port map (
            O => \N__16627\,
            I => \N__16621\
        );

    \I__3271\ : CascadeMux
    port map (
            O => \N__16624\,
            I => \N__16618\
        );

    \I__3270\ : CascadeMux
    port map (
            O => \N__16621\,
            I => \N__16615\
        );

    \I__3269\ : CascadeBuf
    port map (
            O => \N__16618\,
            I => \N__16612\
        );

    \I__3268\ : CascadeBuf
    port map (
            O => \N__16615\,
            I => \N__16609\
        );

    \I__3267\ : CascadeMux
    port map (
            O => \N__16612\,
            I => \N__16606\
        );

    \I__3266\ : CascadeMux
    port map (
            O => \N__16609\,
            I => \N__16603\
        );

    \I__3265\ : CascadeBuf
    port map (
            O => \N__16606\,
            I => \N__16600\
        );

    \I__3264\ : CascadeBuf
    port map (
            O => \N__16603\,
            I => \N__16597\
        );

    \I__3263\ : CascadeMux
    port map (
            O => \N__16600\,
            I => \N__16594\
        );

    \I__3262\ : CascadeMux
    port map (
            O => \N__16597\,
            I => \N__16591\
        );

    \I__3261\ : CascadeBuf
    port map (
            O => \N__16594\,
            I => \N__16588\
        );

    \I__3260\ : CascadeBuf
    port map (
            O => \N__16591\,
            I => \N__16585\
        );

    \I__3259\ : CascadeMux
    port map (
            O => \N__16588\,
            I => \N__16582\
        );

    \I__3258\ : CascadeMux
    port map (
            O => \N__16585\,
            I => \N__16579\
        );

    \I__3257\ : CascadeBuf
    port map (
            O => \N__16582\,
            I => \N__16576\
        );

    \I__3256\ : CascadeBuf
    port map (
            O => \N__16579\,
            I => \N__16573\
        );

    \I__3255\ : CascadeMux
    port map (
            O => \N__16576\,
            I => \N__16570\
        );

    \I__3254\ : CascadeMux
    port map (
            O => \N__16573\,
            I => \N__16567\
        );

    \I__3253\ : CascadeBuf
    port map (
            O => \N__16570\,
            I => \N__16564\
        );

    \I__3252\ : CascadeBuf
    port map (
            O => \N__16567\,
            I => \N__16561\
        );

    \I__3251\ : CascadeMux
    port map (
            O => \N__16564\,
            I => \N__16558\
        );

    \I__3250\ : CascadeMux
    port map (
            O => \N__16561\,
            I => \N__16555\
        );

    \I__3249\ : CascadeBuf
    port map (
            O => \N__16558\,
            I => \N__16552\
        );

    \I__3248\ : CascadeBuf
    port map (
            O => \N__16555\,
            I => \N__16549\
        );

    \I__3247\ : CascadeMux
    port map (
            O => \N__16552\,
            I => \N__16546\
        );

    \I__3246\ : CascadeMux
    port map (
            O => \N__16549\,
            I => \N__16543\
        );

    \I__3245\ : CascadeBuf
    port map (
            O => \N__16546\,
            I => \N__16540\
        );

    \I__3244\ : CascadeBuf
    port map (
            O => \N__16543\,
            I => \N__16537\
        );

    \I__3243\ : CascadeMux
    port map (
            O => \N__16540\,
            I => \N__16534\
        );

    \I__3242\ : CascadeMux
    port map (
            O => \N__16537\,
            I => \N__16531\
        );

    \I__3241\ : CascadeBuf
    port map (
            O => \N__16534\,
            I => \N__16528\
        );

    \I__3240\ : CascadeBuf
    port map (
            O => \N__16531\,
            I => \N__16525\
        );

    \I__3239\ : CascadeMux
    port map (
            O => \N__16528\,
            I => \N__16522\
        );

    \I__3238\ : CascadeMux
    port map (
            O => \N__16525\,
            I => \N__16519\
        );

    \I__3237\ : CascadeBuf
    port map (
            O => \N__16522\,
            I => \N__16516\
        );

    \I__3236\ : CascadeBuf
    port map (
            O => \N__16519\,
            I => \N__16513\
        );

    \I__3235\ : CascadeMux
    port map (
            O => \N__16516\,
            I => \N__16510\
        );

    \I__3234\ : CascadeMux
    port map (
            O => \N__16513\,
            I => \N__16507\
        );

    \I__3233\ : CascadeBuf
    port map (
            O => \N__16510\,
            I => \N__16504\
        );

    \I__3232\ : CascadeBuf
    port map (
            O => \N__16507\,
            I => \N__16501\
        );

    \I__3231\ : CascadeMux
    port map (
            O => \N__16504\,
            I => \N__16498\
        );

    \I__3230\ : CascadeMux
    port map (
            O => \N__16501\,
            I => \N__16495\
        );

    \I__3229\ : CascadeBuf
    port map (
            O => \N__16498\,
            I => \N__16492\
        );

    \I__3228\ : CascadeBuf
    port map (
            O => \N__16495\,
            I => \N__16489\
        );

    \I__3227\ : CascadeMux
    port map (
            O => \N__16492\,
            I => \N__16486\
        );

    \I__3226\ : CascadeMux
    port map (
            O => \N__16489\,
            I => \N__16483\
        );

    \I__3225\ : CascadeBuf
    port map (
            O => \N__16486\,
            I => \N__16480\
        );

    \I__3224\ : CascadeBuf
    port map (
            O => \N__16483\,
            I => \N__16477\
        );

    \I__3223\ : CascadeMux
    port map (
            O => \N__16480\,
            I => \N__16474\
        );

    \I__3222\ : CascadeMux
    port map (
            O => \N__16477\,
            I => \N__16471\
        );

    \I__3221\ : InMux
    port map (
            O => \N__16474\,
            I => \N__16468\
        );

    \I__3220\ : InMux
    port map (
            O => \N__16471\,
            I => \N__16465\
        );

    \I__3219\ : LocalMux
    port map (
            O => \N__16468\,
            I => \N__16461\
        );

    \I__3218\ : LocalMux
    port map (
            O => \N__16465\,
            I => \N__16458\
        );

    \I__3217\ : InMux
    port map (
            O => \N__16464\,
            I => \N__16454\
        );

    \I__3216\ : Span4Mux_h
    port map (
            O => \N__16461\,
            I => \N__16451\
        );

    \I__3215\ : Span4Mux_h
    port map (
            O => \N__16458\,
            I => \N__16448\
        );

    \I__3214\ : CascadeMux
    port map (
            O => \N__16457\,
            I => \N__16445\
        );

    \I__3213\ : LocalMux
    port map (
            O => \N__16454\,
            I => \N__16442\
        );

    \I__3212\ : Sp12to4
    port map (
            O => \N__16451\,
            I => \N__16439\
        );

    \I__3211\ : Sp12to4
    port map (
            O => \N__16448\,
            I => \N__16436\
        );

    \I__3210\ : InMux
    port map (
            O => \N__16445\,
            I => \N__16433\
        );

    \I__3209\ : Span12Mux_v
    port map (
            O => \N__16442\,
            I => \N__16430\
        );

    \I__3208\ : Span12Mux_v
    port map (
            O => \N__16439\,
            I => \N__16425\
        );

    \I__3207\ : Span12Mux_v
    port map (
            O => \N__16436\,
            I => \N__16425\
        );

    \I__3206\ : LocalMux
    port map (
            O => \N__16433\,
            I => \RX_ADDR_7\
        );

    \I__3205\ : Odrv12
    port map (
            O => \N__16430\,
            I => \RX_ADDR_7\
        );

    \I__3204\ : Odrv12
    port map (
            O => \N__16425\,
            I => \RX_ADDR_7\
        );

    \I__3203\ : InMux
    port map (
            O => \N__16418\,
            I => \N__16415\
        );

    \I__3202\ : LocalMux
    port map (
            O => \N__16415\,
            I => \N__16412\
        );

    \I__3201\ : Odrv12
    port map (
            O => \N__16412\,
            I => \transmit_module.ADDR_Y_COMPONENT_3\
        );

    \I__3200\ : InMux
    port map (
            O => \N__16409\,
            I => \N__16406\
        );

    \I__3199\ : LocalMux
    port map (
            O => \N__16406\,
            I => \N__16401\
        );

    \I__3198\ : InMux
    port map (
            O => \N__16405\,
            I => \N__16398\
        );

    \I__3197\ : CascadeMux
    port map (
            O => \N__16404\,
            I => \N__16394\
        );

    \I__3196\ : Span4Mux_v
    port map (
            O => \N__16401\,
            I => \N__16391\
        );

    \I__3195\ : LocalMux
    port map (
            O => \N__16398\,
            I => \N__16388\
        );

    \I__3194\ : InMux
    port map (
            O => \N__16397\,
            I => \N__16385\
        );

    \I__3193\ : InMux
    port map (
            O => \N__16394\,
            I => \N__16382\
        );

    \I__3192\ : Odrv4
    port map (
            O => \N__16391\,
            I => \transmit_module.TX_ADDR_3\
        );

    \I__3191\ : Odrv12
    port map (
            O => \N__16388\,
            I => \transmit_module.TX_ADDR_3\
        );

    \I__3190\ : LocalMux
    port map (
            O => \N__16385\,
            I => \transmit_module.TX_ADDR_3\
        );

    \I__3189\ : LocalMux
    port map (
            O => \N__16382\,
            I => \transmit_module.TX_ADDR_3\
        );

    \I__3188\ : InMux
    port map (
            O => \N__16373\,
            I => \N__16370\
        );

    \I__3187\ : LocalMux
    port map (
            O => \N__16370\,
            I => \N__16367\
        );

    \I__3186\ : Span12Mux_v
    port map (
            O => \N__16367\,
            I => \N__16364\
        );

    \I__3185\ : Odrv12
    port map (
            O => \N__16364\,
            I => \receive_module.n128\
        );

    \I__3184\ : CascadeMux
    port map (
            O => \N__16361\,
            I => \N__16358\
        );

    \I__3183\ : CascadeBuf
    port map (
            O => \N__16358\,
            I => \N__16355\
        );

    \I__3182\ : CascadeMux
    port map (
            O => \N__16355\,
            I => \N__16351\
        );

    \I__3181\ : CascadeMux
    port map (
            O => \N__16354\,
            I => \N__16348\
        );

    \I__3180\ : CascadeBuf
    port map (
            O => \N__16351\,
            I => \N__16345\
        );

    \I__3179\ : CascadeBuf
    port map (
            O => \N__16348\,
            I => \N__16342\
        );

    \I__3178\ : CascadeMux
    port map (
            O => \N__16345\,
            I => \N__16339\
        );

    \I__3177\ : CascadeMux
    port map (
            O => \N__16342\,
            I => \N__16336\
        );

    \I__3176\ : CascadeBuf
    port map (
            O => \N__16339\,
            I => \N__16333\
        );

    \I__3175\ : CascadeBuf
    port map (
            O => \N__16336\,
            I => \N__16330\
        );

    \I__3174\ : CascadeMux
    port map (
            O => \N__16333\,
            I => \N__16327\
        );

    \I__3173\ : CascadeMux
    port map (
            O => \N__16330\,
            I => \N__16324\
        );

    \I__3172\ : CascadeBuf
    port map (
            O => \N__16327\,
            I => \N__16321\
        );

    \I__3171\ : CascadeBuf
    port map (
            O => \N__16324\,
            I => \N__16318\
        );

    \I__3170\ : CascadeMux
    port map (
            O => \N__16321\,
            I => \N__16315\
        );

    \I__3169\ : CascadeMux
    port map (
            O => \N__16318\,
            I => \N__16312\
        );

    \I__3168\ : CascadeBuf
    port map (
            O => \N__16315\,
            I => \N__16309\
        );

    \I__3167\ : CascadeBuf
    port map (
            O => \N__16312\,
            I => \N__16306\
        );

    \I__3166\ : CascadeMux
    port map (
            O => \N__16309\,
            I => \N__16303\
        );

    \I__3165\ : CascadeMux
    port map (
            O => \N__16306\,
            I => \N__16300\
        );

    \I__3164\ : CascadeBuf
    port map (
            O => \N__16303\,
            I => \N__16297\
        );

    \I__3163\ : CascadeBuf
    port map (
            O => \N__16300\,
            I => \N__16294\
        );

    \I__3162\ : CascadeMux
    port map (
            O => \N__16297\,
            I => \N__16291\
        );

    \I__3161\ : CascadeMux
    port map (
            O => \N__16294\,
            I => \N__16288\
        );

    \I__3160\ : CascadeBuf
    port map (
            O => \N__16291\,
            I => \N__16285\
        );

    \I__3159\ : CascadeBuf
    port map (
            O => \N__16288\,
            I => \N__16282\
        );

    \I__3158\ : CascadeMux
    port map (
            O => \N__16285\,
            I => \N__16279\
        );

    \I__3157\ : CascadeMux
    port map (
            O => \N__16282\,
            I => \N__16276\
        );

    \I__3156\ : CascadeBuf
    port map (
            O => \N__16279\,
            I => \N__16273\
        );

    \I__3155\ : CascadeBuf
    port map (
            O => \N__16276\,
            I => \N__16270\
        );

    \I__3154\ : CascadeMux
    port map (
            O => \N__16273\,
            I => \N__16267\
        );

    \I__3153\ : CascadeMux
    port map (
            O => \N__16270\,
            I => \N__16264\
        );

    \I__3152\ : CascadeBuf
    port map (
            O => \N__16267\,
            I => \N__16261\
        );

    \I__3151\ : CascadeBuf
    port map (
            O => \N__16264\,
            I => \N__16258\
        );

    \I__3150\ : CascadeMux
    port map (
            O => \N__16261\,
            I => \N__16255\
        );

    \I__3149\ : CascadeMux
    port map (
            O => \N__16258\,
            I => \N__16252\
        );

    \I__3148\ : CascadeBuf
    port map (
            O => \N__16255\,
            I => \N__16249\
        );

    \I__3147\ : CascadeBuf
    port map (
            O => \N__16252\,
            I => \N__16246\
        );

    \I__3146\ : CascadeMux
    port map (
            O => \N__16249\,
            I => \N__16243\
        );

    \I__3145\ : CascadeMux
    port map (
            O => \N__16246\,
            I => \N__16240\
        );

    \I__3144\ : CascadeBuf
    port map (
            O => \N__16243\,
            I => \N__16237\
        );

    \I__3143\ : CascadeBuf
    port map (
            O => \N__16240\,
            I => \N__16234\
        );

    \I__3142\ : CascadeMux
    port map (
            O => \N__16237\,
            I => \N__16231\
        );

    \I__3141\ : CascadeMux
    port map (
            O => \N__16234\,
            I => \N__16228\
        );

    \I__3140\ : CascadeBuf
    port map (
            O => \N__16231\,
            I => \N__16225\
        );

    \I__3139\ : CascadeBuf
    port map (
            O => \N__16228\,
            I => \N__16222\
        );

    \I__3138\ : CascadeMux
    port map (
            O => \N__16225\,
            I => \N__16219\
        );

    \I__3137\ : CascadeMux
    port map (
            O => \N__16222\,
            I => \N__16216\
        );

    \I__3136\ : CascadeBuf
    port map (
            O => \N__16219\,
            I => \N__16213\
        );

    \I__3135\ : CascadeBuf
    port map (
            O => \N__16216\,
            I => \N__16210\
        );

    \I__3134\ : CascadeMux
    port map (
            O => \N__16213\,
            I => \N__16207\
        );

    \I__3133\ : CascadeMux
    port map (
            O => \N__16210\,
            I => \N__16204\
        );

    \I__3132\ : CascadeBuf
    port map (
            O => \N__16207\,
            I => \N__16201\
        );

    \I__3131\ : CascadeBuf
    port map (
            O => \N__16204\,
            I => \N__16198\
        );

    \I__3130\ : CascadeMux
    port map (
            O => \N__16201\,
            I => \N__16195\
        );

    \I__3129\ : CascadeMux
    port map (
            O => \N__16198\,
            I => \N__16192\
        );

    \I__3128\ : CascadeBuf
    port map (
            O => \N__16195\,
            I => \N__16189\
        );

    \I__3127\ : CascadeBuf
    port map (
            O => \N__16192\,
            I => \N__16186\
        );

    \I__3126\ : CascadeMux
    port map (
            O => \N__16189\,
            I => \N__16183\
        );

    \I__3125\ : CascadeMux
    port map (
            O => \N__16186\,
            I => \N__16180\
        );

    \I__3124\ : InMux
    port map (
            O => \N__16183\,
            I => \N__16177\
        );

    \I__3123\ : CascadeBuf
    port map (
            O => \N__16180\,
            I => \N__16174\
        );

    \I__3122\ : LocalMux
    port map (
            O => \N__16177\,
            I => \N__16170\
        );

    \I__3121\ : CascadeMux
    port map (
            O => \N__16174\,
            I => \N__16167\
        );

    \I__3120\ : InMux
    port map (
            O => \N__16173\,
            I => \N__16164\
        );

    \I__3119\ : Span4Mux_h
    port map (
            O => \N__16170\,
            I => \N__16161\
        );

    \I__3118\ : InMux
    port map (
            O => \N__16167\,
            I => \N__16158\
        );

    \I__3117\ : LocalMux
    port map (
            O => \N__16164\,
            I => \N__16155\
        );

    \I__3116\ : Span4Mux_h
    port map (
            O => \N__16161\,
            I => \N__16152\
        );

    \I__3115\ : LocalMux
    port map (
            O => \N__16158\,
            I => \N__16149\
        );

    \I__3114\ : Span4Mux_v
    port map (
            O => \N__16155\,
            I => \N__16146\
        );

    \I__3113\ : Sp12to4
    port map (
            O => \N__16152\,
            I => \N__16142\
        );

    \I__3112\ : Sp12to4
    port map (
            O => \N__16149\,
            I => \N__16139\
        );

    \I__3111\ : Span4Mux_v
    port map (
            O => \N__16146\,
            I => \N__16136\
        );

    \I__3110\ : InMux
    port map (
            O => \N__16145\,
            I => \N__16133\
        );

    \I__3109\ : Span12Mux_s9_v
    port map (
            O => \N__16142\,
            I => \N__16128\
        );

    \I__3108\ : Span12Mux_s9_v
    port map (
            O => \N__16139\,
            I => \N__16128\
        );

    \I__3107\ : Odrv4
    port map (
            O => \N__16136\,
            I => \RX_ADDR_9\
        );

    \I__3106\ : LocalMux
    port map (
            O => \N__16133\,
            I => \RX_ADDR_9\
        );

    \I__3105\ : Odrv12
    port map (
            O => \N__16128\,
            I => \RX_ADDR_9\
        );

    \I__3104\ : IoInMux
    port map (
            O => \N__16121\,
            I => \N__16117\
        );

    \I__3103\ : IoInMux
    port map (
            O => \N__16120\,
            I => \N__16114\
        );

    \I__3102\ : LocalMux
    port map (
            O => \N__16117\,
            I => \N__16111\
        );

    \I__3101\ : LocalMux
    port map (
            O => \N__16114\,
            I => \N__16108\
        );

    \I__3100\ : Span12Mux_s2_h
    port map (
            O => \N__16111\,
            I => \N__16105\
        );

    \I__3099\ : IoSpan4Mux
    port map (
            O => \N__16108\,
            I => \N__16102\
        );

    \I__3098\ : Span12Mux_v
    port map (
            O => \N__16105\,
            I => \N__16099\
        );

    \I__3097\ : Span4Mux_s1_v
    port map (
            O => \N__16102\,
            I => \N__16096\
        );

    \I__3096\ : Span12Mux_h
    port map (
            O => \N__16099\,
            I => \N__16093\
        );

    \I__3095\ : Span4Mux_v
    port map (
            O => \N__16096\,
            I => \N__16090\
        );

    \I__3094\ : Odrv12
    port map (
            O => \N__16093\,
            I => \GB_BUFFER_DEBUG_c_3_c_THRU_CO\
        );

    \I__3093\ : Odrv4
    port map (
            O => \N__16090\,
            I => \GB_BUFFER_DEBUG_c_3_c_THRU_CO\
        );

    \I__3092\ : IoInMux
    port map (
            O => \N__16085\,
            I => \N__16081\
        );

    \I__3091\ : IoInMux
    port map (
            O => \N__16084\,
            I => \N__16078\
        );

    \I__3090\ : LocalMux
    port map (
            O => \N__16081\,
            I => \N__16075\
        );

    \I__3089\ : LocalMux
    port map (
            O => \N__16078\,
            I => \N__16071\
        );

    \I__3088\ : IoSpan4Mux
    port map (
            O => \N__16075\,
            I => \N__16068\
        );

    \I__3087\ : IoInMux
    port map (
            O => \N__16074\,
            I => \N__16065\
        );

    \I__3086\ : IoSpan4Mux
    port map (
            O => \N__16071\,
            I => \N__16062\
        );

    \I__3085\ : IoSpan4Mux
    port map (
            O => \N__16068\,
            I => \N__16057\
        );

    \I__3084\ : LocalMux
    port map (
            O => \N__16065\,
            I => \N__16057\
        );

    \I__3083\ : Span4Mux_s2_h
    port map (
            O => \N__16062\,
            I => \N__16054\
        );

    \I__3082\ : IoSpan4Mux
    port map (
            O => \N__16057\,
            I => \N__16051\
        );

    \I__3081\ : Sp12to4
    port map (
            O => \N__16054\,
            I => \N__16048\
        );

    \I__3080\ : Span4Mux_s3_v
    port map (
            O => \N__16051\,
            I => \N__16045\
        );

    \I__3079\ : Span12Mux_h
    port map (
            O => \N__16048\,
            I => \N__16042\
        );

    \I__3078\ : Span4Mux_v
    port map (
            O => \N__16045\,
            I => \N__16039\
        );

    \I__3077\ : Odrv12
    port map (
            O => \N__16042\,
            I => n1821
        );

    \I__3076\ : Odrv4
    port map (
            O => \N__16039\,
            I => n1821
        );

    \I__3075\ : InMux
    port map (
            O => \N__16034\,
            I => \N__16031\
        );

    \I__3074\ : LocalMux
    port map (
            O => \N__16031\,
            I => \N__16028\
        );

    \I__3073\ : Span12Mux_v
    port map (
            O => \N__16028\,
            I => \N__16025\
        );

    \I__3072\ : Odrv12
    port map (
            O => \N__16025\,
            I => \receive_module.n129\
        );

    \I__3071\ : CascadeMux
    port map (
            O => \N__16022\,
            I => \N__16018\
        );

    \I__3070\ : CascadeMux
    port map (
            O => \N__16021\,
            I => \N__16015\
        );

    \I__3069\ : CascadeBuf
    port map (
            O => \N__16018\,
            I => \N__16012\
        );

    \I__3068\ : CascadeBuf
    port map (
            O => \N__16015\,
            I => \N__16009\
        );

    \I__3067\ : CascadeMux
    port map (
            O => \N__16012\,
            I => \N__16006\
        );

    \I__3066\ : CascadeMux
    port map (
            O => \N__16009\,
            I => \N__16003\
        );

    \I__3065\ : CascadeBuf
    port map (
            O => \N__16006\,
            I => \N__16000\
        );

    \I__3064\ : CascadeBuf
    port map (
            O => \N__16003\,
            I => \N__15997\
        );

    \I__3063\ : CascadeMux
    port map (
            O => \N__16000\,
            I => \N__15994\
        );

    \I__3062\ : CascadeMux
    port map (
            O => \N__15997\,
            I => \N__15991\
        );

    \I__3061\ : CascadeBuf
    port map (
            O => \N__15994\,
            I => \N__15988\
        );

    \I__3060\ : CascadeBuf
    port map (
            O => \N__15991\,
            I => \N__15985\
        );

    \I__3059\ : CascadeMux
    port map (
            O => \N__15988\,
            I => \N__15982\
        );

    \I__3058\ : CascadeMux
    port map (
            O => \N__15985\,
            I => \N__15979\
        );

    \I__3057\ : CascadeBuf
    port map (
            O => \N__15982\,
            I => \N__15976\
        );

    \I__3056\ : CascadeBuf
    port map (
            O => \N__15979\,
            I => \N__15973\
        );

    \I__3055\ : CascadeMux
    port map (
            O => \N__15976\,
            I => \N__15970\
        );

    \I__3054\ : CascadeMux
    port map (
            O => \N__15973\,
            I => \N__15967\
        );

    \I__3053\ : CascadeBuf
    port map (
            O => \N__15970\,
            I => \N__15964\
        );

    \I__3052\ : CascadeBuf
    port map (
            O => \N__15967\,
            I => \N__15961\
        );

    \I__3051\ : CascadeMux
    port map (
            O => \N__15964\,
            I => \N__15958\
        );

    \I__3050\ : CascadeMux
    port map (
            O => \N__15961\,
            I => \N__15955\
        );

    \I__3049\ : CascadeBuf
    port map (
            O => \N__15958\,
            I => \N__15952\
        );

    \I__3048\ : CascadeBuf
    port map (
            O => \N__15955\,
            I => \N__15949\
        );

    \I__3047\ : CascadeMux
    port map (
            O => \N__15952\,
            I => \N__15946\
        );

    \I__3046\ : CascadeMux
    port map (
            O => \N__15949\,
            I => \N__15943\
        );

    \I__3045\ : CascadeBuf
    port map (
            O => \N__15946\,
            I => \N__15940\
        );

    \I__3044\ : CascadeBuf
    port map (
            O => \N__15943\,
            I => \N__15937\
        );

    \I__3043\ : CascadeMux
    port map (
            O => \N__15940\,
            I => \N__15934\
        );

    \I__3042\ : CascadeMux
    port map (
            O => \N__15937\,
            I => \N__15931\
        );

    \I__3041\ : CascadeBuf
    port map (
            O => \N__15934\,
            I => \N__15928\
        );

    \I__3040\ : CascadeBuf
    port map (
            O => \N__15931\,
            I => \N__15925\
        );

    \I__3039\ : CascadeMux
    port map (
            O => \N__15928\,
            I => \N__15922\
        );

    \I__3038\ : CascadeMux
    port map (
            O => \N__15925\,
            I => \N__15919\
        );

    \I__3037\ : CascadeBuf
    port map (
            O => \N__15922\,
            I => \N__15916\
        );

    \I__3036\ : CascadeBuf
    port map (
            O => \N__15919\,
            I => \N__15913\
        );

    \I__3035\ : CascadeMux
    port map (
            O => \N__15916\,
            I => \N__15910\
        );

    \I__3034\ : CascadeMux
    port map (
            O => \N__15913\,
            I => \N__15907\
        );

    \I__3033\ : CascadeBuf
    port map (
            O => \N__15910\,
            I => \N__15904\
        );

    \I__3032\ : CascadeBuf
    port map (
            O => \N__15907\,
            I => \N__15901\
        );

    \I__3031\ : CascadeMux
    port map (
            O => \N__15904\,
            I => \N__15898\
        );

    \I__3030\ : CascadeMux
    port map (
            O => \N__15901\,
            I => \N__15895\
        );

    \I__3029\ : CascadeBuf
    port map (
            O => \N__15898\,
            I => \N__15892\
        );

    \I__3028\ : CascadeBuf
    port map (
            O => \N__15895\,
            I => \N__15889\
        );

    \I__3027\ : CascadeMux
    port map (
            O => \N__15892\,
            I => \N__15886\
        );

    \I__3026\ : CascadeMux
    port map (
            O => \N__15889\,
            I => \N__15883\
        );

    \I__3025\ : CascadeBuf
    port map (
            O => \N__15886\,
            I => \N__15880\
        );

    \I__3024\ : CascadeBuf
    port map (
            O => \N__15883\,
            I => \N__15877\
        );

    \I__3023\ : CascadeMux
    port map (
            O => \N__15880\,
            I => \N__15874\
        );

    \I__3022\ : CascadeMux
    port map (
            O => \N__15877\,
            I => \N__15871\
        );

    \I__3021\ : CascadeBuf
    port map (
            O => \N__15874\,
            I => \N__15868\
        );

    \I__3020\ : CascadeBuf
    port map (
            O => \N__15871\,
            I => \N__15865\
        );

    \I__3019\ : CascadeMux
    port map (
            O => \N__15868\,
            I => \N__15862\
        );

    \I__3018\ : CascadeMux
    port map (
            O => \N__15865\,
            I => \N__15859\
        );

    \I__3017\ : CascadeBuf
    port map (
            O => \N__15862\,
            I => \N__15856\
        );

    \I__3016\ : CascadeBuf
    port map (
            O => \N__15859\,
            I => \N__15853\
        );

    \I__3015\ : CascadeMux
    port map (
            O => \N__15856\,
            I => \N__15850\
        );

    \I__3014\ : CascadeMux
    port map (
            O => \N__15853\,
            I => \N__15847\
        );

    \I__3013\ : CascadeBuf
    port map (
            O => \N__15850\,
            I => \N__15844\
        );

    \I__3012\ : CascadeBuf
    port map (
            O => \N__15847\,
            I => \N__15841\
        );

    \I__3011\ : CascadeMux
    port map (
            O => \N__15844\,
            I => \N__15838\
        );

    \I__3010\ : CascadeMux
    port map (
            O => \N__15841\,
            I => \N__15835\
        );

    \I__3009\ : InMux
    port map (
            O => \N__15838\,
            I => \N__15832\
        );

    \I__3008\ : InMux
    port map (
            O => \N__15835\,
            I => \N__15829\
        );

    \I__3007\ : LocalMux
    port map (
            O => \N__15832\,
            I => \N__15825\
        );

    \I__3006\ : LocalMux
    port map (
            O => \N__15829\,
            I => \N__15822\
        );

    \I__3005\ : InMux
    port map (
            O => \N__15828\,
            I => \N__15819\
        );

    \I__3004\ : Span4Mux_s1_v
    port map (
            O => \N__15825\,
            I => \N__15816\
        );

    \I__3003\ : Span4Mux_s1_v
    port map (
            O => \N__15822\,
            I => \N__15813\
        );

    \I__3002\ : LocalMux
    port map (
            O => \N__15819\,
            I => \N__15809\
        );

    \I__3001\ : Sp12to4
    port map (
            O => \N__15816\,
            I => \N__15806\
        );

    \I__3000\ : Span4Mux_h
    port map (
            O => \N__15813\,
            I => \N__15803\
        );

    \I__2999\ : InMux
    port map (
            O => \N__15812\,
            I => \N__15800\
        );

    \I__2998\ : Span12Mux_v
    port map (
            O => \N__15809\,
            I => \N__15795\
        );

    \I__2997\ : Span12Mux_h
    port map (
            O => \N__15806\,
            I => \N__15795\
        );

    \I__2996\ : Span4Mux_v
    port map (
            O => \N__15803\,
            I => \N__15792\
        );

    \I__2995\ : LocalMux
    port map (
            O => \N__15800\,
            I => \RX_ADDR_8\
        );

    \I__2994\ : Odrv12
    port map (
            O => \N__15795\,
            I => \RX_ADDR_8\
        );

    \I__2993\ : Odrv4
    port map (
            O => \N__15792\,
            I => \RX_ADDR_8\
        );

    \I__2992\ : CascadeMux
    port map (
            O => \N__15785\,
            I => \transmit_module.n145_cascade_\
        );

    \I__2991\ : InMux
    port map (
            O => \N__15782\,
            I => \N__15779\
        );

    \I__2990\ : LocalMux
    port map (
            O => \N__15779\,
            I => \transmit_module.Y_DELTA_PATTERN_2\
        );

    \I__2989\ : InMux
    port map (
            O => \N__15776\,
            I => \N__15773\
        );

    \I__2988\ : LocalMux
    port map (
            O => \N__15773\,
            I => \N__15770\
        );

    \I__2987\ : Odrv12
    port map (
            O => \N__15770\,
            I => \transmit_module.Y_DELTA_PATTERN_5\
        );

    \I__2986\ : InMux
    port map (
            O => \N__15767\,
            I => \N__15764\
        );

    \I__2985\ : LocalMux
    port map (
            O => \N__15764\,
            I => \transmit_module.Y_DELTA_PATTERN_4\
        );

    \I__2984\ : InMux
    port map (
            O => \N__15761\,
            I => \N__15758\
        );

    \I__2983\ : LocalMux
    port map (
            O => \N__15758\,
            I => \transmit_module.Y_DELTA_PATTERN_3\
        );

    \I__2982\ : InMux
    port map (
            O => \N__15755\,
            I => \N__15752\
        );

    \I__2981\ : LocalMux
    port map (
            O => \N__15752\,
            I => \transmit_module.Y_DELTA_PATTERN_1\
        );

    \I__2980\ : InMux
    port map (
            O => \N__15749\,
            I => \N__15746\
        );

    \I__2979\ : LocalMux
    port map (
            O => \N__15746\,
            I => \N__15743\
        );

    \I__2978\ : Span4Mux_v
    port map (
            O => \N__15743\,
            I => \N__15740\
        );

    \I__2977\ : Span4Mux_v
    port map (
            O => \N__15740\,
            I => \N__15737\
        );

    \I__2976\ : Odrv4
    port map (
            O => \N__15737\,
            I => \receive_module.n136\
        );

    \I__2975\ : CascadeMux
    port map (
            O => \N__15734\,
            I => \N__15730\
        );

    \I__2974\ : CascadeMux
    port map (
            O => \N__15733\,
            I => \N__15727\
        );

    \I__2973\ : CascadeBuf
    port map (
            O => \N__15730\,
            I => \N__15724\
        );

    \I__2972\ : CascadeBuf
    port map (
            O => \N__15727\,
            I => \N__15721\
        );

    \I__2971\ : CascadeMux
    port map (
            O => \N__15724\,
            I => \N__15718\
        );

    \I__2970\ : CascadeMux
    port map (
            O => \N__15721\,
            I => \N__15715\
        );

    \I__2969\ : CascadeBuf
    port map (
            O => \N__15718\,
            I => \N__15712\
        );

    \I__2968\ : CascadeBuf
    port map (
            O => \N__15715\,
            I => \N__15709\
        );

    \I__2967\ : CascadeMux
    port map (
            O => \N__15712\,
            I => \N__15706\
        );

    \I__2966\ : CascadeMux
    port map (
            O => \N__15709\,
            I => \N__15703\
        );

    \I__2965\ : CascadeBuf
    port map (
            O => \N__15706\,
            I => \N__15700\
        );

    \I__2964\ : CascadeBuf
    port map (
            O => \N__15703\,
            I => \N__15697\
        );

    \I__2963\ : CascadeMux
    port map (
            O => \N__15700\,
            I => \N__15694\
        );

    \I__2962\ : CascadeMux
    port map (
            O => \N__15697\,
            I => \N__15691\
        );

    \I__2961\ : CascadeBuf
    port map (
            O => \N__15694\,
            I => \N__15688\
        );

    \I__2960\ : CascadeBuf
    port map (
            O => \N__15691\,
            I => \N__15685\
        );

    \I__2959\ : CascadeMux
    port map (
            O => \N__15688\,
            I => \N__15682\
        );

    \I__2958\ : CascadeMux
    port map (
            O => \N__15685\,
            I => \N__15679\
        );

    \I__2957\ : CascadeBuf
    port map (
            O => \N__15682\,
            I => \N__15676\
        );

    \I__2956\ : CascadeBuf
    port map (
            O => \N__15679\,
            I => \N__15673\
        );

    \I__2955\ : CascadeMux
    port map (
            O => \N__15676\,
            I => \N__15670\
        );

    \I__2954\ : CascadeMux
    port map (
            O => \N__15673\,
            I => \N__15667\
        );

    \I__2953\ : CascadeBuf
    port map (
            O => \N__15670\,
            I => \N__15664\
        );

    \I__2952\ : CascadeBuf
    port map (
            O => \N__15667\,
            I => \N__15661\
        );

    \I__2951\ : CascadeMux
    port map (
            O => \N__15664\,
            I => \N__15658\
        );

    \I__2950\ : CascadeMux
    port map (
            O => \N__15661\,
            I => \N__15655\
        );

    \I__2949\ : CascadeBuf
    port map (
            O => \N__15658\,
            I => \N__15652\
        );

    \I__2948\ : CascadeBuf
    port map (
            O => \N__15655\,
            I => \N__15649\
        );

    \I__2947\ : CascadeMux
    port map (
            O => \N__15652\,
            I => \N__15646\
        );

    \I__2946\ : CascadeMux
    port map (
            O => \N__15649\,
            I => \N__15643\
        );

    \I__2945\ : CascadeBuf
    port map (
            O => \N__15646\,
            I => \N__15640\
        );

    \I__2944\ : CascadeBuf
    port map (
            O => \N__15643\,
            I => \N__15637\
        );

    \I__2943\ : CascadeMux
    port map (
            O => \N__15640\,
            I => \N__15634\
        );

    \I__2942\ : CascadeMux
    port map (
            O => \N__15637\,
            I => \N__15631\
        );

    \I__2941\ : CascadeBuf
    port map (
            O => \N__15634\,
            I => \N__15628\
        );

    \I__2940\ : CascadeBuf
    port map (
            O => \N__15631\,
            I => \N__15625\
        );

    \I__2939\ : CascadeMux
    port map (
            O => \N__15628\,
            I => \N__15622\
        );

    \I__2938\ : CascadeMux
    port map (
            O => \N__15625\,
            I => \N__15619\
        );

    \I__2937\ : CascadeBuf
    port map (
            O => \N__15622\,
            I => \N__15616\
        );

    \I__2936\ : CascadeBuf
    port map (
            O => \N__15619\,
            I => \N__15613\
        );

    \I__2935\ : CascadeMux
    port map (
            O => \N__15616\,
            I => \N__15610\
        );

    \I__2934\ : CascadeMux
    port map (
            O => \N__15613\,
            I => \N__15607\
        );

    \I__2933\ : CascadeBuf
    port map (
            O => \N__15610\,
            I => \N__15604\
        );

    \I__2932\ : CascadeBuf
    port map (
            O => \N__15607\,
            I => \N__15601\
        );

    \I__2931\ : CascadeMux
    port map (
            O => \N__15604\,
            I => \N__15598\
        );

    \I__2930\ : CascadeMux
    port map (
            O => \N__15601\,
            I => \N__15595\
        );

    \I__2929\ : CascadeBuf
    port map (
            O => \N__15598\,
            I => \N__15592\
        );

    \I__2928\ : CascadeBuf
    port map (
            O => \N__15595\,
            I => \N__15589\
        );

    \I__2927\ : CascadeMux
    port map (
            O => \N__15592\,
            I => \N__15586\
        );

    \I__2926\ : CascadeMux
    port map (
            O => \N__15589\,
            I => \N__15583\
        );

    \I__2925\ : CascadeBuf
    port map (
            O => \N__15586\,
            I => \N__15580\
        );

    \I__2924\ : CascadeBuf
    port map (
            O => \N__15583\,
            I => \N__15577\
        );

    \I__2923\ : CascadeMux
    port map (
            O => \N__15580\,
            I => \N__15574\
        );

    \I__2922\ : CascadeMux
    port map (
            O => \N__15577\,
            I => \N__15571\
        );

    \I__2921\ : CascadeBuf
    port map (
            O => \N__15574\,
            I => \N__15568\
        );

    \I__2920\ : CascadeBuf
    port map (
            O => \N__15571\,
            I => \N__15565\
        );

    \I__2919\ : CascadeMux
    port map (
            O => \N__15568\,
            I => \N__15562\
        );

    \I__2918\ : CascadeMux
    port map (
            O => \N__15565\,
            I => \N__15559\
        );

    \I__2917\ : CascadeBuf
    port map (
            O => \N__15562\,
            I => \N__15556\
        );

    \I__2916\ : CascadeBuf
    port map (
            O => \N__15559\,
            I => \N__15553\
        );

    \I__2915\ : CascadeMux
    port map (
            O => \N__15556\,
            I => \N__15550\
        );

    \I__2914\ : CascadeMux
    port map (
            O => \N__15553\,
            I => \N__15547\
        );

    \I__2913\ : InMux
    port map (
            O => \N__15550\,
            I => \N__15544\
        );

    \I__2912\ : InMux
    port map (
            O => \N__15547\,
            I => \N__15541\
        );

    \I__2911\ : LocalMux
    port map (
            O => \N__15544\,
            I => \N__15537\
        );

    \I__2910\ : LocalMux
    port map (
            O => \N__15541\,
            I => \N__15534\
        );

    \I__2909\ : InMux
    port map (
            O => \N__15540\,
            I => \N__15531\
        );

    \I__2908\ : Span4Mux_s1_v
    port map (
            O => \N__15537\,
            I => \N__15528\
        );

    \I__2907\ : Span4Mux_s1_v
    port map (
            O => \N__15534\,
            I => \N__15525\
        );

    \I__2906\ : LocalMux
    port map (
            O => \N__15531\,
            I => \N__15522\
        );

    \I__2905\ : Span4Mux_v
    port map (
            O => \N__15528\,
            I => \N__15519\
        );

    \I__2904\ : Span4Mux_v
    port map (
            O => \N__15525\,
            I => \N__15516\
        );

    \I__2903\ : Span4Mux_v
    port map (
            O => \N__15522\,
            I => \N__15512\
        );

    \I__2902\ : Sp12to4
    port map (
            O => \N__15519\,
            I => \N__15509\
        );

    \I__2901\ : Sp12to4
    port map (
            O => \N__15516\,
            I => \N__15506\
        );

    \I__2900\ : InMux
    port map (
            O => \N__15515\,
            I => \N__15503\
        );

    \I__2899\ : Sp12to4
    port map (
            O => \N__15512\,
            I => \N__15496\
        );

    \I__2898\ : Span12Mux_h
    port map (
            O => \N__15509\,
            I => \N__15496\
        );

    \I__2897\ : Span12Mux_h
    port map (
            O => \N__15506\,
            I => \N__15496\
        );

    \I__2896\ : LocalMux
    port map (
            O => \N__15503\,
            I => \RX_ADDR_1\
        );

    \I__2895\ : Odrv12
    port map (
            O => \N__15496\,
            I => \RX_ADDR_1\
        );

    \I__2894\ : InMux
    port map (
            O => \N__15491\,
            I => \N__15488\
        );

    \I__2893\ : LocalMux
    port map (
            O => \N__15488\,
            I => \N__15485\
        );

    \I__2892\ : Odrv12
    port map (
            O => \N__15485\,
            I => \receive_module.n135\
        );

    \I__2891\ : CascadeMux
    port map (
            O => \N__15482\,
            I => \N__15478\
        );

    \I__2890\ : CascadeMux
    port map (
            O => \N__15481\,
            I => \N__15475\
        );

    \I__2889\ : CascadeBuf
    port map (
            O => \N__15478\,
            I => \N__15472\
        );

    \I__2888\ : CascadeBuf
    port map (
            O => \N__15475\,
            I => \N__15469\
        );

    \I__2887\ : CascadeMux
    port map (
            O => \N__15472\,
            I => \N__15466\
        );

    \I__2886\ : CascadeMux
    port map (
            O => \N__15469\,
            I => \N__15463\
        );

    \I__2885\ : CascadeBuf
    port map (
            O => \N__15466\,
            I => \N__15460\
        );

    \I__2884\ : CascadeBuf
    port map (
            O => \N__15463\,
            I => \N__15457\
        );

    \I__2883\ : CascadeMux
    port map (
            O => \N__15460\,
            I => \N__15454\
        );

    \I__2882\ : CascadeMux
    port map (
            O => \N__15457\,
            I => \N__15451\
        );

    \I__2881\ : CascadeBuf
    port map (
            O => \N__15454\,
            I => \N__15448\
        );

    \I__2880\ : CascadeBuf
    port map (
            O => \N__15451\,
            I => \N__15445\
        );

    \I__2879\ : CascadeMux
    port map (
            O => \N__15448\,
            I => \N__15442\
        );

    \I__2878\ : CascadeMux
    port map (
            O => \N__15445\,
            I => \N__15439\
        );

    \I__2877\ : CascadeBuf
    port map (
            O => \N__15442\,
            I => \N__15436\
        );

    \I__2876\ : CascadeBuf
    port map (
            O => \N__15439\,
            I => \N__15433\
        );

    \I__2875\ : CascadeMux
    port map (
            O => \N__15436\,
            I => \N__15430\
        );

    \I__2874\ : CascadeMux
    port map (
            O => \N__15433\,
            I => \N__15427\
        );

    \I__2873\ : CascadeBuf
    port map (
            O => \N__15430\,
            I => \N__15424\
        );

    \I__2872\ : CascadeBuf
    port map (
            O => \N__15427\,
            I => \N__15421\
        );

    \I__2871\ : CascadeMux
    port map (
            O => \N__15424\,
            I => \N__15418\
        );

    \I__2870\ : CascadeMux
    port map (
            O => \N__15421\,
            I => \N__15415\
        );

    \I__2869\ : CascadeBuf
    port map (
            O => \N__15418\,
            I => \N__15412\
        );

    \I__2868\ : CascadeBuf
    port map (
            O => \N__15415\,
            I => \N__15409\
        );

    \I__2867\ : CascadeMux
    port map (
            O => \N__15412\,
            I => \N__15406\
        );

    \I__2866\ : CascadeMux
    port map (
            O => \N__15409\,
            I => \N__15403\
        );

    \I__2865\ : CascadeBuf
    port map (
            O => \N__15406\,
            I => \N__15400\
        );

    \I__2864\ : CascadeBuf
    port map (
            O => \N__15403\,
            I => \N__15397\
        );

    \I__2863\ : CascadeMux
    port map (
            O => \N__15400\,
            I => \N__15394\
        );

    \I__2862\ : CascadeMux
    port map (
            O => \N__15397\,
            I => \N__15391\
        );

    \I__2861\ : CascadeBuf
    port map (
            O => \N__15394\,
            I => \N__15388\
        );

    \I__2860\ : CascadeBuf
    port map (
            O => \N__15391\,
            I => \N__15385\
        );

    \I__2859\ : CascadeMux
    port map (
            O => \N__15388\,
            I => \N__15382\
        );

    \I__2858\ : CascadeMux
    port map (
            O => \N__15385\,
            I => \N__15379\
        );

    \I__2857\ : CascadeBuf
    port map (
            O => \N__15382\,
            I => \N__15376\
        );

    \I__2856\ : CascadeBuf
    port map (
            O => \N__15379\,
            I => \N__15373\
        );

    \I__2855\ : CascadeMux
    port map (
            O => \N__15376\,
            I => \N__15370\
        );

    \I__2854\ : CascadeMux
    port map (
            O => \N__15373\,
            I => \N__15367\
        );

    \I__2853\ : CascadeBuf
    port map (
            O => \N__15370\,
            I => \N__15364\
        );

    \I__2852\ : CascadeBuf
    port map (
            O => \N__15367\,
            I => \N__15361\
        );

    \I__2851\ : CascadeMux
    port map (
            O => \N__15364\,
            I => \N__15358\
        );

    \I__2850\ : CascadeMux
    port map (
            O => \N__15361\,
            I => \N__15355\
        );

    \I__2849\ : CascadeBuf
    port map (
            O => \N__15358\,
            I => \N__15352\
        );

    \I__2848\ : CascadeBuf
    port map (
            O => \N__15355\,
            I => \N__15349\
        );

    \I__2847\ : CascadeMux
    port map (
            O => \N__15352\,
            I => \N__15346\
        );

    \I__2846\ : CascadeMux
    port map (
            O => \N__15349\,
            I => \N__15343\
        );

    \I__2845\ : CascadeBuf
    port map (
            O => \N__15346\,
            I => \N__15340\
        );

    \I__2844\ : CascadeBuf
    port map (
            O => \N__15343\,
            I => \N__15337\
        );

    \I__2843\ : CascadeMux
    port map (
            O => \N__15340\,
            I => \N__15334\
        );

    \I__2842\ : CascadeMux
    port map (
            O => \N__15337\,
            I => \N__15331\
        );

    \I__2841\ : CascadeBuf
    port map (
            O => \N__15334\,
            I => \N__15328\
        );

    \I__2840\ : CascadeBuf
    port map (
            O => \N__15331\,
            I => \N__15325\
        );

    \I__2839\ : CascadeMux
    port map (
            O => \N__15328\,
            I => \N__15322\
        );

    \I__2838\ : CascadeMux
    port map (
            O => \N__15325\,
            I => \N__15319\
        );

    \I__2837\ : CascadeBuf
    port map (
            O => \N__15322\,
            I => \N__15316\
        );

    \I__2836\ : CascadeBuf
    port map (
            O => \N__15319\,
            I => \N__15313\
        );

    \I__2835\ : CascadeMux
    port map (
            O => \N__15316\,
            I => \N__15310\
        );

    \I__2834\ : CascadeMux
    port map (
            O => \N__15313\,
            I => \N__15307\
        );

    \I__2833\ : CascadeBuf
    port map (
            O => \N__15310\,
            I => \N__15304\
        );

    \I__2832\ : CascadeBuf
    port map (
            O => \N__15307\,
            I => \N__15301\
        );

    \I__2831\ : CascadeMux
    port map (
            O => \N__15304\,
            I => \N__15298\
        );

    \I__2830\ : CascadeMux
    port map (
            O => \N__15301\,
            I => \N__15295\
        );

    \I__2829\ : InMux
    port map (
            O => \N__15298\,
            I => \N__15292\
        );

    \I__2828\ : InMux
    port map (
            O => \N__15295\,
            I => \N__15289\
        );

    \I__2827\ : LocalMux
    port map (
            O => \N__15292\,
            I => \N__15285\
        );

    \I__2826\ : LocalMux
    port map (
            O => \N__15289\,
            I => \N__15282\
        );

    \I__2825\ : InMux
    port map (
            O => \N__15288\,
            I => \N__15279\
        );

    \I__2824\ : Span4Mux_s3_v
    port map (
            O => \N__15285\,
            I => \N__15276\
        );

    \I__2823\ : Span4Mux_s3_v
    port map (
            O => \N__15282\,
            I => \N__15273\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__15279\,
            I => \N__15269\
        );

    \I__2821\ : Sp12to4
    port map (
            O => \N__15276\,
            I => \N__15266\
        );

    \I__2820\ : Sp12to4
    port map (
            O => \N__15273\,
            I => \N__15263\
        );

    \I__2819\ : InMux
    port map (
            O => \N__15272\,
            I => \N__15260\
        );

    \I__2818\ : Span12Mux_v
    port map (
            O => \N__15269\,
            I => \N__15255\
        );

    \I__2817\ : Span12Mux_h
    port map (
            O => \N__15266\,
            I => \N__15255\
        );

    \I__2816\ : Span12Mux_v
    port map (
            O => \N__15263\,
            I => \N__15252\
        );

    \I__2815\ : LocalMux
    port map (
            O => \N__15260\,
            I => \RX_ADDR_2\
        );

    \I__2814\ : Odrv12
    port map (
            O => \N__15255\,
            I => \RX_ADDR_2\
        );

    \I__2813\ : Odrv12
    port map (
            O => \N__15252\,
            I => \RX_ADDR_2\
        );

    \I__2812\ : InMux
    port map (
            O => \N__15245\,
            I => \N__15242\
        );

    \I__2811\ : LocalMux
    port map (
            O => \N__15242\,
            I => \transmit_module.X_DELTA_PATTERN_1\
        );

    \I__2810\ : InMux
    port map (
            O => \N__15239\,
            I => \N__15236\
        );

    \I__2809\ : LocalMux
    port map (
            O => \N__15236\,
            I => \N__15233\
        );

    \I__2808\ : Odrv12
    port map (
            O => \N__15233\,
            I => \transmit_module.X_DELTA_PATTERN_8\
        );

    \I__2807\ : InMux
    port map (
            O => \N__15230\,
            I => \N__15227\
        );

    \I__2806\ : LocalMux
    port map (
            O => \N__15227\,
            I => \transmit_module.X_DELTA_PATTERN_2\
        );

    \I__2805\ : InMux
    port map (
            O => \N__15224\,
            I => \N__15221\
        );

    \I__2804\ : LocalMux
    port map (
            O => \N__15221\,
            I => \transmit_module.X_DELTA_PATTERN_3\
        );

    \I__2803\ : InMux
    port map (
            O => \N__15218\,
            I => \N__15215\
        );

    \I__2802\ : LocalMux
    port map (
            O => \N__15215\,
            I => \transmit_module.X_DELTA_PATTERN_7\
        );

    \I__2801\ : InMux
    port map (
            O => \N__15212\,
            I => \N__15209\
        );

    \I__2800\ : LocalMux
    port map (
            O => \N__15209\,
            I => \transmit_module.X_DELTA_PATTERN_4\
        );

    \I__2799\ : InMux
    port map (
            O => \N__15206\,
            I => \N__15203\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__15203\,
            I => \transmit_module.n129\
        );

    \I__2797\ : InMux
    port map (
            O => \N__15200\,
            I => \N__15196\
        );

    \I__2796\ : InMux
    port map (
            O => \N__15199\,
            I => \N__15193\
        );

    \I__2795\ : LocalMux
    port map (
            O => \N__15196\,
            I => \transmit_module.n110\
        );

    \I__2794\ : LocalMux
    port map (
            O => \N__15193\,
            I => \transmit_module.n110\
        );

    \I__2793\ : InMux
    port map (
            O => \N__15188\,
            I => \N__15185\
        );

    \I__2792\ : LocalMux
    port map (
            O => \N__15185\,
            I => \N__15182\
        );

    \I__2791\ : Odrv4
    port map (
            O => \N__15182\,
            I => \transmit_module.n141\
        );

    \I__2790\ : InMux
    port map (
            O => \N__15179\,
            I => \N__15176\
        );

    \I__2789\ : LocalMux
    port map (
            O => \N__15176\,
            I => \N__15170\
        );

    \I__2788\ : InMux
    port map (
            O => \N__15175\,
            I => \N__15167\
        );

    \I__2787\ : CascadeMux
    port map (
            O => \N__15174\,
            I => \N__15164\
        );

    \I__2786\ : InMux
    port map (
            O => \N__15173\,
            I => \N__15161\
        );

    \I__2785\ : Span4Mux_v
    port map (
            O => \N__15170\,
            I => \N__15156\
        );

    \I__2784\ : LocalMux
    port map (
            O => \N__15167\,
            I => \N__15156\
        );

    \I__2783\ : InMux
    port map (
            O => \N__15164\,
            I => \N__15153\
        );

    \I__2782\ : LocalMux
    port map (
            O => \N__15161\,
            I => \transmit_module.TX_ADDR_6\
        );

    \I__2781\ : Odrv4
    port map (
            O => \N__15156\,
            I => \transmit_module.TX_ADDR_6\
        );

    \I__2780\ : LocalMux
    port map (
            O => \N__15153\,
            I => \transmit_module.TX_ADDR_6\
        );

    \I__2779\ : InMux
    port map (
            O => \N__15146\,
            I => \N__15137\
        );

    \I__2778\ : InMux
    port map (
            O => \N__15145\,
            I => \N__15134\
        );

    \I__2777\ : InMux
    port map (
            O => \N__15144\,
            I => \N__15131\
        );

    \I__2776\ : CascadeMux
    port map (
            O => \N__15143\,
            I => \N__15128\
        );

    \I__2775\ : InMux
    port map (
            O => \N__15142\,
            I => \N__15123\
        );

    \I__2774\ : InMux
    port map (
            O => \N__15141\,
            I => \N__15120\
        );

    \I__2773\ : InMux
    port map (
            O => \N__15140\,
            I => \N__15116\
        );

    \I__2772\ : LocalMux
    port map (
            O => \N__15137\,
            I => \N__15111\
        );

    \I__2771\ : LocalMux
    port map (
            O => \N__15134\,
            I => \N__15106\
        );

    \I__2770\ : LocalMux
    port map (
            O => \N__15131\,
            I => \N__15106\
        );

    \I__2769\ : InMux
    port map (
            O => \N__15128\,
            I => \N__15103\
        );

    \I__2768\ : InMux
    port map (
            O => \N__15127\,
            I => \N__15098\
        );

    \I__2767\ : InMux
    port map (
            O => \N__15126\,
            I => \N__15098\
        );

    \I__2766\ : LocalMux
    port map (
            O => \N__15123\,
            I => \N__15093\
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__15120\,
            I => \N__15090\
        );

    \I__2764\ : InMux
    port map (
            O => \N__15119\,
            I => \N__15087\
        );

    \I__2763\ : LocalMux
    port map (
            O => \N__15116\,
            I => \N__15084\
        );

    \I__2762\ : InMux
    port map (
            O => \N__15115\,
            I => \N__15081\
        );

    \I__2761\ : InMux
    port map (
            O => \N__15114\,
            I => \N__15078\
        );

    \I__2760\ : Span4Mux_h
    port map (
            O => \N__15111\,
            I => \N__15069\
        );

    \I__2759\ : Span4Mux_v
    port map (
            O => \N__15106\,
            I => \N__15069\
        );

    \I__2758\ : LocalMux
    port map (
            O => \N__15103\,
            I => \N__15069\
        );

    \I__2757\ : LocalMux
    port map (
            O => \N__15098\,
            I => \N__15069\
        );

    \I__2756\ : InMux
    port map (
            O => \N__15097\,
            I => \N__15066\
        );

    \I__2755\ : InMux
    port map (
            O => \N__15096\,
            I => \N__15063\
        );

    \I__2754\ : Odrv4
    port map (
            O => \N__15093\,
            I => \transmit_module.VGA_VISIBLE\
        );

    \I__2753\ : Odrv4
    port map (
            O => \N__15090\,
            I => \transmit_module.VGA_VISIBLE\
        );

    \I__2752\ : LocalMux
    port map (
            O => \N__15087\,
            I => \transmit_module.VGA_VISIBLE\
        );

    \I__2751\ : Odrv4
    port map (
            O => \N__15084\,
            I => \transmit_module.VGA_VISIBLE\
        );

    \I__2750\ : LocalMux
    port map (
            O => \N__15081\,
            I => \transmit_module.VGA_VISIBLE\
        );

    \I__2749\ : LocalMux
    port map (
            O => \N__15078\,
            I => \transmit_module.VGA_VISIBLE\
        );

    \I__2748\ : Odrv4
    port map (
            O => \N__15069\,
            I => \transmit_module.VGA_VISIBLE\
        );

    \I__2747\ : LocalMux
    port map (
            O => \N__15066\,
            I => \transmit_module.VGA_VISIBLE\
        );

    \I__2746\ : LocalMux
    port map (
            O => \N__15063\,
            I => \transmit_module.VGA_VISIBLE\
        );

    \I__2745\ : InMux
    port map (
            O => \N__15044\,
            I => \N__15041\
        );

    \I__2744\ : LocalMux
    port map (
            O => \N__15041\,
            I => \transmit_module.n130\
        );

    \I__2743\ : InMux
    port map (
            O => \N__15038\,
            I => \receive_module.n3161\
        );

    \I__2742\ : SRMux
    port map (
            O => \N__15035\,
            I => \N__15032\
        );

    \I__2741\ : LocalMux
    port map (
            O => \N__15032\,
            I => \N__15028\
        );

    \I__2740\ : SRMux
    port map (
            O => \N__15031\,
            I => \N__15025\
        );

    \I__2739\ : Span4Mux_v
    port map (
            O => \N__15028\,
            I => \N__15019\
        );

    \I__2738\ : LocalMux
    port map (
            O => \N__15025\,
            I => \N__15019\
        );

    \I__2737\ : SRMux
    port map (
            O => \N__15024\,
            I => \N__15016\
        );

    \I__2736\ : Span4Mux_v
    port map (
            O => \N__15019\,
            I => \N__15010\
        );

    \I__2735\ : LocalMux
    port map (
            O => \N__15016\,
            I => \N__15010\
        );

    \I__2734\ : SRMux
    port map (
            O => \N__15015\,
            I => \N__15007\
        );

    \I__2733\ : Span4Mux_v
    port map (
            O => \N__15010\,
            I => \N__15002\
        );

    \I__2732\ : LocalMux
    port map (
            O => \N__15007\,
            I => \N__15002\
        );

    \I__2731\ : Span4Mux_h
    port map (
            O => \N__15002\,
            I => \N__14999\
        );

    \I__2730\ : Span4Mux_h
    port map (
            O => \N__14999\,
            I => \N__14996\
        );

    \I__2729\ : Odrv4
    port map (
            O => \N__14996\,
            I => \line_buffer.n606\
        );

    \I__2728\ : SRMux
    port map (
            O => \N__14993\,
            I => \N__14989\
        );

    \I__2727\ : SRMux
    port map (
            O => \N__14992\,
            I => \N__14984\
        );

    \I__2726\ : LocalMux
    port map (
            O => \N__14989\,
            I => \N__14981\
        );

    \I__2725\ : SRMux
    port map (
            O => \N__14988\,
            I => \N__14978\
        );

    \I__2724\ : SRMux
    port map (
            O => \N__14987\,
            I => \N__14975\
        );

    \I__2723\ : LocalMux
    port map (
            O => \N__14984\,
            I => \N__14972\
        );

    \I__2722\ : Span4Mux_s2_v
    port map (
            O => \N__14981\,
            I => \N__14965\
        );

    \I__2721\ : LocalMux
    port map (
            O => \N__14978\,
            I => \N__14965\
        );

    \I__2720\ : LocalMux
    port map (
            O => \N__14975\,
            I => \N__14965\
        );

    \I__2719\ : Span4Mux_h
    port map (
            O => \N__14972\,
            I => \N__14962\
        );

    \I__2718\ : Span4Mux_v
    port map (
            O => \N__14965\,
            I => \N__14959\
        );

    \I__2717\ : Span4Mux_v
    port map (
            O => \N__14962\,
            I => \N__14956\
        );

    \I__2716\ : Sp12to4
    port map (
            O => \N__14959\,
            I => \N__14953\
        );

    \I__2715\ : Span4Mux_h
    port map (
            O => \N__14956\,
            I => \N__14950\
        );

    \I__2714\ : Span12Mux_v
    port map (
            O => \N__14953\,
            I => \N__14947\
        );

    \I__2713\ : Span4Mux_h
    port map (
            O => \N__14950\,
            I => \N__14944\
        );

    \I__2712\ : Odrv12
    port map (
            O => \N__14947\,
            I => \line_buffer.n476\
        );

    \I__2711\ : Odrv4
    port map (
            O => \N__14944\,
            I => \line_buffer.n476\
        );

    \I__2710\ : CEMux
    port map (
            O => \N__14939\,
            I => \N__14936\
        );

    \I__2709\ : LocalMux
    port map (
            O => \N__14936\,
            I => \N__14933\
        );

    \I__2708\ : Span4Mux_h
    port map (
            O => \N__14933\,
            I => \N__14930\
        );

    \I__2707\ : Odrv4
    port map (
            O => \N__14930\,
            I => \receive_module.n3674\
        );

    \I__2706\ : InMux
    port map (
            O => \N__14927\,
            I => \N__14924\
        );

    \I__2705\ : LocalMux
    port map (
            O => \N__14924\,
            I => \N__14913\
        );

    \I__2704\ : InMux
    port map (
            O => \N__14923\,
            I => \N__14910\
        );

    \I__2703\ : InMux
    port map (
            O => \N__14922\,
            I => \N__14903\
        );

    \I__2702\ : InMux
    port map (
            O => \N__14921\,
            I => \N__14903\
        );

    \I__2701\ : InMux
    port map (
            O => \N__14920\,
            I => \N__14903\
        );

    \I__2700\ : InMux
    port map (
            O => \N__14919\,
            I => \N__14896\
        );

    \I__2699\ : InMux
    port map (
            O => \N__14918\,
            I => \N__14896\
        );

    \I__2698\ : InMux
    port map (
            O => \N__14917\,
            I => \N__14896\
        );

    \I__2697\ : InMux
    port map (
            O => \N__14916\,
            I => \N__14893\
        );

    \I__2696\ : Odrv4
    port map (
            O => \N__14913\,
            I => \RX_ADDR_11\
        );

    \I__2695\ : LocalMux
    port map (
            O => \N__14910\,
            I => \RX_ADDR_11\
        );

    \I__2694\ : LocalMux
    port map (
            O => \N__14903\,
            I => \RX_ADDR_11\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__14896\,
            I => \RX_ADDR_11\
        );

    \I__2692\ : LocalMux
    port map (
            O => \N__14893\,
            I => \RX_ADDR_11\
        );

    \I__2691\ : CascadeMux
    port map (
            O => \N__14882\,
            I => \N__14876\
        );

    \I__2690\ : InMux
    port map (
            O => \N__14881\,
            I => \N__14869\
        );

    \I__2689\ : InMux
    port map (
            O => \N__14880\,
            I => \N__14869\
        );

    \I__2688\ : InMux
    port map (
            O => \N__14879\,
            I => \N__14869\
        );

    \I__2687\ : InMux
    port map (
            O => \N__14876\,
            I => \N__14861\
        );

    \I__2686\ : LocalMux
    port map (
            O => \N__14869\,
            I => \N__14858\
        );

    \I__2685\ : InMux
    port map (
            O => \N__14868\,
            I => \N__14855\
        );

    \I__2684\ : InMux
    port map (
            O => \N__14867\,
            I => \N__14852\
        );

    \I__2683\ : InMux
    port map (
            O => \N__14866\,
            I => \N__14847\
        );

    \I__2682\ : InMux
    port map (
            O => \N__14865\,
            I => \N__14847\
        );

    \I__2681\ : InMux
    port map (
            O => \N__14864\,
            I => \N__14844\
        );

    \I__2680\ : LocalMux
    port map (
            O => \N__14861\,
            I => \N__14839\
        );

    \I__2679\ : Span4Mux_v
    port map (
            O => \N__14858\,
            I => \N__14839\
        );

    \I__2678\ : LocalMux
    port map (
            O => \N__14855\,
            I => \RX_ADDR_12\
        );

    \I__2677\ : LocalMux
    port map (
            O => \N__14852\,
            I => \RX_ADDR_12\
        );

    \I__2676\ : LocalMux
    port map (
            O => \N__14847\,
            I => \RX_ADDR_12\
        );

    \I__2675\ : LocalMux
    port map (
            O => \N__14844\,
            I => \RX_ADDR_12\
        );

    \I__2674\ : Odrv4
    port map (
            O => \N__14839\,
            I => \RX_ADDR_12\
        );

    \I__2673\ : InMux
    port map (
            O => \N__14828\,
            I => \N__14818\
        );

    \I__2672\ : CascadeMux
    port map (
            O => \N__14827\,
            I => \N__14814\
        );

    \I__2671\ : CascadeMux
    port map (
            O => \N__14826\,
            I => \N__14811\
        );

    \I__2670\ : CascadeMux
    port map (
            O => \N__14825\,
            I => \N__14808\
        );

    \I__2669\ : CascadeMux
    port map (
            O => \N__14824\,
            I => \N__14805\
        );

    \I__2668\ : CascadeMux
    port map (
            O => \N__14823\,
            I => \N__14802\
        );

    \I__2667\ : CascadeMux
    port map (
            O => \N__14822\,
            I => \N__14799\
        );

    \I__2666\ : CascadeMux
    port map (
            O => \N__14821\,
            I => \N__14796\
        );

    \I__2665\ : LocalMux
    port map (
            O => \N__14818\,
            I => \N__14793\
        );

    \I__2664\ : InMux
    port map (
            O => \N__14817\,
            I => \N__14790\
        );

    \I__2663\ : InMux
    port map (
            O => \N__14814\,
            I => \N__14787\
        );

    \I__2662\ : InMux
    port map (
            O => \N__14811\,
            I => \N__14784\
        );

    \I__2661\ : InMux
    port map (
            O => \N__14808\,
            I => \N__14781\
        );

    \I__2660\ : InMux
    port map (
            O => \N__14805\,
            I => \N__14776\
        );

    \I__2659\ : InMux
    port map (
            O => \N__14802\,
            I => \N__14776\
        );

    \I__2658\ : InMux
    port map (
            O => \N__14799\,
            I => \N__14771\
        );

    \I__2657\ : InMux
    port map (
            O => \N__14796\,
            I => \N__14771\
        );

    \I__2656\ : Span4Mux_v
    port map (
            O => \N__14793\,
            I => \N__14768\
        );

    \I__2655\ : LocalMux
    port map (
            O => \N__14790\,
            I => \RX_ADDR_13\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__14787\,
            I => \RX_ADDR_13\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__14784\,
            I => \RX_ADDR_13\
        );

    \I__2652\ : LocalMux
    port map (
            O => \N__14781\,
            I => \RX_ADDR_13\
        );

    \I__2651\ : LocalMux
    port map (
            O => \N__14776\,
            I => \RX_ADDR_13\
        );

    \I__2650\ : LocalMux
    port map (
            O => \N__14771\,
            I => \RX_ADDR_13\
        );

    \I__2649\ : Odrv4
    port map (
            O => \N__14768\,
            I => \RX_ADDR_13\
        );

    \I__2648\ : SRMux
    port map (
            O => \N__14753\,
            I => \N__14750\
        );

    \I__2647\ : LocalMux
    port map (
            O => \N__14750\,
            I => \N__14745\
        );

    \I__2646\ : SRMux
    port map (
            O => \N__14749\,
            I => \N__14742\
        );

    \I__2645\ : SRMux
    port map (
            O => \N__14748\,
            I => \N__14738\
        );

    \I__2644\ : Span4Mux_h
    port map (
            O => \N__14745\,
            I => \N__14735\
        );

    \I__2643\ : LocalMux
    port map (
            O => \N__14742\,
            I => \N__14732\
        );

    \I__2642\ : SRMux
    port map (
            O => \N__14741\,
            I => \N__14729\
        );

    \I__2641\ : LocalMux
    port map (
            O => \N__14738\,
            I => \N__14726\
        );

    \I__2640\ : Span4Mux_h
    port map (
            O => \N__14735\,
            I => \N__14723\
        );

    \I__2639\ : Span4Mux_h
    port map (
            O => \N__14732\,
            I => \N__14720\
        );

    \I__2638\ : LocalMux
    port map (
            O => \N__14729\,
            I => \N__14717\
        );

    \I__2637\ : Span4Mux_h
    port map (
            O => \N__14726\,
            I => \N__14714\
        );

    \I__2636\ : Span4Mux_v
    port map (
            O => \N__14723\,
            I => \N__14711\
        );

    \I__2635\ : Span4Mux_v
    port map (
            O => \N__14720\,
            I => \N__14706\
        );

    \I__2634\ : Span4Mux_h
    port map (
            O => \N__14717\,
            I => \N__14706\
        );

    \I__2633\ : Span4Mux_h
    port map (
            O => \N__14714\,
            I => \N__14703\
        );

    \I__2632\ : Span4Mux_v
    port map (
            O => \N__14711\,
            I => \N__14698\
        );

    \I__2631\ : Span4Mux_h
    port map (
            O => \N__14706\,
            I => \N__14698\
        );

    \I__2630\ : Odrv4
    port map (
            O => \N__14703\,
            I => \line_buffer.n574\
        );

    \I__2629\ : Odrv4
    port map (
            O => \N__14698\,
            I => \line_buffer.n574\
        );

    \I__2628\ : InMux
    port map (
            O => \N__14693\,
            I => \N__14690\
        );

    \I__2627\ : LocalMux
    port map (
            O => \N__14690\,
            I => \N__14687\
        );

    \I__2626\ : Span4Mux_v
    port map (
            O => \N__14687\,
            I => \N__14684\
        );

    \I__2625\ : Odrv4
    port map (
            O => \N__14684\,
            I => \tvp_vs_buffer.BUFFER_1_0\
        );

    \I__2624\ : InMux
    port map (
            O => \N__14681\,
            I => \N__14678\
        );

    \I__2623\ : LocalMux
    port map (
            O => \N__14678\,
            I => \tvp_vs_buffer.BUFFER_2_0\
        );

    \I__2622\ : InMux
    port map (
            O => \N__14675\,
            I => \N__14672\
        );

    \I__2621\ : LocalMux
    port map (
            O => \N__14672\,
            I => \N__14668\
        );

    \I__2620\ : CascadeMux
    port map (
            O => \N__14671\,
            I => \N__14665\
        );

    \I__2619\ : Span4Mux_h
    port map (
            O => \N__14668\,
            I => \N__14662\
        );

    \I__2618\ : InMux
    port map (
            O => \N__14665\,
            I => \N__14659\
        );

    \I__2617\ : Odrv4
    port map (
            O => \N__14662\,
            I => \transmit_module.X_DELTA_PATTERN_0\
        );

    \I__2616\ : LocalMux
    port map (
            O => \N__14659\,
            I => \transmit_module.X_DELTA_PATTERN_0\
        );

    \I__2615\ : InMux
    port map (
            O => \N__14654\,
            I => \receive_module.n3152\
        );

    \I__2614\ : InMux
    port map (
            O => \N__14651\,
            I => \receive_module.n3153\
        );

    \I__2613\ : InMux
    port map (
            O => \N__14648\,
            I => \receive_module.n3154\
        );

    \I__2612\ : InMux
    port map (
            O => \N__14645\,
            I => \receive_module.n3155\
        );

    \I__2611\ : InMux
    port map (
            O => \N__14642\,
            I => \bfn_15_12_0_\
        );

    \I__2610\ : InMux
    port map (
            O => \N__14639\,
            I => \receive_module.n3157\
        );

    \I__2609\ : InMux
    port map (
            O => \N__14636\,
            I => \receive_module.n3158\
        );

    \I__2608\ : InMux
    port map (
            O => \N__14633\,
            I => \receive_module.n3159\
        );

    \I__2607\ : InMux
    port map (
            O => \N__14630\,
            I => \receive_module.n3160\
        );

    \I__2606\ : InMux
    port map (
            O => \N__14627\,
            I => \N__14624\
        );

    \I__2605\ : LocalMux
    port map (
            O => \N__14624\,
            I => \transmit_module.X_DELTA_PATTERN_10\
        );

    \I__2604\ : InMux
    port map (
            O => \N__14621\,
            I => \N__14618\
        );

    \I__2603\ : LocalMux
    port map (
            O => \N__14618\,
            I => \transmit_module.X_DELTA_PATTERN_9\
        );

    \I__2602\ : InMux
    port map (
            O => \N__14615\,
            I => \N__14612\
        );

    \I__2601\ : LocalMux
    port map (
            O => \N__14612\,
            I => \transmit_module.X_DELTA_PATTERN_11\
        );

    \I__2600\ : InMux
    port map (
            O => \N__14609\,
            I => \N__14606\
        );

    \I__2599\ : LocalMux
    port map (
            O => \N__14606\,
            I => \N__14603\
        );

    \I__2598\ : Span4Mux_h
    port map (
            O => \N__14603\,
            I => \N__14600\
        );

    \I__2597\ : Odrv4
    port map (
            O => \N__14600\,
            I => \transmit_module.X_DELTA_PATTERN_13\
        );

    \I__2596\ : InMux
    port map (
            O => \N__14597\,
            I => \N__14594\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__14594\,
            I => \transmit_module.X_DELTA_PATTERN_12\
        );

    \I__2594\ : InMux
    port map (
            O => \N__14591\,
            I => \bfn_15_11_0_\
        );

    \I__2593\ : InMux
    port map (
            O => \N__14588\,
            I => \receive_module.n3149\
        );

    \I__2592\ : InMux
    port map (
            O => \N__14585\,
            I => \receive_module.n3150\
        );

    \I__2591\ : InMux
    port map (
            O => \N__14582\,
            I => \receive_module.n3151\
        );

    \I__2590\ : InMux
    port map (
            O => \N__14579\,
            I => \N__14575\
        );

    \I__2589\ : CascadeMux
    port map (
            O => \N__14578\,
            I => \N__14570\
        );

    \I__2588\ : LocalMux
    port map (
            O => \N__14575\,
            I => \N__14567\
        );

    \I__2587\ : InMux
    port map (
            O => \N__14574\,
            I => \N__14564\
        );

    \I__2586\ : InMux
    port map (
            O => \N__14573\,
            I => \N__14561\
        );

    \I__2585\ : InMux
    port map (
            O => \N__14570\,
            I => \N__14558\
        );

    \I__2584\ : Odrv4
    port map (
            O => \N__14567\,
            I => \transmit_module.TX_ADDR_10\
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__14564\,
            I => \transmit_module.TX_ADDR_10\
        );

    \I__2582\ : LocalMux
    port map (
            O => \N__14561\,
            I => \transmit_module.TX_ADDR_10\
        );

    \I__2581\ : LocalMux
    port map (
            O => \N__14558\,
            I => \transmit_module.TX_ADDR_10\
        );

    \I__2580\ : InMux
    port map (
            O => \N__14549\,
            I => \N__14546\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__14546\,
            I => \N__14543\
        );

    \I__2578\ : Odrv4
    port map (
            O => \N__14543\,
            I => \transmit_module.ADDR_Y_COMPONENT_10\
        );

    \I__2577\ : InMux
    port map (
            O => \N__14540\,
            I => \N__14536\
        );

    \I__2576\ : CascadeMux
    port map (
            O => \N__14539\,
            I => \N__14531\
        );

    \I__2575\ : LocalMux
    port map (
            O => \N__14536\,
            I => \N__14528\
        );

    \I__2574\ : InMux
    port map (
            O => \N__14535\,
            I => \N__14523\
        );

    \I__2573\ : InMux
    port map (
            O => \N__14534\,
            I => \N__14523\
        );

    \I__2572\ : InMux
    port map (
            O => \N__14531\,
            I => \N__14520\
        );

    \I__2571\ : Odrv4
    port map (
            O => \N__14528\,
            I => \transmit_module.TX_ADDR_8\
        );

    \I__2570\ : LocalMux
    port map (
            O => \N__14523\,
            I => \transmit_module.TX_ADDR_8\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__14520\,
            I => \transmit_module.TX_ADDR_8\
        );

    \I__2568\ : InMux
    port map (
            O => \N__14513\,
            I => \N__14510\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__14510\,
            I => \N__14507\
        );

    \I__2566\ : Odrv4
    port map (
            O => \N__14507\,
            I => \transmit_module.ADDR_Y_COMPONENT_8\
        );

    \I__2565\ : InMux
    port map (
            O => \N__14504\,
            I => \N__14499\
        );

    \I__2564\ : InMux
    port map (
            O => \N__14503\,
            I => \N__14496\
        );

    \I__2563\ : InMux
    port map (
            O => \N__14502\,
            I => \N__14493\
        );

    \I__2562\ : LocalMux
    port map (
            O => \N__14499\,
            I => \N__14489\
        );

    \I__2561\ : LocalMux
    port map (
            O => \N__14496\,
            I => \N__14486\
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__14493\,
            I => \N__14483\
        );

    \I__2559\ : InMux
    port map (
            O => \N__14492\,
            I => \N__14480\
        );

    \I__2558\ : Odrv12
    port map (
            O => \N__14489\,
            I => \transmit_module.TX_ADDR_1\
        );

    \I__2557\ : Odrv4
    port map (
            O => \N__14486\,
            I => \transmit_module.TX_ADDR_1\
        );

    \I__2556\ : Odrv4
    port map (
            O => \N__14483\,
            I => \transmit_module.TX_ADDR_1\
        );

    \I__2555\ : LocalMux
    port map (
            O => \N__14480\,
            I => \transmit_module.TX_ADDR_1\
        );

    \I__2554\ : InMux
    port map (
            O => \N__14471\,
            I => \N__14468\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__14468\,
            I => \transmit_module.ADDR_Y_COMPONENT_1\
        );

    \I__2552\ : InMux
    port map (
            O => \N__14465\,
            I => \N__14462\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__14462\,
            I => \N__14457\
        );

    \I__2550\ : InMux
    port map (
            O => \N__14461\,
            I => \N__14454\
        );

    \I__2549\ : InMux
    port map (
            O => \N__14460\,
            I => \N__14451\
        );

    \I__2548\ : Span12Mux_v
    port map (
            O => \N__14457\,
            I => \N__14443\
        );

    \I__2547\ : LocalMux
    port map (
            O => \N__14454\,
            I => \N__14443\
        );

    \I__2546\ : LocalMux
    port map (
            O => \N__14451\,
            I => \N__14443\
        );

    \I__2545\ : InMux
    port map (
            O => \N__14450\,
            I => \N__14440\
        );

    \I__2544\ : Odrv12
    port map (
            O => \N__14443\,
            I => \transmit_module.TX_ADDR_0\
        );

    \I__2543\ : LocalMux
    port map (
            O => \N__14440\,
            I => \transmit_module.TX_ADDR_0\
        );

    \I__2542\ : InMux
    port map (
            O => \N__14435\,
            I => \N__14432\
        );

    \I__2541\ : LocalMux
    port map (
            O => \N__14432\,
            I => \N__14429\
        );

    \I__2540\ : Odrv4
    port map (
            O => \N__14429\,
            I => \transmit_module.ADDR_Y_COMPONENT_0\
        );

    \I__2539\ : IoInMux
    port map (
            O => \N__14426\,
            I => \N__14423\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__14423\,
            I => \N__14420\
        );

    \I__2537\ : IoSpan4Mux
    port map (
            O => \N__14420\,
            I => \N__14417\
        );

    \I__2536\ : Span4Mux_s1_h
    port map (
            O => \N__14417\,
            I => \N__14414\
        );

    \I__2535\ : Sp12to4
    port map (
            O => \N__14414\,
            I => \N__14410\
        );

    \I__2534\ : InMux
    port map (
            O => \N__14413\,
            I => \N__14407\
        );

    \I__2533\ : Span12Mux_h
    port map (
            O => \N__14410\,
            I => \N__14402\
        );

    \I__2532\ : LocalMux
    port map (
            O => \N__14407\,
            I => \N__14402\
        );

    \I__2531\ : Odrv12
    port map (
            O => \N__14402\,
            I => \DEBUG_c_1_c\
        );

    \I__2530\ : IoInMux
    port map (
            O => \N__14399\,
            I => \N__14396\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__14396\,
            I => \N__14393\
        );

    \I__2528\ : IoSpan4Mux
    port map (
            O => \N__14393\,
            I => \N__14390\
        );

    \I__2527\ : Span4Mux_s0_h
    port map (
            O => \N__14390\,
            I => \N__14386\
        );

    \I__2526\ : InMux
    port map (
            O => \N__14389\,
            I => \N__14383\
        );

    \I__2525\ : Sp12to4
    port map (
            O => \N__14386\,
            I => \N__14380\
        );

    \I__2524\ : LocalMux
    port map (
            O => \N__14383\,
            I => \N__14377\
        );

    \I__2523\ : Span12Mux_s11_h
    port map (
            O => \N__14380\,
            I => \N__14374\
        );

    \I__2522\ : Span4Mux_h
    port map (
            O => \N__14377\,
            I => \N__14371\
        );

    \I__2521\ : Span12Mux_v
    port map (
            O => \N__14374\,
            I => \N__14368\
        );

    \I__2520\ : Span4Mux_v
    port map (
            O => \N__14371\,
            I => \N__14365\
        );

    \I__2519\ : Odrv12
    port map (
            O => \N__14368\,
            I => \DEBUG_c_6_c\
        );

    \I__2518\ : Odrv4
    port map (
            O => \N__14365\,
            I => \DEBUG_c_6_c\
        );

    \I__2517\ : InMux
    port map (
            O => \N__14360\,
            I => \N__14357\
        );

    \I__2516\ : LocalMux
    port map (
            O => \N__14357\,
            I => \N__14354\
        );

    \I__2515\ : Odrv4
    port map (
            O => \N__14354\,
            I => \tvp_vs_buffer.BUFFER_0_0\
        );

    \I__2514\ : InMux
    port map (
            O => \N__14351\,
            I => \N__14348\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__14348\,
            I => \tvp_video_buffer.BUFFER_0_6\
        );

    \I__2512\ : CascadeMux
    port map (
            O => \N__14345\,
            I => \N__14341\
        );

    \I__2511\ : InMux
    port map (
            O => \N__14344\,
            I => \N__14336\
        );

    \I__2510\ : InMux
    port map (
            O => \N__14341\,
            I => \N__14336\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__14336\,
            I => \N__14332\
        );

    \I__2508\ : InMux
    port map (
            O => \N__14335\,
            I => \N__14329\
        );

    \I__2507\ : Odrv4
    port map (
            O => \N__14332\,
            I => \TVP_HSYNC_buff\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__14329\,
            I => \TVP_HSYNC_buff\
        );

    \I__2505\ : InMux
    port map (
            O => \N__14324\,
            I => \N__14321\
        );

    \I__2504\ : LocalMux
    port map (
            O => \N__14321\,
            I => \N__14318\
        );

    \I__2503\ : Span4Mux_h
    port map (
            O => \N__14318\,
            I => \N__14315\
        );

    \I__2502\ : Odrv4
    port map (
            O => \N__14315\,
            I => \transmit_module.n138\
        );

    \I__2501\ : InMux
    port map (
            O => \N__14312\,
            I => \N__14309\
        );

    \I__2500\ : LocalMux
    port map (
            O => \N__14309\,
            I => \N__14306\
        );

    \I__2499\ : Span4Mux_h
    port map (
            O => \N__14306\,
            I => \N__14302\
        );

    \I__2498\ : InMux
    port map (
            O => \N__14305\,
            I => \N__14299\
        );

    \I__2497\ : Odrv4
    port map (
            O => \N__14302\,
            I => \transmit_module.video_signal_controller.n3382\
        );

    \I__2496\ : LocalMux
    port map (
            O => \N__14299\,
            I => \transmit_module.video_signal_controller.n3382\
        );

    \I__2495\ : InMux
    port map (
            O => \N__14294\,
            I => \N__14291\
        );

    \I__2494\ : LocalMux
    port map (
            O => \N__14291\,
            I => \transmit_module.video_signal_controller.n3017\
        );

    \I__2493\ : CascadeMux
    port map (
            O => \N__14288\,
            I => \N__14284\
        );

    \I__2492\ : CascadeMux
    port map (
            O => \N__14287\,
            I => \N__14281\
        );

    \I__2491\ : InMux
    port map (
            O => \N__14284\,
            I => \N__14278\
        );

    \I__2490\ : InMux
    port map (
            O => \N__14281\,
            I => \N__14274\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__14278\,
            I => \N__14270\
        );

    \I__2488\ : InMux
    port map (
            O => \N__14277\,
            I => \N__14266\
        );

    \I__2487\ : LocalMux
    port map (
            O => \N__14274\,
            I => \N__14263\
        );

    \I__2486\ : InMux
    port map (
            O => \N__14273\,
            I => \N__14260\
        );

    \I__2485\ : Span4Mux_h
    port map (
            O => \N__14270\,
            I => \N__14257\
        );

    \I__2484\ : InMux
    port map (
            O => \N__14269\,
            I => \N__14254\
        );

    \I__2483\ : LocalMux
    port map (
            O => \N__14266\,
            I => \N__14247\
        );

    \I__2482\ : Span4Mux_v
    port map (
            O => \N__14263\,
            I => \N__14247\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__14260\,
            I => \N__14247\
        );

    \I__2480\ : Odrv4
    port map (
            O => \N__14257\,
            I => \transmit_module.video_signal_controller.VGA_X_11\
        );

    \I__2479\ : LocalMux
    port map (
            O => \N__14254\,
            I => \transmit_module.video_signal_controller.VGA_X_11\
        );

    \I__2478\ : Odrv4
    port map (
            O => \N__14247\,
            I => \transmit_module.video_signal_controller.VGA_X_11\
        );

    \I__2477\ : InMux
    port map (
            O => \N__14240\,
            I => \N__14237\
        );

    \I__2476\ : LocalMux
    port map (
            O => \N__14237\,
            I => \transmit_module.video_signal_controller.n7_adj_624\
        );

    \I__2475\ : InMux
    port map (
            O => \N__14234\,
            I => \N__14231\
        );

    \I__2474\ : LocalMux
    port map (
            O => \N__14231\,
            I => \N__14228\
        );

    \I__2473\ : Odrv12
    port map (
            O => \N__14228\,
            I => \transmit_module.n132\
        );

    \I__2472\ : InMux
    port map (
            O => \N__14225\,
            I => \N__14222\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__14222\,
            I => \N__14219\
        );

    \I__2470\ : Odrv12
    port map (
            O => \N__14219\,
            I => \transmit_module.ADDR_Y_COMPONENT_9\
        );

    \I__2469\ : InMux
    port map (
            O => \N__14216\,
            I => \N__14213\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__14213\,
            I => \N__14207\
        );

    \I__2467\ : InMux
    port map (
            O => \N__14212\,
            I => \N__14204\
        );

    \I__2466\ : InMux
    port map (
            O => \N__14211\,
            I => \N__14201\
        );

    \I__2465\ : CascadeMux
    port map (
            O => \N__14210\,
            I => \N__14198\
        );

    \I__2464\ : Span4Mux_h
    port map (
            O => \N__14207\,
            I => \N__14195\
        );

    \I__2463\ : LocalMux
    port map (
            O => \N__14204\,
            I => \N__14190\
        );

    \I__2462\ : LocalMux
    port map (
            O => \N__14201\,
            I => \N__14190\
        );

    \I__2461\ : InMux
    port map (
            O => \N__14198\,
            I => \N__14187\
        );

    \I__2460\ : Odrv4
    port map (
            O => \N__14195\,
            I => \transmit_module.TX_ADDR_9\
        );

    \I__2459\ : Odrv4
    port map (
            O => \N__14190\,
            I => \transmit_module.TX_ADDR_9\
        );

    \I__2458\ : LocalMux
    port map (
            O => \N__14187\,
            I => \transmit_module.TX_ADDR_9\
        );

    \I__2457\ : InMux
    port map (
            O => \N__14180\,
            I => \N__14177\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__14177\,
            I => \N__14173\
        );

    \I__2455\ : InMux
    port map (
            O => \N__14176\,
            I => \N__14170\
        );

    \I__2454\ : Odrv4
    port map (
            O => \N__14173\,
            I => \transmit_module.n107\
        );

    \I__2453\ : LocalMux
    port map (
            O => \N__14170\,
            I => \transmit_module.n107\
        );

    \I__2452\ : InMux
    port map (
            O => \N__14165\,
            I => \N__14161\
        );

    \I__2451\ : InMux
    port map (
            O => \N__14164\,
            I => \N__14158\
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__14161\,
            I => \N__14155\
        );

    \I__2449\ : LocalMux
    port map (
            O => \N__14158\,
            I => \N__14152\
        );

    \I__2448\ : Span4Mux_h
    port map (
            O => \N__14155\,
            I => \N__14149\
        );

    \I__2447\ : Odrv4
    port map (
            O => \N__14152\,
            I => \transmit_module.n115\
        );

    \I__2446\ : Odrv4
    port map (
            O => \N__14149\,
            I => \transmit_module.n115\
        );

    \I__2445\ : InMux
    port map (
            O => \N__14144\,
            I => \N__14141\
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__14141\,
            I => \N__14138\
        );

    \I__2443\ : Span4Mux_v
    port map (
            O => \N__14138\,
            I => \N__14135\
        );

    \I__2442\ : Odrv4
    port map (
            O => \N__14135\,
            I => \transmit_module.n116\
        );

    \I__2441\ : CascadeMux
    port map (
            O => \N__14132\,
            I => \transmit_module.n116_cascade_\
        );

    \I__2440\ : InMux
    port map (
            O => \N__14129\,
            I => \N__14126\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__14126\,
            I => \N__14122\
        );

    \I__2438\ : InMux
    port map (
            O => \N__14125\,
            I => \N__14119\
        );

    \I__2437\ : Odrv12
    port map (
            O => \N__14122\,
            I => \transmit_module.n147\
        );

    \I__2436\ : LocalMux
    port map (
            O => \N__14119\,
            I => \transmit_module.n147\
        );

    \I__2435\ : CascadeMux
    port map (
            O => \N__14114\,
            I => \N__14110\
        );

    \I__2434\ : CascadeMux
    port map (
            O => \N__14113\,
            I => \N__14107\
        );

    \I__2433\ : CascadeBuf
    port map (
            O => \N__14110\,
            I => \N__14104\
        );

    \I__2432\ : CascadeBuf
    port map (
            O => \N__14107\,
            I => \N__14101\
        );

    \I__2431\ : CascadeMux
    port map (
            O => \N__14104\,
            I => \N__14098\
        );

    \I__2430\ : CascadeMux
    port map (
            O => \N__14101\,
            I => \N__14095\
        );

    \I__2429\ : CascadeBuf
    port map (
            O => \N__14098\,
            I => \N__14092\
        );

    \I__2428\ : CascadeBuf
    port map (
            O => \N__14095\,
            I => \N__14089\
        );

    \I__2427\ : CascadeMux
    port map (
            O => \N__14092\,
            I => \N__14086\
        );

    \I__2426\ : CascadeMux
    port map (
            O => \N__14089\,
            I => \N__14083\
        );

    \I__2425\ : CascadeBuf
    port map (
            O => \N__14086\,
            I => \N__14080\
        );

    \I__2424\ : CascadeBuf
    port map (
            O => \N__14083\,
            I => \N__14077\
        );

    \I__2423\ : CascadeMux
    port map (
            O => \N__14080\,
            I => \N__14074\
        );

    \I__2422\ : CascadeMux
    port map (
            O => \N__14077\,
            I => \N__14071\
        );

    \I__2421\ : CascadeBuf
    port map (
            O => \N__14074\,
            I => \N__14068\
        );

    \I__2420\ : CascadeBuf
    port map (
            O => \N__14071\,
            I => \N__14065\
        );

    \I__2419\ : CascadeMux
    port map (
            O => \N__14068\,
            I => \N__14062\
        );

    \I__2418\ : CascadeMux
    port map (
            O => \N__14065\,
            I => \N__14059\
        );

    \I__2417\ : CascadeBuf
    port map (
            O => \N__14062\,
            I => \N__14056\
        );

    \I__2416\ : CascadeBuf
    port map (
            O => \N__14059\,
            I => \N__14053\
        );

    \I__2415\ : CascadeMux
    port map (
            O => \N__14056\,
            I => \N__14050\
        );

    \I__2414\ : CascadeMux
    port map (
            O => \N__14053\,
            I => \N__14047\
        );

    \I__2413\ : CascadeBuf
    port map (
            O => \N__14050\,
            I => \N__14044\
        );

    \I__2412\ : CascadeBuf
    port map (
            O => \N__14047\,
            I => \N__14041\
        );

    \I__2411\ : CascadeMux
    port map (
            O => \N__14044\,
            I => \N__14038\
        );

    \I__2410\ : CascadeMux
    port map (
            O => \N__14041\,
            I => \N__14035\
        );

    \I__2409\ : CascadeBuf
    port map (
            O => \N__14038\,
            I => \N__14032\
        );

    \I__2408\ : CascadeBuf
    port map (
            O => \N__14035\,
            I => \N__14029\
        );

    \I__2407\ : CascadeMux
    port map (
            O => \N__14032\,
            I => \N__14026\
        );

    \I__2406\ : CascadeMux
    port map (
            O => \N__14029\,
            I => \N__14023\
        );

    \I__2405\ : CascadeBuf
    port map (
            O => \N__14026\,
            I => \N__14020\
        );

    \I__2404\ : CascadeBuf
    port map (
            O => \N__14023\,
            I => \N__14017\
        );

    \I__2403\ : CascadeMux
    port map (
            O => \N__14020\,
            I => \N__14014\
        );

    \I__2402\ : CascadeMux
    port map (
            O => \N__14017\,
            I => \N__14011\
        );

    \I__2401\ : CascadeBuf
    port map (
            O => \N__14014\,
            I => \N__14008\
        );

    \I__2400\ : CascadeBuf
    port map (
            O => \N__14011\,
            I => \N__14005\
        );

    \I__2399\ : CascadeMux
    port map (
            O => \N__14008\,
            I => \N__14002\
        );

    \I__2398\ : CascadeMux
    port map (
            O => \N__14005\,
            I => \N__13999\
        );

    \I__2397\ : CascadeBuf
    port map (
            O => \N__14002\,
            I => \N__13996\
        );

    \I__2396\ : CascadeBuf
    port map (
            O => \N__13999\,
            I => \N__13993\
        );

    \I__2395\ : CascadeMux
    port map (
            O => \N__13996\,
            I => \N__13990\
        );

    \I__2394\ : CascadeMux
    port map (
            O => \N__13993\,
            I => \N__13987\
        );

    \I__2393\ : CascadeBuf
    port map (
            O => \N__13990\,
            I => \N__13984\
        );

    \I__2392\ : CascadeBuf
    port map (
            O => \N__13987\,
            I => \N__13981\
        );

    \I__2391\ : CascadeMux
    port map (
            O => \N__13984\,
            I => \N__13978\
        );

    \I__2390\ : CascadeMux
    port map (
            O => \N__13981\,
            I => \N__13975\
        );

    \I__2389\ : CascadeBuf
    port map (
            O => \N__13978\,
            I => \N__13972\
        );

    \I__2388\ : CascadeBuf
    port map (
            O => \N__13975\,
            I => \N__13969\
        );

    \I__2387\ : CascadeMux
    port map (
            O => \N__13972\,
            I => \N__13966\
        );

    \I__2386\ : CascadeMux
    port map (
            O => \N__13969\,
            I => \N__13963\
        );

    \I__2385\ : CascadeBuf
    port map (
            O => \N__13966\,
            I => \N__13960\
        );

    \I__2384\ : CascadeBuf
    port map (
            O => \N__13963\,
            I => \N__13957\
        );

    \I__2383\ : CascadeMux
    port map (
            O => \N__13960\,
            I => \N__13954\
        );

    \I__2382\ : CascadeMux
    port map (
            O => \N__13957\,
            I => \N__13951\
        );

    \I__2381\ : CascadeBuf
    port map (
            O => \N__13954\,
            I => \N__13948\
        );

    \I__2380\ : CascadeBuf
    port map (
            O => \N__13951\,
            I => \N__13945\
        );

    \I__2379\ : CascadeMux
    port map (
            O => \N__13948\,
            I => \N__13942\
        );

    \I__2378\ : CascadeMux
    port map (
            O => \N__13945\,
            I => \N__13939\
        );

    \I__2377\ : CascadeBuf
    port map (
            O => \N__13942\,
            I => \N__13936\
        );

    \I__2376\ : CascadeBuf
    port map (
            O => \N__13939\,
            I => \N__13933\
        );

    \I__2375\ : CascadeMux
    port map (
            O => \N__13936\,
            I => \N__13930\
        );

    \I__2374\ : CascadeMux
    port map (
            O => \N__13933\,
            I => \N__13927\
        );

    \I__2373\ : InMux
    port map (
            O => \N__13930\,
            I => \N__13924\
        );

    \I__2372\ : InMux
    port map (
            O => \N__13927\,
            I => \N__13921\
        );

    \I__2371\ : LocalMux
    port map (
            O => \N__13924\,
            I => \N__13918\
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__13921\,
            I => \N__13915\
        );

    \I__2369\ : Span4Mux_h
    port map (
            O => \N__13918\,
            I => \N__13912\
        );

    \I__2368\ : Span12Mux_h
    port map (
            O => \N__13915\,
            I => \N__13909\
        );

    \I__2367\ : Sp12to4
    port map (
            O => \N__13912\,
            I => \N__13906\
        );

    \I__2366\ : Span12Mux_v
    port map (
            O => \N__13909\,
            I => \N__13903\
        );

    \I__2365\ : Span12Mux_v
    port map (
            O => \N__13906\,
            I => \N__13900\
        );

    \I__2364\ : Odrv12
    port map (
            O => \N__13903\,
            I => n28
        );

    \I__2363\ : Odrv12
    port map (
            O => \N__13900\,
            I => n28
        );

    \I__2362\ : InMux
    port map (
            O => \N__13895\,
            I => \N__13891\
        );

    \I__2361\ : InMux
    port map (
            O => \N__13894\,
            I => \N__13888\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__13891\,
            I => \transmit_module.n106\
        );

    \I__2359\ : LocalMux
    port map (
            O => \N__13888\,
            I => \transmit_module.n106\
        );

    \I__2358\ : InMux
    port map (
            O => \N__13883\,
            I => \N__13880\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__13880\,
            I => \N__13877\
        );

    \I__2356\ : Odrv4
    port map (
            O => \N__13877\,
            I => \transmit_module.n137\
        );

    \I__2355\ : CascadeMux
    port map (
            O => \N__13874\,
            I => \N__13871\
        );

    \I__2354\ : CascadeBuf
    port map (
            O => \N__13871\,
            I => \N__13867\
        );

    \I__2353\ : CascadeMux
    port map (
            O => \N__13870\,
            I => \N__13864\
        );

    \I__2352\ : CascadeMux
    port map (
            O => \N__13867\,
            I => \N__13861\
        );

    \I__2351\ : CascadeBuf
    port map (
            O => \N__13864\,
            I => \N__13858\
        );

    \I__2350\ : CascadeBuf
    port map (
            O => \N__13861\,
            I => \N__13855\
        );

    \I__2349\ : CascadeMux
    port map (
            O => \N__13858\,
            I => \N__13852\
        );

    \I__2348\ : CascadeMux
    port map (
            O => \N__13855\,
            I => \N__13849\
        );

    \I__2347\ : CascadeBuf
    port map (
            O => \N__13852\,
            I => \N__13846\
        );

    \I__2346\ : CascadeBuf
    port map (
            O => \N__13849\,
            I => \N__13843\
        );

    \I__2345\ : CascadeMux
    port map (
            O => \N__13846\,
            I => \N__13840\
        );

    \I__2344\ : CascadeMux
    port map (
            O => \N__13843\,
            I => \N__13837\
        );

    \I__2343\ : CascadeBuf
    port map (
            O => \N__13840\,
            I => \N__13834\
        );

    \I__2342\ : CascadeBuf
    port map (
            O => \N__13837\,
            I => \N__13831\
        );

    \I__2341\ : CascadeMux
    port map (
            O => \N__13834\,
            I => \N__13828\
        );

    \I__2340\ : CascadeMux
    port map (
            O => \N__13831\,
            I => \N__13825\
        );

    \I__2339\ : CascadeBuf
    port map (
            O => \N__13828\,
            I => \N__13822\
        );

    \I__2338\ : CascadeBuf
    port map (
            O => \N__13825\,
            I => \N__13819\
        );

    \I__2337\ : CascadeMux
    port map (
            O => \N__13822\,
            I => \N__13816\
        );

    \I__2336\ : CascadeMux
    port map (
            O => \N__13819\,
            I => \N__13813\
        );

    \I__2335\ : CascadeBuf
    port map (
            O => \N__13816\,
            I => \N__13810\
        );

    \I__2334\ : CascadeBuf
    port map (
            O => \N__13813\,
            I => \N__13807\
        );

    \I__2333\ : CascadeMux
    port map (
            O => \N__13810\,
            I => \N__13804\
        );

    \I__2332\ : CascadeMux
    port map (
            O => \N__13807\,
            I => \N__13801\
        );

    \I__2331\ : CascadeBuf
    port map (
            O => \N__13804\,
            I => \N__13798\
        );

    \I__2330\ : CascadeBuf
    port map (
            O => \N__13801\,
            I => \N__13795\
        );

    \I__2329\ : CascadeMux
    port map (
            O => \N__13798\,
            I => \N__13792\
        );

    \I__2328\ : CascadeMux
    port map (
            O => \N__13795\,
            I => \N__13789\
        );

    \I__2327\ : CascadeBuf
    port map (
            O => \N__13792\,
            I => \N__13786\
        );

    \I__2326\ : CascadeBuf
    port map (
            O => \N__13789\,
            I => \N__13783\
        );

    \I__2325\ : CascadeMux
    port map (
            O => \N__13786\,
            I => \N__13780\
        );

    \I__2324\ : CascadeMux
    port map (
            O => \N__13783\,
            I => \N__13777\
        );

    \I__2323\ : CascadeBuf
    port map (
            O => \N__13780\,
            I => \N__13774\
        );

    \I__2322\ : CascadeBuf
    port map (
            O => \N__13777\,
            I => \N__13771\
        );

    \I__2321\ : CascadeMux
    port map (
            O => \N__13774\,
            I => \N__13768\
        );

    \I__2320\ : CascadeMux
    port map (
            O => \N__13771\,
            I => \N__13765\
        );

    \I__2319\ : CascadeBuf
    port map (
            O => \N__13768\,
            I => \N__13762\
        );

    \I__2318\ : CascadeBuf
    port map (
            O => \N__13765\,
            I => \N__13759\
        );

    \I__2317\ : CascadeMux
    port map (
            O => \N__13762\,
            I => \N__13756\
        );

    \I__2316\ : CascadeMux
    port map (
            O => \N__13759\,
            I => \N__13753\
        );

    \I__2315\ : CascadeBuf
    port map (
            O => \N__13756\,
            I => \N__13750\
        );

    \I__2314\ : CascadeBuf
    port map (
            O => \N__13753\,
            I => \N__13747\
        );

    \I__2313\ : CascadeMux
    port map (
            O => \N__13750\,
            I => \N__13744\
        );

    \I__2312\ : CascadeMux
    port map (
            O => \N__13747\,
            I => \N__13741\
        );

    \I__2311\ : CascadeBuf
    port map (
            O => \N__13744\,
            I => \N__13738\
        );

    \I__2310\ : CascadeBuf
    port map (
            O => \N__13741\,
            I => \N__13735\
        );

    \I__2309\ : CascadeMux
    port map (
            O => \N__13738\,
            I => \N__13732\
        );

    \I__2308\ : CascadeMux
    port map (
            O => \N__13735\,
            I => \N__13729\
        );

    \I__2307\ : CascadeBuf
    port map (
            O => \N__13732\,
            I => \N__13726\
        );

    \I__2306\ : CascadeBuf
    port map (
            O => \N__13729\,
            I => \N__13723\
        );

    \I__2305\ : CascadeMux
    port map (
            O => \N__13726\,
            I => \N__13720\
        );

    \I__2304\ : CascadeMux
    port map (
            O => \N__13723\,
            I => \N__13717\
        );

    \I__2303\ : CascadeBuf
    port map (
            O => \N__13720\,
            I => \N__13714\
        );

    \I__2302\ : CascadeBuf
    port map (
            O => \N__13717\,
            I => \N__13711\
        );

    \I__2301\ : CascadeMux
    port map (
            O => \N__13714\,
            I => \N__13708\
        );

    \I__2300\ : CascadeMux
    port map (
            O => \N__13711\,
            I => \N__13705\
        );

    \I__2299\ : CascadeBuf
    port map (
            O => \N__13708\,
            I => \N__13702\
        );

    \I__2298\ : CascadeBuf
    port map (
            O => \N__13705\,
            I => \N__13699\
        );

    \I__2297\ : CascadeMux
    port map (
            O => \N__13702\,
            I => \N__13696\
        );

    \I__2296\ : CascadeMux
    port map (
            O => \N__13699\,
            I => \N__13693\
        );

    \I__2295\ : CascadeBuf
    port map (
            O => \N__13696\,
            I => \N__13690\
        );

    \I__2294\ : InMux
    port map (
            O => \N__13693\,
            I => \N__13687\
        );

    \I__2293\ : CascadeMux
    port map (
            O => \N__13690\,
            I => \N__13684\
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__13687\,
            I => \N__13681\
        );

    \I__2291\ : InMux
    port map (
            O => \N__13684\,
            I => \N__13678\
        );

    \I__2290\ : Span4Mux_h
    port map (
            O => \N__13681\,
            I => \N__13675\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__13678\,
            I => \N__13672\
        );

    \I__2288\ : Sp12to4
    port map (
            O => \N__13675\,
            I => \N__13669\
        );

    \I__2287\ : Sp12to4
    port map (
            O => \N__13672\,
            I => \N__13666\
        );

    \I__2286\ : Span12Mux_h
    port map (
            O => \N__13669\,
            I => \N__13661\
        );

    \I__2285\ : Span12Mux_s9_h
    port map (
            O => \N__13666\,
            I => \N__13661\
        );

    \I__2284\ : Span12Mux_v
    port map (
            O => \N__13661\,
            I => \N__13658\
        );

    \I__2283\ : Odrv12
    port map (
            O => \N__13658\,
            I => n18
        );

    \I__2282\ : InMux
    port map (
            O => \N__13655\,
            I => \N__13652\
        );

    \I__2281\ : LocalMux
    port map (
            O => \N__13652\,
            I => \N__13649\
        );

    \I__2280\ : Odrv4
    port map (
            O => \N__13649\,
            I => \transmit_module.n121\
        );

    \I__2279\ : InMux
    port map (
            O => \N__13646\,
            I => \transmit_module.n3172\
        );

    \I__2278\ : InMux
    port map (
            O => \N__13643\,
            I => \N__13640\
        );

    \I__2277\ : LocalMux
    port map (
            O => \N__13640\,
            I => \N__13637\
        );

    \I__2276\ : Odrv4
    port map (
            O => \N__13637\,
            I => \transmit_module.n120\
        );

    \I__2275\ : InMux
    port map (
            O => \N__13634\,
            I => \transmit_module.n3173\
        );

    \I__2274\ : InMux
    port map (
            O => \N__13631\,
            I => \transmit_module.n3174\
        );

    \I__2273\ : InMux
    port map (
            O => \N__13628\,
            I => \N__13625\
        );

    \I__2272\ : LocalMux
    port map (
            O => \N__13625\,
            I => \N__13622\
        );

    \I__2271\ : Span4Mux_h
    port map (
            O => \N__13622\,
            I => \N__13619\
        );

    \I__2270\ : Odrv4
    port map (
            O => \N__13619\,
            I => \transmit_module.n119\
        );

    \I__2269\ : InMux
    port map (
            O => \N__13616\,
            I => \N__13612\
        );

    \I__2268\ : InMux
    port map (
            O => \N__13615\,
            I => \N__13609\
        );

    \I__2267\ : LocalMux
    port map (
            O => \N__13612\,
            I => \transmit_module.n112\
        );

    \I__2266\ : LocalMux
    port map (
            O => \N__13609\,
            I => \transmit_module.n112\
        );

    \I__2265\ : InMux
    port map (
            O => \N__13604\,
            I => \N__13601\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__13601\,
            I => \N__13597\
        );

    \I__2263\ : InMux
    port map (
            O => \N__13600\,
            I => \N__13594\
        );

    \I__2262\ : Span4Mux_h
    port map (
            O => \N__13597\,
            I => \N__13591\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__13594\,
            I => \transmit_module.n146\
        );

    \I__2260\ : Odrv4
    port map (
            O => \N__13591\,
            I => \transmit_module.n146\
        );

    \I__2259\ : InMux
    port map (
            O => \N__13586\,
            I => \N__13583\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__13583\,
            I => \N__13580\
        );

    \I__2257\ : Odrv12
    port map (
            O => \N__13580\,
            I => \sync_buffer.BUFFER_1_0\
        );

    \I__2256\ : InMux
    port map (
            O => \N__13577\,
            I => \N__13574\
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__13574\,
            I => \N__13571\
        );

    \I__2254\ : Odrv4
    port map (
            O => \N__13571\,
            I => \RX_TX_SYNC_BUFF\
        );

    \I__2253\ : InMux
    port map (
            O => \N__13568\,
            I => \N__13565\
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__13565\,
            I => \transmit_module.n122\
        );

    \I__2251\ : CascadeMux
    port map (
            O => \N__13562\,
            I => \transmit_module.n137_cascade_\
        );

    \I__2250\ : InMux
    port map (
            O => \N__13559\,
            I => \transmit_module.n3163\
        );

    \I__2249\ : InMux
    port map (
            O => \N__13556\,
            I => \transmit_module.n3164\
        );

    \I__2248\ : CascadeMux
    port map (
            O => \N__13553\,
            I => \N__13550\
        );

    \I__2247\ : InMux
    port map (
            O => \N__13550\,
            I => \N__13547\
        );

    \I__2246\ : LocalMux
    port map (
            O => \N__13547\,
            I => \N__13544\
        );

    \I__2245\ : Odrv4
    port map (
            O => \N__13544\,
            I => \transmit_module.n128\
        );

    \I__2244\ : InMux
    port map (
            O => \N__13541\,
            I => \transmit_module.n3165\
        );

    \I__2243\ : InMux
    port map (
            O => \N__13538\,
            I => \N__13535\
        );

    \I__2242\ : LocalMux
    port map (
            O => \N__13535\,
            I => \N__13529\
        );

    \I__2241\ : InMux
    port map (
            O => \N__13534\,
            I => \N__13526\
        );

    \I__2240\ : InMux
    port map (
            O => \N__13533\,
            I => \N__13523\
        );

    \I__2239\ : InMux
    port map (
            O => \N__13532\,
            I => \N__13520\
        );

    \I__2238\ : Odrv4
    port map (
            O => \N__13529\,
            I => \transmit_module.TX_ADDR_5\
        );

    \I__2237\ : LocalMux
    port map (
            O => \N__13526\,
            I => \transmit_module.TX_ADDR_5\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__13523\,
            I => \transmit_module.TX_ADDR_5\
        );

    \I__2235\ : LocalMux
    port map (
            O => \N__13520\,
            I => \transmit_module.TX_ADDR_5\
        );

    \I__2234\ : CascadeMux
    port map (
            O => \N__13511\,
            I => \N__13508\
        );

    \I__2233\ : InMux
    port map (
            O => \N__13508\,
            I => \N__13505\
        );

    \I__2232\ : LocalMux
    port map (
            O => \N__13505\,
            I => \transmit_module.n127\
        );

    \I__2231\ : InMux
    port map (
            O => \N__13502\,
            I => \transmit_module.n3166\
        );

    \I__2230\ : InMux
    port map (
            O => \N__13499\,
            I => \N__13496\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__13496\,
            I => \transmit_module.n126\
        );

    \I__2228\ : InMux
    port map (
            O => \N__13493\,
            I => \transmit_module.n3167\
        );

    \I__2227\ : InMux
    port map (
            O => \N__13490\,
            I => \N__13487\
        );

    \I__2226\ : LocalMux
    port map (
            O => \N__13487\,
            I => \N__13483\
        );

    \I__2225\ : CascadeMux
    port map (
            O => \N__13486\,
            I => \N__13479\
        );

    \I__2224\ : Span4Mux_v
    port map (
            O => \N__13483\,
            I => \N__13475\
        );

    \I__2223\ : InMux
    port map (
            O => \N__13482\,
            I => \N__13472\
        );

    \I__2222\ : InMux
    port map (
            O => \N__13479\,
            I => \N__13469\
        );

    \I__2221\ : InMux
    port map (
            O => \N__13478\,
            I => \N__13466\
        );

    \I__2220\ : Odrv4
    port map (
            O => \N__13475\,
            I => \transmit_module.TX_ADDR_7\
        );

    \I__2219\ : LocalMux
    port map (
            O => \N__13472\,
            I => \transmit_module.TX_ADDR_7\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__13469\,
            I => \transmit_module.TX_ADDR_7\
        );

    \I__2217\ : LocalMux
    port map (
            O => \N__13466\,
            I => \transmit_module.TX_ADDR_7\
        );

    \I__2216\ : InMux
    port map (
            O => \N__13457\,
            I => \N__13454\
        );

    \I__2215\ : LocalMux
    port map (
            O => \N__13454\,
            I => \transmit_module.n125\
        );

    \I__2214\ : InMux
    port map (
            O => \N__13451\,
            I => \transmit_module.n3168\
        );

    \I__2213\ : InMux
    port map (
            O => \N__13448\,
            I => \N__13445\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__13445\,
            I => \N__13442\
        );

    \I__2211\ : Odrv4
    port map (
            O => \N__13442\,
            I => \transmit_module.n124\
        );

    \I__2210\ : InMux
    port map (
            O => \N__13439\,
            I => \bfn_14_16_0_\
        );

    \I__2209\ : InMux
    port map (
            O => \N__13436\,
            I => \N__13433\
        );

    \I__2208\ : LocalMux
    port map (
            O => \N__13433\,
            I => \N__13430\
        );

    \I__2207\ : Span4Mux_v
    port map (
            O => \N__13430\,
            I => \N__13427\
        );

    \I__2206\ : Odrv4
    port map (
            O => \N__13427\,
            I => \transmit_module.n123\
        );

    \I__2205\ : InMux
    port map (
            O => \N__13424\,
            I => \transmit_module.n3170\
        );

    \I__2204\ : InMux
    port map (
            O => \N__13421\,
            I => \transmit_module.n3171\
        );

    \I__2203\ : SRMux
    port map (
            O => \N__13418\,
            I => \N__13415\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__13415\,
            I => \N__13410\
        );

    \I__2201\ : SRMux
    port map (
            O => \N__13414\,
            I => \N__13407\
        );

    \I__2200\ : SRMux
    port map (
            O => \N__13413\,
            I => \N__13404\
        );

    \I__2199\ : Span4Mux_s2_v
    port map (
            O => \N__13410\,
            I => \N__13396\
        );

    \I__2198\ : LocalMux
    port map (
            O => \N__13407\,
            I => \N__13396\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__13404\,
            I => \N__13396\
        );

    \I__2196\ : SRMux
    port map (
            O => \N__13403\,
            I => \N__13393\
        );

    \I__2195\ : Span4Mux_v
    port map (
            O => \N__13396\,
            I => \N__13390\
        );

    \I__2194\ : LocalMux
    port map (
            O => \N__13393\,
            I => \N__13387\
        );

    \I__2193\ : Sp12to4
    port map (
            O => \N__13390\,
            I => \N__13384\
        );

    \I__2192\ : Span4Mux_h
    port map (
            O => \N__13387\,
            I => \N__13381\
        );

    \I__2191\ : Span12Mux_v
    port map (
            O => \N__13384\,
            I => \N__13378\
        );

    \I__2190\ : Span4Mux_h
    port map (
            O => \N__13381\,
            I => \N__13375\
        );

    \I__2189\ : Odrv12
    port map (
            O => \N__13378\,
            I => \line_buffer.n605\
        );

    \I__2188\ : Odrv4
    port map (
            O => \N__13375\,
            I => \line_buffer.n605\
        );

    \I__2187\ : InMux
    port map (
            O => \N__13370\,
            I => \N__13367\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__13367\,
            I => \N__13364\
        );

    \I__2185\ : Span4Mux_h
    port map (
            O => \N__13364\,
            I => \N__13361\
        );

    \I__2184\ : Span4Mux_h
    port map (
            O => \N__13361\,
            I => \N__13358\
        );

    \I__2183\ : Span4Mux_v
    port map (
            O => \N__13358\,
            I => \N__13355\
        );

    \I__2182\ : Odrv4
    port map (
            O => \N__13355\,
            I => \line_buffer.n568\
        );

    \I__2181\ : InMux
    port map (
            O => \N__13352\,
            I => \N__13349\
        );

    \I__2180\ : LocalMux
    port map (
            O => \N__13349\,
            I => \N__13346\
        );

    \I__2179\ : Span4Mux_h
    port map (
            O => \N__13346\,
            I => \N__13343\
        );

    \I__2178\ : Span4Mux_h
    port map (
            O => \N__13343\,
            I => \N__13340\
        );

    \I__2177\ : Odrv4
    port map (
            O => \N__13340\,
            I => \line_buffer.n560\
        );

    \I__2176\ : InMux
    port map (
            O => \N__13337\,
            I => \N__13334\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__13334\,
            I => \sync_buffer.BUFFER_0_0\
        );

    \I__2174\ : InMux
    port map (
            O => \N__13331\,
            I => \N__13328\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__13328\,
            I => \N__13325\
        );

    \I__2172\ : Odrv4
    port map (
            O => \N__13325\,
            I => \transmit_module.ADDR_Y_COMPONENT_6\
        );

    \I__2171\ : InMux
    port map (
            O => \N__13322\,
            I => \N__13319\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__13319\,
            I => \transmit_module.n131\
        );

    \I__2169\ : InMux
    port map (
            O => \N__13316\,
            I => \transmit_module.n3162\
        );

    \I__2168\ : CascadeMux
    port map (
            O => \N__13313\,
            I => \receive_module.rx_counter.n5_cascade_\
        );

    \I__2167\ : InMux
    port map (
            O => \N__13310\,
            I => \N__13306\
        );

    \I__2166\ : InMux
    port map (
            O => \N__13309\,
            I => \N__13301\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__13306\,
            I => \N__13298\
        );

    \I__2164\ : InMux
    port map (
            O => \N__13305\,
            I => \N__13293\
        );

    \I__2163\ : InMux
    port map (
            O => \N__13304\,
            I => \N__13293\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__13301\,
            I => \receive_module.rx_counter.Y_7\
        );

    \I__2161\ : Odrv4
    port map (
            O => \N__13298\,
            I => \receive_module.rx_counter.Y_7\
        );

    \I__2160\ : LocalMux
    port map (
            O => \N__13293\,
            I => \receive_module.rx_counter.Y_7\
        );

    \I__2159\ : CascadeMux
    port map (
            O => \N__13286\,
            I => \receive_module.rx_counter.n3455_cascade_\
        );

    \I__2158\ : InMux
    port map (
            O => \N__13283\,
            I => \N__13280\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__13280\,
            I => \N__13276\
        );

    \I__2156\ : InMux
    port map (
            O => \N__13279\,
            I => \N__13273\
        );

    \I__2155\ : Odrv4
    port map (
            O => \N__13276\,
            I => \receive_module.rx_counter.n3680\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__13273\,
            I => \receive_module.rx_counter.n3680\
        );

    \I__2153\ : CascadeMux
    port map (
            O => \N__13268\,
            I => \N__13265\
        );

    \I__2152\ : InMux
    port map (
            O => \N__13265\,
            I => \N__13259\
        );

    \I__2151\ : InMux
    port map (
            O => \N__13264\,
            I => \N__13256\
        );

    \I__2150\ : InMux
    port map (
            O => \N__13263\,
            I => \N__13253\
        );

    \I__2149\ : InMux
    port map (
            O => \N__13262\,
            I => \N__13250\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__13259\,
            I => \N__13247\
        );

    \I__2147\ : LocalMux
    port map (
            O => \N__13256\,
            I => \receive_module.rx_counter.Y_8\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__13253\,
            I => \receive_module.rx_counter.Y_8\
        );

    \I__2145\ : LocalMux
    port map (
            O => \N__13250\,
            I => \receive_module.rx_counter.Y_8\
        );

    \I__2144\ : Odrv4
    port map (
            O => \N__13247\,
            I => \receive_module.rx_counter.Y_8\
        );

    \I__2143\ : InMux
    port map (
            O => \N__13238\,
            I => \N__13235\
        );

    \I__2142\ : LocalMux
    port map (
            O => \N__13235\,
            I => \receive_module.rx_counter.n3481\
        );

    \I__2141\ : CascadeMux
    port map (
            O => \N__13232\,
            I => \receive_module.rx_counter.n4_adj_612_cascade_\
        );

    \I__2140\ : InMux
    port map (
            O => \N__13229\,
            I => \N__13226\
        );

    \I__2139\ : LocalMux
    port map (
            O => \N__13226\,
            I => \receive_module.rx_counter.n54\
        );

    \I__2138\ : InMux
    port map (
            O => \N__13223\,
            I => \N__13220\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__13220\,
            I => \N__13214\
        );

    \I__2136\ : InMux
    port map (
            O => \N__13219\,
            I => \N__13211\
        );

    \I__2135\ : InMux
    port map (
            O => \N__13218\,
            I => \N__13206\
        );

    \I__2134\ : InMux
    port map (
            O => \N__13217\,
            I => \N__13206\
        );

    \I__2133\ : Odrv4
    port map (
            O => \N__13214\,
            I => \receive_module.rx_counter.Y_1\
        );

    \I__2132\ : LocalMux
    port map (
            O => \N__13211\,
            I => \receive_module.rx_counter.Y_1\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__13206\,
            I => \receive_module.rx_counter.Y_1\
        );

    \I__2130\ : InMux
    port map (
            O => \N__13199\,
            I => \N__13195\
        );

    \I__2129\ : CascadeMux
    port map (
            O => \N__13198\,
            I => \N__13190\
        );

    \I__2128\ : LocalMux
    port map (
            O => \N__13195\,
            I => \N__13187\
        );

    \I__2127\ : InMux
    port map (
            O => \N__13194\,
            I => \N__13184\
        );

    \I__2126\ : InMux
    port map (
            O => \N__13193\,
            I => \N__13181\
        );

    \I__2125\ : InMux
    port map (
            O => \N__13190\,
            I => \N__13178\
        );

    \I__2124\ : Odrv4
    port map (
            O => \N__13187\,
            I => \receive_module.rx_counter.Y_0\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__13184\,
            I => \receive_module.rx_counter.Y_0\
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__13181\,
            I => \receive_module.rx_counter.Y_0\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__13178\,
            I => \receive_module.rx_counter.Y_0\
        );

    \I__2120\ : InMux
    port map (
            O => \N__13169\,
            I => \N__13166\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__13166\,
            I => \N__13160\
        );

    \I__2118\ : InMux
    port map (
            O => \N__13165\,
            I => \N__13157\
        );

    \I__2117\ : InMux
    port map (
            O => \N__13164\,
            I => \N__13152\
        );

    \I__2116\ : InMux
    port map (
            O => \N__13163\,
            I => \N__13152\
        );

    \I__2115\ : Odrv4
    port map (
            O => \N__13160\,
            I => \receive_module.rx_counter.Y_2\
        );

    \I__2114\ : LocalMux
    port map (
            O => \N__13157\,
            I => \receive_module.rx_counter.Y_2\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__13152\,
            I => \receive_module.rx_counter.Y_2\
        );

    \I__2112\ : InMux
    port map (
            O => \N__13145\,
            I => \N__13142\
        );

    \I__2111\ : LocalMux
    port map (
            O => \N__13142\,
            I => \receive_module.rx_counter.n3453\
        );

    \I__2110\ : InMux
    port map (
            O => \N__13139\,
            I => \N__13136\
        );

    \I__2109\ : LocalMux
    port map (
            O => \N__13136\,
            I => \N__13130\
        );

    \I__2108\ : InMux
    port map (
            O => \N__13135\,
            I => \N__13127\
        );

    \I__2107\ : InMux
    port map (
            O => \N__13134\,
            I => \N__13122\
        );

    \I__2106\ : InMux
    port map (
            O => \N__13133\,
            I => \N__13122\
        );

    \I__2105\ : Odrv4
    port map (
            O => \N__13130\,
            I => \receive_module.rx_counter.Y_3\
        );

    \I__2104\ : LocalMux
    port map (
            O => \N__13127\,
            I => \receive_module.rx_counter.Y_3\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__13122\,
            I => \receive_module.rx_counter.Y_3\
        );

    \I__2102\ : InMux
    port map (
            O => \N__13115\,
            I => \N__13111\
        );

    \I__2101\ : InMux
    port map (
            O => \N__13114\,
            I => \N__13106\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__13111\,
            I => \N__13103\
        );

    \I__2099\ : InMux
    port map (
            O => \N__13110\,
            I => \N__13100\
        );

    \I__2098\ : InMux
    port map (
            O => \N__13109\,
            I => \N__13097\
        );

    \I__2097\ : LocalMux
    port map (
            O => \N__13106\,
            I => \receive_module.rx_counter.Y_4\
        );

    \I__2096\ : Odrv4
    port map (
            O => \N__13103\,
            I => \receive_module.rx_counter.Y_4\
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__13100\,
            I => \receive_module.rx_counter.Y_4\
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__13097\,
            I => \receive_module.rx_counter.Y_4\
        );

    \I__2093\ : InMux
    port map (
            O => \N__13088\,
            I => \N__13085\
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__13085\,
            I => \receive_module.rx_counter.n4\
        );

    \I__2091\ : InMux
    port map (
            O => \N__13082\,
            I => \N__13079\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__13079\,
            I => \RX_TX_SYNC\
        );

    \I__2089\ : SRMux
    port map (
            O => \N__13076\,
            I => \N__13073\
        );

    \I__2088\ : LocalMux
    port map (
            O => \N__13073\,
            I => \N__13068\
        );

    \I__2087\ : SRMux
    port map (
            O => \N__13072\,
            I => \N__13065\
        );

    \I__2086\ : SRMux
    port map (
            O => \N__13071\,
            I => \N__13062\
        );

    \I__2085\ : Span4Mux_v
    port map (
            O => \N__13068\,
            I => \N__13054\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__13065\,
            I => \N__13054\
        );

    \I__2083\ : LocalMux
    port map (
            O => \N__13062\,
            I => \N__13054\
        );

    \I__2082\ : SRMux
    port map (
            O => \N__13061\,
            I => \N__13051\
        );

    \I__2081\ : Span4Mux_v
    port map (
            O => \N__13054\,
            I => \N__13048\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__13051\,
            I => \N__13045\
        );

    \I__2079\ : Span4Mux_h
    port map (
            O => \N__13048\,
            I => \N__13040\
        );

    \I__2078\ : Span4Mux_h
    port map (
            O => \N__13045\,
            I => \N__13040\
        );

    \I__2077\ : Span4Mux_h
    port map (
            O => \N__13040\,
            I => \N__13037\
        );

    \I__2076\ : Span4Mux_h
    port map (
            O => \N__13037\,
            I => \N__13034\
        );

    \I__2075\ : Span4Mux_v
    port map (
            O => \N__13034\,
            I => \N__13031\
        );

    \I__2074\ : Odrv4
    port map (
            O => \N__13031\,
            I => \line_buffer.n477\
        );

    \I__2073\ : SRMux
    port map (
            O => \N__13028\,
            I => \N__13025\
        );

    \I__2072\ : LocalMux
    port map (
            O => \N__13025\,
            I => \N__13021\
        );

    \I__2071\ : SRMux
    port map (
            O => \N__13024\,
            I => \N__13018\
        );

    \I__2070\ : Span4Mux_v
    port map (
            O => \N__13021\,
            I => \N__13011\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__13018\,
            I => \N__13011\
        );

    \I__2068\ : SRMux
    port map (
            O => \N__13017\,
            I => \N__13008\
        );

    \I__2067\ : SRMux
    port map (
            O => \N__13016\,
            I => \N__13005\
        );

    \I__2066\ : Span4Mux_v
    port map (
            O => \N__13011\,
            I => \N__12998\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__13008\,
            I => \N__12998\
        );

    \I__2064\ : LocalMux
    port map (
            O => \N__13005\,
            I => \N__12998\
        );

    \I__2063\ : Span4Mux_v
    port map (
            O => \N__12998\,
            I => \N__12995\
        );

    \I__2062\ : Sp12to4
    port map (
            O => \N__12995\,
            I => \N__12992\
        );

    \I__2061\ : Odrv12
    port map (
            O => \N__12992\,
            I => \line_buffer.n541\
        );

    \I__2060\ : InMux
    port map (
            O => \N__12989\,
            I => \N__12984\
        );

    \I__2059\ : InMux
    port map (
            O => \N__12988\,
            I => \N__12981\
        );

    \I__2058\ : InMux
    port map (
            O => \N__12987\,
            I => \N__12978\
        );

    \I__2057\ : LocalMux
    port map (
            O => \N__12984\,
            I => \receive_module.rx_counter.X_3\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__12981\,
            I => \receive_module.rx_counter.X_3\
        );

    \I__2055\ : LocalMux
    port map (
            O => \N__12978\,
            I => \receive_module.rx_counter.X_3\
        );

    \I__2054\ : InMux
    port map (
            O => \N__12971\,
            I => \N__12966\
        );

    \I__2053\ : InMux
    port map (
            O => \N__12970\,
            I => \N__12963\
        );

    \I__2052\ : InMux
    port map (
            O => \N__12969\,
            I => \N__12960\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__12966\,
            I => \receive_module.rx_counter.X_5\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__12963\,
            I => \receive_module.rx_counter.X_5\
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__12960\,
            I => \receive_module.rx_counter.X_5\
        );

    \I__2048\ : InMux
    port map (
            O => \N__12953\,
            I => \N__12948\
        );

    \I__2047\ : InMux
    port map (
            O => \N__12952\,
            I => \N__12945\
        );

    \I__2046\ : InMux
    port map (
            O => \N__12951\,
            I => \N__12942\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__12948\,
            I => \receive_module.rx_counter.X_7\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__12945\,
            I => \receive_module.rx_counter.X_7\
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__12942\,
            I => \receive_module.rx_counter.X_7\
        );

    \I__2042\ : InMux
    port map (
            O => \N__12935\,
            I => \N__12932\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__12932\,
            I => \receive_module.rx_counter.n6\
        );

    \I__2040\ : CascadeMux
    port map (
            O => \N__12929\,
            I => \receive_module.rx_counter.n7_cascade_\
        );

    \I__2039\ : InMux
    port map (
            O => \N__12926\,
            I => \N__12923\
        );

    \I__2038\ : LocalMux
    port map (
            O => \N__12923\,
            I => \receive_module.rx_counter.n3225\
        );

    \I__2037\ : InMux
    port map (
            O => \N__12920\,
            I => \N__12917\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__12917\,
            I => \receive_module.rx_counter.old_HS\
        );

    \I__2035\ : CEMux
    port map (
            O => \N__12914\,
            I => \N__12910\
        );

    \I__2034\ : CEMux
    port map (
            O => \N__12913\,
            I => \N__12907\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__12910\,
            I => \receive_module.rx_counter.n2081\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__12907\,
            I => \receive_module.rx_counter.n2081\
        );

    \I__2031\ : SRMux
    port map (
            O => \N__12902\,
            I => \N__12897\
        );

    \I__2030\ : SRMux
    port map (
            O => \N__12901\,
            I => \N__12894\
        );

    \I__2029\ : SRMux
    port map (
            O => \N__12900\,
            I => \N__12891\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__12897\,
            I => \N__12887\
        );

    \I__2027\ : LocalMux
    port map (
            O => \N__12894\,
            I => \N__12882\
        );

    \I__2026\ : LocalMux
    port map (
            O => \N__12891\,
            I => \N__12882\
        );

    \I__2025\ : SRMux
    port map (
            O => \N__12890\,
            I => \N__12879\
        );

    \I__2024\ : Span4Mux_v
    port map (
            O => \N__12887\,
            I => \N__12876\
        );

    \I__2023\ : Span4Mux_v
    port map (
            O => \N__12882\,
            I => \N__12871\
        );

    \I__2022\ : LocalMux
    port map (
            O => \N__12879\,
            I => \N__12871\
        );

    \I__2021\ : Span4Mux_v
    port map (
            O => \N__12876\,
            I => \N__12866\
        );

    \I__2020\ : Span4Mux_v
    port map (
            O => \N__12871\,
            I => \N__12866\
        );

    \I__2019\ : Sp12to4
    port map (
            O => \N__12866\,
            I => \N__12863\
        );

    \I__2018\ : Odrv12
    port map (
            O => \N__12863\,
            I => \line_buffer.n573\
        );

    \I__2017\ : InMux
    port map (
            O => \N__12860\,
            I => \N__12857\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__12857\,
            I => \receive_module.rx_counter.n3429\
        );

    \I__2015\ : InMux
    port map (
            O => \N__12854\,
            I => \N__12849\
        );

    \I__2014\ : InMux
    port map (
            O => \N__12853\,
            I => \N__12846\
        );

    \I__2013\ : InMux
    port map (
            O => \N__12852\,
            I => \N__12843\
        );

    \I__2012\ : LocalMux
    port map (
            O => \N__12849\,
            I => \receive_module.rx_counter.X_8\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__12846\,
            I => \receive_module.rx_counter.X_8\
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__12843\,
            I => \receive_module.rx_counter.X_8\
        );

    \I__2009\ : CascadeMux
    port map (
            O => \N__12836\,
            I => \N__12832\
        );

    \I__2008\ : InMux
    port map (
            O => \N__12835\,
            I => \N__12829\
        );

    \I__2007\ : InMux
    port map (
            O => \N__12832\,
            I => \N__12826\
        );

    \I__2006\ : LocalMux
    port map (
            O => \N__12829\,
            I => \receive_module.rx_counter.X_9\
        );

    \I__2005\ : LocalMux
    port map (
            O => \N__12826\,
            I => \receive_module.rx_counter.X_9\
        );

    \I__2004\ : InMux
    port map (
            O => \N__12821\,
            I => \N__12818\
        );

    \I__2003\ : LocalMux
    port map (
            O => \N__12818\,
            I => \N__12815\
        );

    \I__2002\ : Odrv4
    port map (
            O => \N__12815\,
            I => \receive_module.rx_counter.n39\
        );

    \I__2001\ : InMux
    port map (
            O => \N__12812\,
            I => \N__12807\
        );

    \I__2000\ : InMux
    port map (
            O => \N__12811\,
            I => \N__12804\
        );

    \I__1999\ : InMux
    port map (
            O => \N__12810\,
            I => \N__12801\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__12807\,
            I => \receive_module.rx_counter.Y_6\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__12804\,
            I => \receive_module.rx_counter.Y_6\
        );

    \I__1996\ : LocalMux
    port map (
            O => \N__12801\,
            I => \receive_module.rx_counter.Y_6\
        );

    \I__1995\ : InMux
    port map (
            O => \N__12794\,
            I => \N__12789\
        );

    \I__1994\ : InMux
    port map (
            O => \N__12793\,
            I => \N__12786\
        );

    \I__1993\ : InMux
    port map (
            O => \N__12792\,
            I => \N__12783\
        );

    \I__1992\ : LocalMux
    port map (
            O => \N__12789\,
            I => \receive_module.rx_counter.Y_5\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__12786\,
            I => \receive_module.rx_counter.Y_5\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__12783\,
            I => \receive_module.rx_counter.Y_5\
        );

    \I__1989\ : InMux
    port map (
            O => \N__12776\,
            I => \N__12773\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__12773\,
            I => \N__12770\
        );

    \I__1987\ : Span4Mux_h
    port map (
            O => \N__12770\,
            I => \N__12767\
        );

    \I__1986\ : Span4Mux_h
    port map (
            O => \N__12767\,
            I => \N__12764\
        );

    \I__1985\ : Odrv4
    port map (
            O => \N__12764\,
            I => \line_buffer.n571\
        );

    \I__1984\ : InMux
    port map (
            O => \N__12761\,
            I => \N__12758\
        );

    \I__1983\ : LocalMux
    port map (
            O => \N__12758\,
            I => \N__12755\
        );

    \I__1982\ : Span12Mux_v
    port map (
            O => \N__12755\,
            I => \N__12752\
        );

    \I__1981\ : Span12Mux_v
    port map (
            O => \N__12752\,
            I => \N__12749\
        );

    \I__1980\ : Span12Mux_h
    port map (
            O => \N__12749\,
            I => \N__12746\
        );

    \I__1979\ : Odrv12
    port map (
            O => \N__12746\,
            I => \line_buffer.n563\
        );

    \I__1978\ : InMux
    port map (
            O => \N__12743\,
            I => \N__12740\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__12740\,
            I => \line_buffer.n3534\
        );

    \I__1976\ : InMux
    port map (
            O => \N__12737\,
            I => \N__12734\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__12734\,
            I => \N__12731\
        );

    \I__1974\ : Odrv4
    port map (
            O => \N__12731\,
            I => \TX_DATA_7\
        );

    \I__1973\ : IoInMux
    port map (
            O => \N__12728\,
            I => \N__12723\
        );

    \I__1972\ : IoInMux
    port map (
            O => \N__12727\,
            I => \N__12720\
        );

    \I__1971\ : IoInMux
    port map (
            O => \N__12726\,
            I => \N__12717\
        );

    \I__1970\ : LocalMux
    port map (
            O => \N__12723\,
            I => \N__12714\
        );

    \I__1969\ : LocalMux
    port map (
            O => \N__12720\,
            I => \N__12711\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__12717\,
            I => \N__12708\
        );

    \I__1967\ : IoSpan4Mux
    port map (
            O => \N__12714\,
            I => \N__12705\
        );

    \I__1966\ : IoSpan4Mux
    port map (
            O => \N__12711\,
            I => \N__12702\
        );

    \I__1965\ : Span12Mux_s8_v
    port map (
            O => \N__12708\,
            I => \N__12699\
        );

    \I__1964\ : Sp12to4
    port map (
            O => \N__12705\,
            I => \N__12696\
        );

    \I__1963\ : Span4Mux_s2_v
    port map (
            O => \N__12702\,
            I => \N__12693\
        );

    \I__1962\ : Span12Mux_h
    port map (
            O => \N__12699\,
            I => \N__12690\
        );

    \I__1961\ : Span12Mux_h
    port map (
            O => \N__12696\,
            I => \N__12687\
        );

    \I__1960\ : Sp12to4
    port map (
            O => \N__12693\,
            I => \N__12684\
        );

    \I__1959\ : Odrv12
    port map (
            O => \N__12690\,
            I => \ADV_B_c\
        );

    \I__1958\ : Odrv12
    port map (
            O => \N__12687\,
            I => \ADV_B_c\
        );

    \I__1957\ : Odrv12
    port map (
            O => \N__12684\,
            I => \ADV_B_c\
        );

    \I__1956\ : InMux
    port map (
            O => \N__12677\,
            I => \N__12674\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__12674\,
            I => \N__12671\
        );

    \I__1954\ : Span12Mux_h
    port map (
            O => \N__12671\,
            I => \N__12668\
        );

    \I__1953\ : Odrv12
    port map (
            O => \N__12668\,
            I => \line_buffer.n474\
        );

    \I__1952\ : InMux
    port map (
            O => \N__12665\,
            I => \N__12662\
        );

    \I__1951\ : LocalMux
    port map (
            O => \N__12662\,
            I => \N__12659\
        );

    \I__1950\ : Span4Mux_h
    port map (
            O => \N__12659\,
            I => \N__12656\
        );

    \I__1949\ : Span4Mux_h
    port map (
            O => \N__12656\,
            I => \N__12653\
        );

    \I__1948\ : Odrv4
    port map (
            O => \N__12653\,
            I => \line_buffer.n466\
        );

    \I__1947\ : InMux
    port map (
            O => \N__12650\,
            I => \N__12647\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__12647\,
            I => \N__12644\
        );

    \I__1945\ : Odrv12
    port map (
            O => \N__12644\,
            I => \line_buffer.n3533\
        );

    \I__1944\ : SRMux
    port map (
            O => \N__12641\,
            I => \N__12636\
        );

    \I__1943\ : SRMux
    port map (
            O => \N__12640\,
            I => \N__12633\
        );

    \I__1942\ : SRMux
    port map (
            O => \N__12639\,
            I => \N__12630\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__12636\,
            I => \N__12627\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__12633\,
            I => \N__12623\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__12630\,
            I => \N__12620\
        );

    \I__1938\ : Span4Mux_h
    port map (
            O => \N__12627\,
            I => \N__12617\
        );

    \I__1937\ : SRMux
    port map (
            O => \N__12626\,
            I => \N__12614\
        );

    \I__1936\ : Span4Mux_v
    port map (
            O => \N__12623\,
            I => \N__12611\
        );

    \I__1935\ : Span4Mux_h
    port map (
            O => \N__12620\,
            I => \N__12608\
        );

    \I__1934\ : Span4Mux_v
    port map (
            O => \N__12617\,
            I => \N__12603\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__12614\,
            I => \N__12603\
        );

    \I__1932\ : Sp12to4
    port map (
            O => \N__12611\,
            I => \N__12600\
        );

    \I__1931\ : Span4Mux_h
    port map (
            O => \N__12608\,
            I => \N__12597\
        );

    \I__1930\ : Span4Mux_h
    port map (
            O => \N__12603\,
            I => \N__12594\
        );

    \I__1929\ : Span12Mux_v
    port map (
            O => \N__12600\,
            I => \N__12591\
        );

    \I__1928\ : Span4Mux_v
    port map (
            O => \N__12597\,
            I => \N__12588\
        );

    \I__1927\ : Span4Mux_h
    port map (
            O => \N__12594\,
            I => \N__12585\
        );

    \I__1926\ : Odrv12
    port map (
            O => \N__12591\,
            I => \line_buffer.n542\
        );

    \I__1925\ : Odrv4
    port map (
            O => \N__12588\,
            I => \line_buffer.n542\
        );

    \I__1924\ : Odrv4
    port map (
            O => \N__12585\,
            I => \line_buffer.n542\
        );

    \I__1923\ : InMux
    port map (
            O => \N__12578\,
            I => \N__12574\
        );

    \I__1922\ : InMux
    port map (
            O => \N__12577\,
            I => \N__12571\
        );

    \I__1921\ : LocalMux
    port map (
            O => \N__12574\,
            I => \receive_module.rx_counter.X_1\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__12571\,
            I => \receive_module.rx_counter.X_1\
        );

    \I__1919\ : InMux
    port map (
            O => \N__12566\,
            I => \N__12562\
        );

    \I__1918\ : InMux
    port map (
            O => \N__12565\,
            I => \N__12559\
        );

    \I__1917\ : LocalMux
    port map (
            O => \N__12562\,
            I => \receive_module.rx_counter.X_0\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__12559\,
            I => \receive_module.rx_counter.X_0\
        );

    \I__1915\ : InMux
    port map (
            O => \N__12554\,
            I => \N__12550\
        );

    \I__1914\ : InMux
    port map (
            O => \N__12553\,
            I => \N__12547\
        );

    \I__1913\ : LocalMux
    port map (
            O => \N__12550\,
            I => \receive_module.rx_counter.X_2\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__12547\,
            I => \receive_module.rx_counter.X_2\
        );

    \I__1911\ : CascadeMux
    port map (
            O => \N__12542\,
            I => \receive_module.rx_counter.n3225_cascade_\
        );

    \I__1910\ : CascadeMux
    port map (
            O => \N__12539\,
            I => \receive_module.rx_counter.n3458_cascade_\
        );

    \I__1909\ : InMux
    port map (
            O => \N__12536\,
            I => \N__12531\
        );

    \I__1908\ : InMux
    port map (
            O => \N__12535\,
            I => \N__12526\
        );

    \I__1907\ : InMux
    port map (
            O => \N__12534\,
            I => \N__12526\
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__12531\,
            I => \receive_module.rx_counter.X_4\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__12526\,
            I => \receive_module.rx_counter.X_4\
        );

    \I__1904\ : InMux
    port map (
            O => \N__12521\,
            I => \N__12516\
        );

    \I__1903\ : InMux
    port map (
            O => \N__12520\,
            I => \N__12511\
        );

    \I__1902\ : InMux
    port map (
            O => \N__12519\,
            I => \N__12511\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__12516\,
            I => \receive_module.rx_counter.X_6\
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__12511\,
            I => \receive_module.rx_counter.X_6\
        );

    \I__1899\ : SRMux
    port map (
            O => \N__12506\,
            I => \N__12503\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__12503\,
            I => \N__12499\
        );

    \I__1897\ : SRMux
    port map (
            O => \N__12502\,
            I => \N__12496\
        );

    \I__1896\ : Span4Mux_h
    port map (
            O => \N__12499\,
            I => \N__12493\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__12496\,
            I => \N__12490\
        );

    \I__1894\ : Odrv4
    port map (
            O => \N__12493\,
            I => \receive_module.rx_counter.n3\
        );

    \I__1893\ : Odrv12
    port map (
            O => \N__12490\,
            I => \receive_module.rx_counter.n3\
        );

    \I__1892\ : InMux
    port map (
            O => \N__12485\,
            I => \N__12480\
        );

    \I__1891\ : InMux
    port map (
            O => \N__12484\,
            I => \N__12477\
        );

    \I__1890\ : CascadeMux
    port map (
            O => \N__12483\,
            I => \N__12474\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__12480\,
            I => \N__12468\
        );

    \I__1888\ : LocalMux
    port map (
            O => \N__12477\,
            I => \N__12468\
        );

    \I__1887\ : InMux
    port map (
            O => \N__12474\,
            I => \N__12463\
        );

    \I__1886\ : InMux
    port map (
            O => \N__12473\,
            I => \N__12463\
        );

    \I__1885\ : Odrv4
    port map (
            O => \N__12468\,
            I => \transmit_module.video_signal_controller.VGA_X_2\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__12463\,
            I => \transmit_module.video_signal_controller.VGA_X_2\
        );

    \I__1883\ : InMux
    port map (
            O => \N__12458\,
            I => \N__12452\
        );

    \I__1882\ : InMux
    port map (
            O => \N__12457\,
            I => \N__12449\
        );

    \I__1881\ : InMux
    port map (
            O => \N__12456\,
            I => \N__12444\
        );

    \I__1880\ : InMux
    port map (
            O => \N__12455\,
            I => \N__12444\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__12452\,
            I => \N__12439\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__12449\,
            I => \N__12439\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__12444\,
            I => \transmit_module.video_signal_controller.VGA_X_1\
        );

    \I__1876\ : Odrv4
    port map (
            O => \N__12439\,
            I => \transmit_module.video_signal_controller.VGA_X_1\
        );

    \I__1875\ : InMux
    port map (
            O => \N__12434\,
            I => \N__12431\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__12431\,
            I => \transmit_module.video_signal_controller.n3679\
        );

    \I__1873\ : InMux
    port map (
            O => \N__12428\,
            I => \N__12424\
        );

    \I__1872\ : InMux
    port map (
            O => \N__12427\,
            I => \N__12421\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__12424\,
            I => \transmit_module.n108\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__12421\,
            I => \transmit_module.n108\
        );

    \I__1869\ : InMux
    port map (
            O => \N__12416\,
            I => \N__12412\
        );

    \I__1868\ : InMux
    port map (
            O => \N__12415\,
            I => \N__12409\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__12412\,
            I => \N__12403\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__12409\,
            I => \N__12400\
        );

    \I__1865\ : InMux
    port map (
            O => \N__12408\,
            I => \N__12397\
        );

    \I__1864\ : InMux
    port map (
            O => \N__12407\,
            I => \N__12394\
        );

    \I__1863\ : InMux
    port map (
            O => \N__12406\,
            I => \N__12391\
        );

    \I__1862\ : Span4Mux_v
    port map (
            O => \N__12403\,
            I => \N__12384\
        );

    \I__1861\ : Span4Mux_v
    port map (
            O => \N__12400\,
            I => \N__12384\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__12397\,
            I => \N__12384\
        );

    \I__1859\ : LocalMux
    port map (
            O => \N__12394\,
            I => \transmit_module.video_signal_controller.VGA_X_9\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__12391\,
            I => \transmit_module.video_signal_controller.VGA_X_9\
        );

    \I__1857\ : Odrv4
    port map (
            O => \N__12384\,
            I => \transmit_module.video_signal_controller.VGA_X_9\
        );

    \I__1856\ : InMux
    port map (
            O => \N__12377\,
            I => \N__12374\
        );

    \I__1855\ : LocalMux
    port map (
            O => \N__12374\,
            I => \transmit_module.video_signal_controller.n6_adj_623\
        );

    \I__1854\ : InMux
    port map (
            O => \N__12371\,
            I => \N__12367\
        );

    \I__1853\ : InMux
    port map (
            O => \N__12370\,
            I => \N__12364\
        );

    \I__1852\ : LocalMux
    port map (
            O => \N__12367\,
            I => \transmit_module.n139\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__12364\,
            I => \transmit_module.n139\
        );

    \I__1850\ : CascadeMux
    port map (
            O => \N__12359\,
            I => \transmit_module.n138_cascade_\
        );

    \I__1849\ : CascadeMux
    port map (
            O => \N__12356\,
            I => \N__12352\
        );

    \I__1848\ : CascadeMux
    port map (
            O => \N__12355\,
            I => \N__12349\
        );

    \I__1847\ : CascadeBuf
    port map (
            O => \N__12352\,
            I => \N__12346\
        );

    \I__1846\ : CascadeBuf
    port map (
            O => \N__12349\,
            I => \N__12343\
        );

    \I__1845\ : CascadeMux
    port map (
            O => \N__12346\,
            I => \N__12340\
        );

    \I__1844\ : CascadeMux
    port map (
            O => \N__12343\,
            I => \N__12337\
        );

    \I__1843\ : CascadeBuf
    port map (
            O => \N__12340\,
            I => \N__12334\
        );

    \I__1842\ : CascadeBuf
    port map (
            O => \N__12337\,
            I => \N__12331\
        );

    \I__1841\ : CascadeMux
    port map (
            O => \N__12334\,
            I => \N__12328\
        );

    \I__1840\ : CascadeMux
    port map (
            O => \N__12331\,
            I => \N__12325\
        );

    \I__1839\ : CascadeBuf
    port map (
            O => \N__12328\,
            I => \N__12322\
        );

    \I__1838\ : CascadeBuf
    port map (
            O => \N__12325\,
            I => \N__12319\
        );

    \I__1837\ : CascadeMux
    port map (
            O => \N__12322\,
            I => \N__12316\
        );

    \I__1836\ : CascadeMux
    port map (
            O => \N__12319\,
            I => \N__12313\
        );

    \I__1835\ : CascadeBuf
    port map (
            O => \N__12316\,
            I => \N__12310\
        );

    \I__1834\ : CascadeBuf
    port map (
            O => \N__12313\,
            I => \N__12307\
        );

    \I__1833\ : CascadeMux
    port map (
            O => \N__12310\,
            I => \N__12304\
        );

    \I__1832\ : CascadeMux
    port map (
            O => \N__12307\,
            I => \N__12301\
        );

    \I__1831\ : CascadeBuf
    port map (
            O => \N__12304\,
            I => \N__12298\
        );

    \I__1830\ : CascadeBuf
    port map (
            O => \N__12301\,
            I => \N__12295\
        );

    \I__1829\ : CascadeMux
    port map (
            O => \N__12298\,
            I => \N__12292\
        );

    \I__1828\ : CascadeMux
    port map (
            O => \N__12295\,
            I => \N__12289\
        );

    \I__1827\ : CascadeBuf
    port map (
            O => \N__12292\,
            I => \N__12286\
        );

    \I__1826\ : CascadeBuf
    port map (
            O => \N__12289\,
            I => \N__12283\
        );

    \I__1825\ : CascadeMux
    port map (
            O => \N__12286\,
            I => \N__12280\
        );

    \I__1824\ : CascadeMux
    port map (
            O => \N__12283\,
            I => \N__12277\
        );

    \I__1823\ : CascadeBuf
    port map (
            O => \N__12280\,
            I => \N__12274\
        );

    \I__1822\ : CascadeBuf
    port map (
            O => \N__12277\,
            I => \N__12271\
        );

    \I__1821\ : CascadeMux
    port map (
            O => \N__12274\,
            I => \N__12268\
        );

    \I__1820\ : CascadeMux
    port map (
            O => \N__12271\,
            I => \N__12265\
        );

    \I__1819\ : CascadeBuf
    port map (
            O => \N__12268\,
            I => \N__12262\
        );

    \I__1818\ : CascadeBuf
    port map (
            O => \N__12265\,
            I => \N__12259\
        );

    \I__1817\ : CascadeMux
    port map (
            O => \N__12262\,
            I => \N__12256\
        );

    \I__1816\ : CascadeMux
    port map (
            O => \N__12259\,
            I => \N__12253\
        );

    \I__1815\ : CascadeBuf
    port map (
            O => \N__12256\,
            I => \N__12250\
        );

    \I__1814\ : CascadeBuf
    port map (
            O => \N__12253\,
            I => \N__12247\
        );

    \I__1813\ : CascadeMux
    port map (
            O => \N__12250\,
            I => \N__12244\
        );

    \I__1812\ : CascadeMux
    port map (
            O => \N__12247\,
            I => \N__12241\
        );

    \I__1811\ : CascadeBuf
    port map (
            O => \N__12244\,
            I => \N__12238\
        );

    \I__1810\ : CascadeBuf
    port map (
            O => \N__12241\,
            I => \N__12235\
        );

    \I__1809\ : CascadeMux
    port map (
            O => \N__12238\,
            I => \N__12232\
        );

    \I__1808\ : CascadeMux
    port map (
            O => \N__12235\,
            I => \N__12229\
        );

    \I__1807\ : CascadeBuf
    port map (
            O => \N__12232\,
            I => \N__12226\
        );

    \I__1806\ : CascadeBuf
    port map (
            O => \N__12229\,
            I => \N__12223\
        );

    \I__1805\ : CascadeMux
    port map (
            O => \N__12226\,
            I => \N__12220\
        );

    \I__1804\ : CascadeMux
    port map (
            O => \N__12223\,
            I => \N__12217\
        );

    \I__1803\ : CascadeBuf
    port map (
            O => \N__12220\,
            I => \N__12214\
        );

    \I__1802\ : CascadeBuf
    port map (
            O => \N__12217\,
            I => \N__12211\
        );

    \I__1801\ : CascadeMux
    port map (
            O => \N__12214\,
            I => \N__12208\
        );

    \I__1800\ : CascadeMux
    port map (
            O => \N__12211\,
            I => \N__12205\
        );

    \I__1799\ : CascadeBuf
    port map (
            O => \N__12208\,
            I => \N__12202\
        );

    \I__1798\ : CascadeBuf
    port map (
            O => \N__12205\,
            I => \N__12199\
        );

    \I__1797\ : CascadeMux
    port map (
            O => \N__12202\,
            I => \N__12196\
        );

    \I__1796\ : CascadeMux
    port map (
            O => \N__12199\,
            I => \N__12193\
        );

    \I__1795\ : CascadeBuf
    port map (
            O => \N__12196\,
            I => \N__12190\
        );

    \I__1794\ : CascadeBuf
    port map (
            O => \N__12193\,
            I => \N__12187\
        );

    \I__1793\ : CascadeMux
    port map (
            O => \N__12190\,
            I => \N__12184\
        );

    \I__1792\ : CascadeMux
    port map (
            O => \N__12187\,
            I => \N__12181\
        );

    \I__1791\ : CascadeBuf
    port map (
            O => \N__12184\,
            I => \N__12178\
        );

    \I__1790\ : CascadeBuf
    port map (
            O => \N__12181\,
            I => \N__12175\
        );

    \I__1789\ : CascadeMux
    port map (
            O => \N__12178\,
            I => \N__12172\
        );

    \I__1788\ : CascadeMux
    port map (
            O => \N__12175\,
            I => \N__12169\
        );

    \I__1787\ : InMux
    port map (
            O => \N__12172\,
            I => \N__12166\
        );

    \I__1786\ : InMux
    port map (
            O => \N__12169\,
            I => \N__12163\
        );

    \I__1785\ : LocalMux
    port map (
            O => \N__12166\,
            I => \N__12160\
        );

    \I__1784\ : LocalMux
    port map (
            O => \N__12163\,
            I => \N__12157\
        );

    \I__1783\ : Span12Mux_s7_v
    port map (
            O => \N__12160\,
            I => \N__12154\
        );

    \I__1782\ : Span12Mux_h
    port map (
            O => \N__12157\,
            I => \N__12151\
        );

    \I__1781\ : Span12Mux_h
    port map (
            O => \N__12154\,
            I => \N__12148\
        );

    \I__1780\ : Span12Mux_v
    port map (
            O => \N__12151\,
            I => \N__12145\
        );

    \I__1779\ : Odrv12
    port map (
            O => \N__12148\,
            I => n19
        );

    \I__1778\ : Odrv12
    port map (
            O => \N__12145\,
            I => n19
        );

    \I__1777\ : InMux
    port map (
            O => \N__12140\,
            I => \N__12137\
        );

    \I__1776\ : LocalMux
    port map (
            O => \N__12137\,
            I => \N__12134\
        );

    \I__1775\ : Odrv12
    port map (
            O => \N__12134\,
            I => \line_buffer.n3531\
        );

    \I__1774\ : InMux
    port map (
            O => \N__12131\,
            I => \N__12128\
        );

    \I__1773\ : LocalMux
    port map (
            O => \N__12128\,
            I => \N__12125\
        );

    \I__1772\ : Span4Mux_v
    port map (
            O => \N__12125\,
            I => \N__12122\
        );

    \I__1771\ : Odrv4
    port map (
            O => \N__12122\,
            I => \line_buffer.n3530\
        );

    \I__1770\ : InMux
    port map (
            O => \N__12119\,
            I => \N__12116\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__12116\,
            I => \line_buffer.n3620\
        );

    \I__1768\ : InMux
    port map (
            O => \N__12113\,
            I => \N__12110\
        );

    \I__1767\ : LocalMux
    port map (
            O => \N__12110\,
            I => \transmit_module.n142\
        );

    \I__1766\ : CascadeMux
    port map (
            O => \N__12107\,
            I => \transmit_module.n142_cascade_\
        );

    \I__1765\ : InMux
    port map (
            O => \N__12104\,
            I => \N__12098\
        );

    \I__1764\ : InMux
    port map (
            O => \N__12103\,
            I => \N__12098\
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__12098\,
            I => \transmit_module.n111\
        );

    \I__1762\ : CascadeMux
    port map (
            O => \N__12095\,
            I => \N__12092\
        );

    \I__1761\ : CascadeBuf
    port map (
            O => \N__12092\,
            I => \N__12088\
        );

    \I__1760\ : CascadeMux
    port map (
            O => \N__12091\,
            I => \N__12085\
        );

    \I__1759\ : CascadeMux
    port map (
            O => \N__12088\,
            I => \N__12082\
        );

    \I__1758\ : CascadeBuf
    port map (
            O => \N__12085\,
            I => \N__12079\
        );

    \I__1757\ : CascadeBuf
    port map (
            O => \N__12082\,
            I => \N__12076\
        );

    \I__1756\ : CascadeMux
    port map (
            O => \N__12079\,
            I => \N__12073\
        );

    \I__1755\ : CascadeMux
    port map (
            O => \N__12076\,
            I => \N__12070\
        );

    \I__1754\ : CascadeBuf
    port map (
            O => \N__12073\,
            I => \N__12067\
        );

    \I__1753\ : CascadeBuf
    port map (
            O => \N__12070\,
            I => \N__12064\
        );

    \I__1752\ : CascadeMux
    port map (
            O => \N__12067\,
            I => \N__12061\
        );

    \I__1751\ : CascadeMux
    port map (
            O => \N__12064\,
            I => \N__12058\
        );

    \I__1750\ : CascadeBuf
    port map (
            O => \N__12061\,
            I => \N__12055\
        );

    \I__1749\ : CascadeBuf
    port map (
            O => \N__12058\,
            I => \N__12052\
        );

    \I__1748\ : CascadeMux
    port map (
            O => \N__12055\,
            I => \N__12049\
        );

    \I__1747\ : CascadeMux
    port map (
            O => \N__12052\,
            I => \N__12046\
        );

    \I__1746\ : CascadeBuf
    port map (
            O => \N__12049\,
            I => \N__12043\
        );

    \I__1745\ : CascadeBuf
    port map (
            O => \N__12046\,
            I => \N__12040\
        );

    \I__1744\ : CascadeMux
    port map (
            O => \N__12043\,
            I => \N__12037\
        );

    \I__1743\ : CascadeMux
    port map (
            O => \N__12040\,
            I => \N__12034\
        );

    \I__1742\ : CascadeBuf
    port map (
            O => \N__12037\,
            I => \N__12031\
        );

    \I__1741\ : CascadeBuf
    port map (
            O => \N__12034\,
            I => \N__12028\
        );

    \I__1740\ : CascadeMux
    port map (
            O => \N__12031\,
            I => \N__12025\
        );

    \I__1739\ : CascadeMux
    port map (
            O => \N__12028\,
            I => \N__12022\
        );

    \I__1738\ : CascadeBuf
    port map (
            O => \N__12025\,
            I => \N__12019\
        );

    \I__1737\ : CascadeBuf
    port map (
            O => \N__12022\,
            I => \N__12016\
        );

    \I__1736\ : CascadeMux
    port map (
            O => \N__12019\,
            I => \N__12013\
        );

    \I__1735\ : CascadeMux
    port map (
            O => \N__12016\,
            I => \N__12010\
        );

    \I__1734\ : CascadeBuf
    port map (
            O => \N__12013\,
            I => \N__12007\
        );

    \I__1733\ : CascadeBuf
    port map (
            O => \N__12010\,
            I => \N__12004\
        );

    \I__1732\ : CascadeMux
    port map (
            O => \N__12007\,
            I => \N__12001\
        );

    \I__1731\ : CascadeMux
    port map (
            O => \N__12004\,
            I => \N__11998\
        );

    \I__1730\ : CascadeBuf
    port map (
            O => \N__12001\,
            I => \N__11995\
        );

    \I__1729\ : CascadeBuf
    port map (
            O => \N__11998\,
            I => \N__11992\
        );

    \I__1728\ : CascadeMux
    port map (
            O => \N__11995\,
            I => \N__11989\
        );

    \I__1727\ : CascadeMux
    port map (
            O => \N__11992\,
            I => \N__11986\
        );

    \I__1726\ : CascadeBuf
    port map (
            O => \N__11989\,
            I => \N__11983\
        );

    \I__1725\ : CascadeBuf
    port map (
            O => \N__11986\,
            I => \N__11980\
        );

    \I__1724\ : CascadeMux
    port map (
            O => \N__11983\,
            I => \N__11977\
        );

    \I__1723\ : CascadeMux
    port map (
            O => \N__11980\,
            I => \N__11974\
        );

    \I__1722\ : CascadeBuf
    port map (
            O => \N__11977\,
            I => \N__11971\
        );

    \I__1721\ : CascadeBuf
    port map (
            O => \N__11974\,
            I => \N__11968\
        );

    \I__1720\ : CascadeMux
    port map (
            O => \N__11971\,
            I => \N__11965\
        );

    \I__1719\ : CascadeMux
    port map (
            O => \N__11968\,
            I => \N__11962\
        );

    \I__1718\ : CascadeBuf
    port map (
            O => \N__11965\,
            I => \N__11959\
        );

    \I__1717\ : CascadeBuf
    port map (
            O => \N__11962\,
            I => \N__11956\
        );

    \I__1716\ : CascadeMux
    port map (
            O => \N__11959\,
            I => \N__11953\
        );

    \I__1715\ : CascadeMux
    port map (
            O => \N__11956\,
            I => \N__11950\
        );

    \I__1714\ : CascadeBuf
    port map (
            O => \N__11953\,
            I => \N__11947\
        );

    \I__1713\ : CascadeBuf
    port map (
            O => \N__11950\,
            I => \N__11944\
        );

    \I__1712\ : CascadeMux
    port map (
            O => \N__11947\,
            I => \N__11941\
        );

    \I__1711\ : CascadeMux
    port map (
            O => \N__11944\,
            I => \N__11938\
        );

    \I__1710\ : CascadeBuf
    port map (
            O => \N__11941\,
            I => \N__11935\
        );

    \I__1709\ : CascadeBuf
    port map (
            O => \N__11938\,
            I => \N__11932\
        );

    \I__1708\ : CascadeMux
    port map (
            O => \N__11935\,
            I => \N__11929\
        );

    \I__1707\ : CascadeMux
    port map (
            O => \N__11932\,
            I => \N__11926\
        );

    \I__1706\ : CascadeBuf
    port map (
            O => \N__11929\,
            I => \N__11923\
        );

    \I__1705\ : CascadeBuf
    port map (
            O => \N__11926\,
            I => \N__11920\
        );

    \I__1704\ : CascadeMux
    port map (
            O => \N__11923\,
            I => \N__11917\
        );

    \I__1703\ : CascadeMux
    port map (
            O => \N__11920\,
            I => \N__11914\
        );

    \I__1702\ : CascadeBuf
    port map (
            O => \N__11917\,
            I => \N__11911\
        );

    \I__1701\ : InMux
    port map (
            O => \N__11914\,
            I => \N__11908\
        );

    \I__1700\ : CascadeMux
    port map (
            O => \N__11911\,
            I => \N__11905\
        );

    \I__1699\ : LocalMux
    port map (
            O => \N__11908\,
            I => \N__11902\
        );

    \I__1698\ : InMux
    port map (
            O => \N__11905\,
            I => \N__11899\
        );

    \I__1697\ : Span4Mux_v
    port map (
            O => \N__11902\,
            I => \N__11896\
        );

    \I__1696\ : LocalMux
    port map (
            O => \N__11899\,
            I => \N__11893\
        );

    \I__1695\ : Span4Mux_v
    port map (
            O => \N__11896\,
            I => \N__11890\
        );

    \I__1694\ : Span12Mux_s9_v
    port map (
            O => \N__11893\,
            I => \N__11887\
        );

    \I__1693\ : Span4Mux_v
    port map (
            O => \N__11890\,
            I => \N__11884\
        );

    \I__1692\ : Span12Mux_h
    port map (
            O => \N__11887\,
            I => \N__11881\
        );

    \I__1691\ : Span4Mux_h
    port map (
            O => \N__11884\,
            I => \N__11878\
        );

    \I__1690\ : Odrv12
    port map (
            O => \N__11881\,
            I => n23
        );

    \I__1689\ : Odrv4
    port map (
            O => \N__11878\,
            I => n23
        );

    \I__1688\ : InMux
    port map (
            O => \N__11873\,
            I => \N__11869\
        );

    \I__1687\ : InMux
    port map (
            O => \N__11872\,
            I => \N__11866\
        );

    \I__1686\ : LocalMux
    port map (
            O => \N__11869\,
            I => \transmit_module.video_signal_controller.n3366\
        );

    \I__1685\ : LocalMux
    port map (
            O => \N__11866\,
            I => \transmit_module.video_signal_controller.n3366\
        );

    \I__1684\ : CascadeMux
    port map (
            O => \N__11861\,
            I => \N__11857\
        );

    \I__1683\ : InMux
    port map (
            O => \N__11860\,
            I => \N__11853\
        );

    \I__1682\ : InMux
    port map (
            O => \N__11857\,
            I => \N__11850\
        );

    \I__1681\ : InMux
    port map (
            O => \N__11856\,
            I => \N__11847\
        );

    \I__1680\ : LocalMux
    port map (
            O => \N__11853\,
            I => \N__11843\
        );

    \I__1679\ : LocalMux
    port map (
            O => \N__11850\,
            I => \N__11840\
        );

    \I__1678\ : LocalMux
    port map (
            O => \N__11847\,
            I => \N__11837\
        );

    \I__1677\ : InMux
    port map (
            O => \N__11846\,
            I => \N__11834\
        );

    \I__1676\ : Span4Mux_v
    port map (
            O => \N__11843\,
            I => \N__11829\
        );

    \I__1675\ : Span4Mux_v
    port map (
            O => \N__11840\,
            I => \N__11829\
        );

    \I__1674\ : Span4Mux_h
    port map (
            O => \N__11837\,
            I => \N__11826\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__11834\,
            I => \transmit_module.video_signal_controller.VGA_X_8\
        );

    \I__1672\ : Odrv4
    port map (
            O => \N__11829\,
            I => \transmit_module.video_signal_controller.VGA_X_8\
        );

    \I__1671\ : Odrv4
    port map (
            O => \N__11826\,
            I => \transmit_module.video_signal_controller.VGA_X_8\
        );

    \I__1670\ : InMux
    port map (
            O => \N__11819\,
            I => \N__11815\
        );

    \I__1669\ : InMux
    port map (
            O => \N__11818\,
            I => \N__11812\
        );

    \I__1668\ : LocalMux
    port map (
            O => \N__11815\,
            I => \N__11809\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__11812\,
            I => \transmit_module.video_signal_controller.n2017\
        );

    \I__1666\ : Odrv4
    port map (
            O => \N__11809\,
            I => \transmit_module.video_signal_controller.n2017\
        );

    \I__1665\ : CascadeMux
    port map (
            O => \N__11804\,
            I => \transmit_module.video_signal_controller.n3007_cascade_\
        );

    \I__1664\ : InMux
    port map (
            O => \N__11801\,
            I => \N__11797\
        );

    \I__1663\ : InMux
    port map (
            O => \N__11800\,
            I => \N__11794\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__11797\,
            I => \transmit_module.video_signal_controller.VGA_VISIBLE_N_588\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__11794\,
            I => \transmit_module.video_signal_controller.VGA_VISIBLE_N_588\
        );

    \I__1660\ : InMux
    port map (
            O => \N__11789\,
            I => \N__11786\
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__11786\,
            I => \transmit_module.n143\
        );

    \I__1658\ : CascadeMux
    port map (
            O => \N__11783\,
            I => \transmit_module.n143_cascade_\
        );

    \I__1657\ : CascadeMux
    port map (
            O => \N__11780\,
            I => \N__11776\
        );

    \I__1656\ : CascadeMux
    port map (
            O => \N__11779\,
            I => \N__11773\
        );

    \I__1655\ : CascadeBuf
    port map (
            O => \N__11776\,
            I => \N__11770\
        );

    \I__1654\ : CascadeBuf
    port map (
            O => \N__11773\,
            I => \N__11767\
        );

    \I__1653\ : CascadeMux
    port map (
            O => \N__11770\,
            I => \N__11764\
        );

    \I__1652\ : CascadeMux
    port map (
            O => \N__11767\,
            I => \N__11761\
        );

    \I__1651\ : CascadeBuf
    port map (
            O => \N__11764\,
            I => \N__11758\
        );

    \I__1650\ : CascadeBuf
    port map (
            O => \N__11761\,
            I => \N__11755\
        );

    \I__1649\ : CascadeMux
    port map (
            O => \N__11758\,
            I => \N__11752\
        );

    \I__1648\ : CascadeMux
    port map (
            O => \N__11755\,
            I => \N__11749\
        );

    \I__1647\ : CascadeBuf
    port map (
            O => \N__11752\,
            I => \N__11746\
        );

    \I__1646\ : CascadeBuf
    port map (
            O => \N__11749\,
            I => \N__11743\
        );

    \I__1645\ : CascadeMux
    port map (
            O => \N__11746\,
            I => \N__11740\
        );

    \I__1644\ : CascadeMux
    port map (
            O => \N__11743\,
            I => \N__11737\
        );

    \I__1643\ : CascadeBuf
    port map (
            O => \N__11740\,
            I => \N__11734\
        );

    \I__1642\ : CascadeBuf
    port map (
            O => \N__11737\,
            I => \N__11731\
        );

    \I__1641\ : CascadeMux
    port map (
            O => \N__11734\,
            I => \N__11728\
        );

    \I__1640\ : CascadeMux
    port map (
            O => \N__11731\,
            I => \N__11725\
        );

    \I__1639\ : CascadeBuf
    port map (
            O => \N__11728\,
            I => \N__11722\
        );

    \I__1638\ : CascadeBuf
    port map (
            O => \N__11725\,
            I => \N__11719\
        );

    \I__1637\ : CascadeMux
    port map (
            O => \N__11722\,
            I => \N__11716\
        );

    \I__1636\ : CascadeMux
    port map (
            O => \N__11719\,
            I => \N__11713\
        );

    \I__1635\ : CascadeBuf
    port map (
            O => \N__11716\,
            I => \N__11710\
        );

    \I__1634\ : CascadeBuf
    port map (
            O => \N__11713\,
            I => \N__11707\
        );

    \I__1633\ : CascadeMux
    port map (
            O => \N__11710\,
            I => \N__11704\
        );

    \I__1632\ : CascadeMux
    port map (
            O => \N__11707\,
            I => \N__11701\
        );

    \I__1631\ : CascadeBuf
    port map (
            O => \N__11704\,
            I => \N__11698\
        );

    \I__1630\ : CascadeBuf
    port map (
            O => \N__11701\,
            I => \N__11695\
        );

    \I__1629\ : CascadeMux
    port map (
            O => \N__11698\,
            I => \N__11692\
        );

    \I__1628\ : CascadeMux
    port map (
            O => \N__11695\,
            I => \N__11689\
        );

    \I__1627\ : CascadeBuf
    port map (
            O => \N__11692\,
            I => \N__11686\
        );

    \I__1626\ : CascadeBuf
    port map (
            O => \N__11689\,
            I => \N__11683\
        );

    \I__1625\ : CascadeMux
    port map (
            O => \N__11686\,
            I => \N__11680\
        );

    \I__1624\ : CascadeMux
    port map (
            O => \N__11683\,
            I => \N__11677\
        );

    \I__1623\ : CascadeBuf
    port map (
            O => \N__11680\,
            I => \N__11674\
        );

    \I__1622\ : CascadeBuf
    port map (
            O => \N__11677\,
            I => \N__11671\
        );

    \I__1621\ : CascadeMux
    port map (
            O => \N__11674\,
            I => \N__11668\
        );

    \I__1620\ : CascadeMux
    port map (
            O => \N__11671\,
            I => \N__11665\
        );

    \I__1619\ : CascadeBuf
    port map (
            O => \N__11668\,
            I => \N__11662\
        );

    \I__1618\ : CascadeBuf
    port map (
            O => \N__11665\,
            I => \N__11659\
        );

    \I__1617\ : CascadeMux
    port map (
            O => \N__11662\,
            I => \N__11656\
        );

    \I__1616\ : CascadeMux
    port map (
            O => \N__11659\,
            I => \N__11653\
        );

    \I__1615\ : CascadeBuf
    port map (
            O => \N__11656\,
            I => \N__11650\
        );

    \I__1614\ : CascadeBuf
    port map (
            O => \N__11653\,
            I => \N__11647\
        );

    \I__1613\ : CascadeMux
    port map (
            O => \N__11650\,
            I => \N__11644\
        );

    \I__1612\ : CascadeMux
    port map (
            O => \N__11647\,
            I => \N__11641\
        );

    \I__1611\ : CascadeBuf
    port map (
            O => \N__11644\,
            I => \N__11638\
        );

    \I__1610\ : CascadeBuf
    port map (
            O => \N__11641\,
            I => \N__11635\
        );

    \I__1609\ : CascadeMux
    port map (
            O => \N__11638\,
            I => \N__11632\
        );

    \I__1608\ : CascadeMux
    port map (
            O => \N__11635\,
            I => \N__11629\
        );

    \I__1607\ : CascadeBuf
    port map (
            O => \N__11632\,
            I => \N__11626\
        );

    \I__1606\ : CascadeBuf
    port map (
            O => \N__11629\,
            I => \N__11623\
        );

    \I__1605\ : CascadeMux
    port map (
            O => \N__11626\,
            I => \N__11620\
        );

    \I__1604\ : CascadeMux
    port map (
            O => \N__11623\,
            I => \N__11617\
        );

    \I__1603\ : CascadeBuf
    port map (
            O => \N__11620\,
            I => \N__11614\
        );

    \I__1602\ : CascadeBuf
    port map (
            O => \N__11617\,
            I => \N__11611\
        );

    \I__1601\ : CascadeMux
    port map (
            O => \N__11614\,
            I => \N__11608\
        );

    \I__1600\ : CascadeMux
    port map (
            O => \N__11611\,
            I => \N__11605\
        );

    \I__1599\ : CascadeBuf
    port map (
            O => \N__11608\,
            I => \N__11602\
        );

    \I__1598\ : CascadeBuf
    port map (
            O => \N__11605\,
            I => \N__11599\
        );

    \I__1597\ : CascadeMux
    port map (
            O => \N__11602\,
            I => \N__11596\
        );

    \I__1596\ : CascadeMux
    port map (
            O => \N__11599\,
            I => \N__11593\
        );

    \I__1595\ : InMux
    port map (
            O => \N__11596\,
            I => \N__11590\
        );

    \I__1594\ : InMux
    port map (
            O => \N__11593\,
            I => \N__11587\
        );

    \I__1593\ : LocalMux
    port map (
            O => \N__11590\,
            I => \N__11584\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__11587\,
            I => \N__11581\
        );

    \I__1591\ : Span4Mux_v
    port map (
            O => \N__11584\,
            I => \N__11578\
        );

    \I__1590\ : Span4Mux_v
    port map (
            O => \N__11581\,
            I => \N__11575\
        );

    \I__1589\ : Span4Mux_v
    port map (
            O => \N__11578\,
            I => \N__11572\
        );

    \I__1588\ : Sp12to4
    port map (
            O => \N__11575\,
            I => \N__11569\
        );

    \I__1587\ : Span4Mux_v
    port map (
            O => \N__11572\,
            I => \N__11566\
        );

    \I__1586\ : Span12Mux_v
    port map (
            O => \N__11569\,
            I => \N__11563\
        );

    \I__1585\ : Span4Mux_h
    port map (
            O => \N__11566\,
            I => \N__11560\
        );

    \I__1584\ : Odrv12
    port map (
            O => \N__11563\,
            I => n24
        );

    \I__1583\ : Odrv4
    port map (
            O => \N__11560\,
            I => n24
        );

    \I__1582\ : InMux
    port map (
            O => \N__11555\,
            I => \N__11549\
        );

    \I__1581\ : InMux
    port map (
            O => \N__11554\,
            I => \N__11549\
        );

    \I__1580\ : LocalMux
    port map (
            O => \N__11549\,
            I => \N__11545\
        );

    \I__1579\ : InMux
    port map (
            O => \N__11548\,
            I => \N__11540\
        );

    \I__1578\ : Span4Mux_h
    port map (
            O => \N__11545\,
            I => \N__11537\
        );

    \I__1577\ : InMux
    port map (
            O => \N__11544\,
            I => \N__11534\
        );

    \I__1576\ : InMux
    port map (
            O => \N__11543\,
            I => \N__11531\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__11540\,
            I => \transmit_module.video_signal_controller.VGA_X_10\
        );

    \I__1574\ : Odrv4
    port map (
            O => \N__11537\,
            I => \transmit_module.video_signal_controller.VGA_X_10\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__11534\,
            I => \transmit_module.video_signal_controller.VGA_X_10\
        );

    \I__1572\ : LocalMux
    port map (
            O => \N__11531\,
            I => \transmit_module.video_signal_controller.VGA_X_10\
        );

    \I__1571\ : InMux
    port map (
            O => \N__11522\,
            I => \N__11519\
        );

    \I__1570\ : LocalMux
    port map (
            O => \N__11519\,
            I => \transmit_module.video_signal_controller.n3007\
        );

    \I__1569\ : CascadeMux
    port map (
            O => \N__11516\,
            I => \transmit_module.n141_cascade_\
        );

    \I__1568\ : CascadeMux
    port map (
            O => \N__11513\,
            I => \N__11510\
        );

    \I__1567\ : CascadeBuf
    port map (
            O => \N__11510\,
            I => \N__11507\
        );

    \I__1566\ : CascadeMux
    port map (
            O => \N__11507\,
            I => \N__11504\
        );

    \I__1565\ : CascadeBuf
    port map (
            O => \N__11504\,
            I => \N__11500\
        );

    \I__1564\ : CascadeMux
    port map (
            O => \N__11503\,
            I => \N__11497\
        );

    \I__1563\ : CascadeMux
    port map (
            O => \N__11500\,
            I => \N__11494\
        );

    \I__1562\ : CascadeBuf
    port map (
            O => \N__11497\,
            I => \N__11491\
        );

    \I__1561\ : CascadeBuf
    port map (
            O => \N__11494\,
            I => \N__11488\
        );

    \I__1560\ : CascadeMux
    port map (
            O => \N__11491\,
            I => \N__11485\
        );

    \I__1559\ : CascadeMux
    port map (
            O => \N__11488\,
            I => \N__11482\
        );

    \I__1558\ : CascadeBuf
    port map (
            O => \N__11485\,
            I => \N__11479\
        );

    \I__1557\ : CascadeBuf
    port map (
            O => \N__11482\,
            I => \N__11476\
        );

    \I__1556\ : CascadeMux
    port map (
            O => \N__11479\,
            I => \N__11473\
        );

    \I__1555\ : CascadeMux
    port map (
            O => \N__11476\,
            I => \N__11470\
        );

    \I__1554\ : CascadeBuf
    port map (
            O => \N__11473\,
            I => \N__11467\
        );

    \I__1553\ : CascadeBuf
    port map (
            O => \N__11470\,
            I => \N__11464\
        );

    \I__1552\ : CascadeMux
    port map (
            O => \N__11467\,
            I => \N__11461\
        );

    \I__1551\ : CascadeMux
    port map (
            O => \N__11464\,
            I => \N__11458\
        );

    \I__1550\ : CascadeBuf
    port map (
            O => \N__11461\,
            I => \N__11455\
        );

    \I__1549\ : CascadeBuf
    port map (
            O => \N__11458\,
            I => \N__11452\
        );

    \I__1548\ : CascadeMux
    port map (
            O => \N__11455\,
            I => \N__11449\
        );

    \I__1547\ : CascadeMux
    port map (
            O => \N__11452\,
            I => \N__11446\
        );

    \I__1546\ : CascadeBuf
    port map (
            O => \N__11449\,
            I => \N__11443\
        );

    \I__1545\ : CascadeBuf
    port map (
            O => \N__11446\,
            I => \N__11440\
        );

    \I__1544\ : CascadeMux
    port map (
            O => \N__11443\,
            I => \N__11437\
        );

    \I__1543\ : CascadeMux
    port map (
            O => \N__11440\,
            I => \N__11434\
        );

    \I__1542\ : CascadeBuf
    port map (
            O => \N__11437\,
            I => \N__11431\
        );

    \I__1541\ : CascadeBuf
    port map (
            O => \N__11434\,
            I => \N__11428\
        );

    \I__1540\ : CascadeMux
    port map (
            O => \N__11431\,
            I => \N__11425\
        );

    \I__1539\ : CascadeMux
    port map (
            O => \N__11428\,
            I => \N__11422\
        );

    \I__1538\ : CascadeBuf
    port map (
            O => \N__11425\,
            I => \N__11419\
        );

    \I__1537\ : CascadeBuf
    port map (
            O => \N__11422\,
            I => \N__11416\
        );

    \I__1536\ : CascadeMux
    port map (
            O => \N__11419\,
            I => \N__11413\
        );

    \I__1535\ : CascadeMux
    port map (
            O => \N__11416\,
            I => \N__11410\
        );

    \I__1534\ : CascadeBuf
    port map (
            O => \N__11413\,
            I => \N__11407\
        );

    \I__1533\ : CascadeBuf
    port map (
            O => \N__11410\,
            I => \N__11404\
        );

    \I__1532\ : CascadeMux
    port map (
            O => \N__11407\,
            I => \N__11401\
        );

    \I__1531\ : CascadeMux
    port map (
            O => \N__11404\,
            I => \N__11398\
        );

    \I__1530\ : CascadeBuf
    port map (
            O => \N__11401\,
            I => \N__11395\
        );

    \I__1529\ : CascadeBuf
    port map (
            O => \N__11398\,
            I => \N__11392\
        );

    \I__1528\ : CascadeMux
    port map (
            O => \N__11395\,
            I => \N__11389\
        );

    \I__1527\ : CascadeMux
    port map (
            O => \N__11392\,
            I => \N__11386\
        );

    \I__1526\ : CascadeBuf
    port map (
            O => \N__11389\,
            I => \N__11383\
        );

    \I__1525\ : CascadeBuf
    port map (
            O => \N__11386\,
            I => \N__11380\
        );

    \I__1524\ : CascadeMux
    port map (
            O => \N__11383\,
            I => \N__11377\
        );

    \I__1523\ : CascadeMux
    port map (
            O => \N__11380\,
            I => \N__11374\
        );

    \I__1522\ : CascadeBuf
    port map (
            O => \N__11377\,
            I => \N__11371\
        );

    \I__1521\ : CascadeBuf
    port map (
            O => \N__11374\,
            I => \N__11368\
        );

    \I__1520\ : CascadeMux
    port map (
            O => \N__11371\,
            I => \N__11365\
        );

    \I__1519\ : CascadeMux
    port map (
            O => \N__11368\,
            I => \N__11362\
        );

    \I__1518\ : CascadeBuf
    port map (
            O => \N__11365\,
            I => \N__11359\
        );

    \I__1517\ : CascadeBuf
    port map (
            O => \N__11362\,
            I => \N__11356\
        );

    \I__1516\ : CascadeMux
    port map (
            O => \N__11359\,
            I => \N__11353\
        );

    \I__1515\ : CascadeMux
    port map (
            O => \N__11356\,
            I => \N__11350\
        );

    \I__1514\ : CascadeBuf
    port map (
            O => \N__11353\,
            I => \N__11347\
        );

    \I__1513\ : CascadeBuf
    port map (
            O => \N__11350\,
            I => \N__11344\
        );

    \I__1512\ : CascadeMux
    port map (
            O => \N__11347\,
            I => \N__11341\
        );

    \I__1511\ : CascadeMux
    port map (
            O => \N__11344\,
            I => \N__11338\
        );

    \I__1510\ : CascadeBuf
    port map (
            O => \N__11341\,
            I => \N__11335\
        );

    \I__1509\ : InMux
    port map (
            O => \N__11338\,
            I => \N__11332\
        );

    \I__1508\ : CascadeMux
    port map (
            O => \N__11335\,
            I => \N__11329\
        );

    \I__1507\ : LocalMux
    port map (
            O => \N__11332\,
            I => \N__11326\
        );

    \I__1506\ : CascadeBuf
    port map (
            O => \N__11329\,
            I => \N__11323\
        );

    \I__1505\ : Span4Mux_v
    port map (
            O => \N__11326\,
            I => \N__11320\
        );

    \I__1504\ : CascadeMux
    port map (
            O => \N__11323\,
            I => \N__11317\
        );

    \I__1503\ : Span4Mux_v
    port map (
            O => \N__11320\,
            I => \N__11314\
        );

    \I__1502\ : InMux
    port map (
            O => \N__11317\,
            I => \N__11311\
        );

    \I__1501\ : Span4Mux_h
    port map (
            O => \N__11314\,
            I => \N__11308\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__11311\,
            I => \N__11305\
        );

    \I__1499\ : Span4Mux_h
    port map (
            O => \N__11308\,
            I => \N__11302\
        );

    \I__1498\ : Span4Mux_v
    port map (
            O => \N__11305\,
            I => \N__11299\
        );

    \I__1497\ : Span4Mux_h
    port map (
            O => \N__11302\,
            I => \N__11296\
        );

    \I__1496\ : Span4Mux_h
    port map (
            O => \N__11299\,
            I => \N__11293\
        );

    \I__1495\ : Sp12to4
    port map (
            O => \N__11296\,
            I => \N__11288\
        );

    \I__1494\ : Sp12to4
    port map (
            O => \N__11293\,
            I => \N__11288\
        );

    \I__1493\ : Odrv12
    port map (
            O => \N__11288\,
            I => n22
        );

    \I__1492\ : InMux
    port map (
            O => \N__11285\,
            I => \N__11278\
        );

    \I__1491\ : InMux
    port map (
            O => \N__11284\,
            I => \N__11278\
        );

    \I__1490\ : CascadeMux
    port map (
            O => \N__11283\,
            I => \N__11275\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__11278\,
            I => \N__11271\
        );

    \I__1488\ : InMux
    port map (
            O => \N__11275\,
            I => \N__11266\
        );

    \I__1487\ : InMux
    port map (
            O => \N__11274\,
            I => \N__11266\
        );

    \I__1486\ : Odrv4
    port map (
            O => \N__11271\,
            I => \transmit_module.VGA_VISIBLE_Y\
        );

    \I__1485\ : LocalMux
    port map (
            O => \N__11266\,
            I => \transmit_module.VGA_VISIBLE_Y\
        );

    \I__1484\ : InMux
    port map (
            O => \N__11261\,
            I => \N__11258\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__11258\,
            I => \transmit_module.n140\
        );

    \I__1482\ : CascadeMux
    port map (
            O => \N__11255\,
            I => \transmit_module.n140_cascade_\
        );

    \I__1481\ : InMux
    port map (
            O => \N__11252\,
            I => \N__11246\
        );

    \I__1480\ : InMux
    port map (
            O => \N__11251\,
            I => \N__11246\
        );

    \I__1479\ : LocalMux
    port map (
            O => \N__11246\,
            I => \transmit_module.n109\
        );

    \I__1478\ : CascadeMux
    port map (
            O => \N__11243\,
            I => \N__11240\
        );

    \I__1477\ : CascadeBuf
    port map (
            O => \N__11240\,
            I => \N__11236\
        );

    \I__1476\ : CascadeMux
    port map (
            O => \N__11239\,
            I => \N__11233\
        );

    \I__1475\ : CascadeMux
    port map (
            O => \N__11236\,
            I => \N__11230\
        );

    \I__1474\ : CascadeBuf
    port map (
            O => \N__11233\,
            I => \N__11227\
        );

    \I__1473\ : CascadeBuf
    port map (
            O => \N__11230\,
            I => \N__11224\
        );

    \I__1472\ : CascadeMux
    port map (
            O => \N__11227\,
            I => \N__11221\
        );

    \I__1471\ : CascadeMux
    port map (
            O => \N__11224\,
            I => \N__11218\
        );

    \I__1470\ : CascadeBuf
    port map (
            O => \N__11221\,
            I => \N__11215\
        );

    \I__1469\ : CascadeBuf
    port map (
            O => \N__11218\,
            I => \N__11212\
        );

    \I__1468\ : CascadeMux
    port map (
            O => \N__11215\,
            I => \N__11209\
        );

    \I__1467\ : CascadeMux
    port map (
            O => \N__11212\,
            I => \N__11206\
        );

    \I__1466\ : CascadeBuf
    port map (
            O => \N__11209\,
            I => \N__11203\
        );

    \I__1465\ : CascadeBuf
    port map (
            O => \N__11206\,
            I => \N__11200\
        );

    \I__1464\ : CascadeMux
    port map (
            O => \N__11203\,
            I => \N__11197\
        );

    \I__1463\ : CascadeMux
    port map (
            O => \N__11200\,
            I => \N__11194\
        );

    \I__1462\ : CascadeBuf
    port map (
            O => \N__11197\,
            I => \N__11191\
        );

    \I__1461\ : CascadeBuf
    port map (
            O => \N__11194\,
            I => \N__11188\
        );

    \I__1460\ : CascadeMux
    port map (
            O => \N__11191\,
            I => \N__11185\
        );

    \I__1459\ : CascadeMux
    port map (
            O => \N__11188\,
            I => \N__11182\
        );

    \I__1458\ : CascadeBuf
    port map (
            O => \N__11185\,
            I => \N__11179\
        );

    \I__1457\ : CascadeBuf
    port map (
            O => \N__11182\,
            I => \N__11176\
        );

    \I__1456\ : CascadeMux
    port map (
            O => \N__11179\,
            I => \N__11173\
        );

    \I__1455\ : CascadeMux
    port map (
            O => \N__11176\,
            I => \N__11170\
        );

    \I__1454\ : CascadeBuf
    port map (
            O => \N__11173\,
            I => \N__11167\
        );

    \I__1453\ : CascadeBuf
    port map (
            O => \N__11170\,
            I => \N__11164\
        );

    \I__1452\ : CascadeMux
    port map (
            O => \N__11167\,
            I => \N__11161\
        );

    \I__1451\ : CascadeMux
    port map (
            O => \N__11164\,
            I => \N__11158\
        );

    \I__1450\ : CascadeBuf
    port map (
            O => \N__11161\,
            I => \N__11155\
        );

    \I__1449\ : CascadeBuf
    port map (
            O => \N__11158\,
            I => \N__11152\
        );

    \I__1448\ : CascadeMux
    port map (
            O => \N__11155\,
            I => \N__11149\
        );

    \I__1447\ : CascadeMux
    port map (
            O => \N__11152\,
            I => \N__11146\
        );

    \I__1446\ : CascadeBuf
    port map (
            O => \N__11149\,
            I => \N__11143\
        );

    \I__1445\ : CascadeBuf
    port map (
            O => \N__11146\,
            I => \N__11140\
        );

    \I__1444\ : CascadeMux
    port map (
            O => \N__11143\,
            I => \N__11137\
        );

    \I__1443\ : CascadeMux
    port map (
            O => \N__11140\,
            I => \N__11134\
        );

    \I__1442\ : CascadeBuf
    port map (
            O => \N__11137\,
            I => \N__11131\
        );

    \I__1441\ : CascadeBuf
    port map (
            O => \N__11134\,
            I => \N__11128\
        );

    \I__1440\ : CascadeMux
    port map (
            O => \N__11131\,
            I => \N__11125\
        );

    \I__1439\ : CascadeMux
    port map (
            O => \N__11128\,
            I => \N__11122\
        );

    \I__1438\ : CascadeBuf
    port map (
            O => \N__11125\,
            I => \N__11119\
        );

    \I__1437\ : CascadeBuf
    port map (
            O => \N__11122\,
            I => \N__11116\
        );

    \I__1436\ : CascadeMux
    port map (
            O => \N__11119\,
            I => \N__11113\
        );

    \I__1435\ : CascadeMux
    port map (
            O => \N__11116\,
            I => \N__11110\
        );

    \I__1434\ : CascadeBuf
    port map (
            O => \N__11113\,
            I => \N__11107\
        );

    \I__1433\ : CascadeBuf
    port map (
            O => \N__11110\,
            I => \N__11104\
        );

    \I__1432\ : CascadeMux
    port map (
            O => \N__11107\,
            I => \N__11101\
        );

    \I__1431\ : CascadeMux
    port map (
            O => \N__11104\,
            I => \N__11098\
        );

    \I__1430\ : CascadeBuf
    port map (
            O => \N__11101\,
            I => \N__11095\
        );

    \I__1429\ : CascadeBuf
    port map (
            O => \N__11098\,
            I => \N__11092\
        );

    \I__1428\ : CascadeMux
    port map (
            O => \N__11095\,
            I => \N__11089\
        );

    \I__1427\ : CascadeMux
    port map (
            O => \N__11092\,
            I => \N__11086\
        );

    \I__1426\ : CascadeBuf
    port map (
            O => \N__11089\,
            I => \N__11083\
        );

    \I__1425\ : CascadeBuf
    port map (
            O => \N__11086\,
            I => \N__11080\
        );

    \I__1424\ : CascadeMux
    port map (
            O => \N__11083\,
            I => \N__11077\
        );

    \I__1423\ : CascadeMux
    port map (
            O => \N__11080\,
            I => \N__11074\
        );

    \I__1422\ : CascadeBuf
    port map (
            O => \N__11077\,
            I => \N__11071\
        );

    \I__1421\ : CascadeBuf
    port map (
            O => \N__11074\,
            I => \N__11068\
        );

    \I__1420\ : CascadeMux
    port map (
            O => \N__11071\,
            I => \N__11065\
        );

    \I__1419\ : CascadeMux
    port map (
            O => \N__11068\,
            I => \N__11062\
        );

    \I__1418\ : CascadeBuf
    port map (
            O => \N__11065\,
            I => \N__11059\
        );

    \I__1417\ : InMux
    port map (
            O => \N__11062\,
            I => \N__11056\
        );

    \I__1416\ : CascadeMux
    port map (
            O => \N__11059\,
            I => \N__11053\
        );

    \I__1415\ : LocalMux
    port map (
            O => \N__11056\,
            I => \N__11050\
        );

    \I__1414\ : InMux
    port map (
            O => \N__11053\,
            I => \N__11047\
        );

    \I__1413\ : Span4Mux_s2_v
    port map (
            O => \N__11050\,
            I => \N__11044\
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__11047\,
            I => \N__11041\
        );

    \I__1411\ : Span4Mux_v
    port map (
            O => \N__11044\,
            I => \N__11038\
        );

    \I__1410\ : Sp12to4
    port map (
            O => \N__11041\,
            I => \N__11035\
        );

    \I__1409\ : Span4Mux_v
    port map (
            O => \N__11038\,
            I => \N__11032\
        );

    \I__1408\ : Span12Mux_s11_v
    port map (
            O => \N__11035\,
            I => \N__11029\
        );

    \I__1407\ : Span4Mux_v
    port map (
            O => \N__11032\,
            I => \N__11026\
        );

    \I__1406\ : Span12Mux_h
    port map (
            O => \N__11029\,
            I => \N__11023\
        );

    \I__1405\ : Span4Mux_h
    port map (
            O => \N__11026\,
            I => \N__11020\
        );

    \I__1404\ : Odrv12
    port map (
            O => \N__11023\,
            I => n21
        );

    \I__1403\ : Odrv4
    port map (
            O => \N__11020\,
            I => n21
        );

    \I__1402\ : InMux
    port map (
            O => \N__11015\,
            I => \N__11010\
        );

    \I__1401\ : InMux
    port map (
            O => \N__11014\,
            I => \N__11006\
        );

    \I__1400\ : InMux
    port map (
            O => \N__11013\,
            I => \N__11003\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__11010\,
            I => \N__11000\
        );

    \I__1398\ : InMux
    port map (
            O => \N__11009\,
            I => \N__10997\
        );

    \I__1397\ : LocalMux
    port map (
            O => \N__11006\,
            I => \transmit_module.video_signal_controller.VGA_Y_1\
        );

    \I__1396\ : LocalMux
    port map (
            O => \N__11003\,
            I => \transmit_module.video_signal_controller.VGA_Y_1\
        );

    \I__1395\ : Odrv4
    port map (
            O => \N__11000\,
            I => \transmit_module.video_signal_controller.VGA_Y_1\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__10997\,
            I => \transmit_module.video_signal_controller.VGA_Y_1\
        );

    \I__1393\ : InMux
    port map (
            O => \N__10988\,
            I => \N__10985\
        );

    \I__1392\ : LocalMux
    port map (
            O => \N__10985\,
            I => \N__10982\
        );

    \I__1391\ : Odrv4
    port map (
            O => \N__10982\,
            I => \transmit_module.video_signal_controller.n3520\
        );

    \I__1390\ : CascadeMux
    port map (
            O => \N__10979\,
            I => \N__10976\
        );

    \I__1389\ : InMux
    port map (
            O => \N__10976\,
            I => \N__10972\
        );

    \I__1388\ : InMux
    port map (
            O => \N__10975\,
            I => \N__10969\
        );

    \I__1387\ : LocalMux
    port map (
            O => \N__10972\,
            I => \transmit_module.video_signal_controller.VGA_Y_0\
        );

    \I__1386\ : LocalMux
    port map (
            O => \N__10969\,
            I => \transmit_module.video_signal_controller.VGA_Y_0\
        );

    \I__1385\ : InMux
    port map (
            O => \N__10964\,
            I => \N__10959\
        );

    \I__1384\ : InMux
    port map (
            O => \N__10963\,
            I => \N__10955\
        );

    \I__1383\ : InMux
    port map (
            O => \N__10962\,
            I => \N__10952\
        );

    \I__1382\ : LocalMux
    port map (
            O => \N__10959\,
            I => \N__10949\
        );

    \I__1381\ : InMux
    port map (
            O => \N__10958\,
            I => \N__10946\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__10955\,
            I => \transmit_module.video_signal_controller.VGA_Y_2\
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__10952\,
            I => \transmit_module.video_signal_controller.VGA_Y_2\
        );

    \I__1378\ : Odrv4
    port map (
            O => \N__10949\,
            I => \transmit_module.video_signal_controller.VGA_Y_2\
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__10946\,
            I => \transmit_module.video_signal_controller.VGA_Y_2\
        );

    \I__1376\ : CascadeMux
    port map (
            O => \N__10937\,
            I => \N__10934\
        );

    \I__1375\ : InMux
    port map (
            O => \N__10934\,
            I => \N__10931\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__10931\,
            I => \N__10928\
        );

    \I__1373\ : Odrv4
    port map (
            O => \N__10928\,
            I => \transmit_module.video_signal_controller.n2958\
        );

    \I__1372\ : CascadeMux
    port map (
            O => \N__10925\,
            I => \N__10922\
        );

    \I__1371\ : InMux
    port map (
            O => \N__10922\,
            I => \N__10919\
        );

    \I__1370\ : LocalMux
    port map (
            O => \N__10919\,
            I => \N__10916\
        );

    \I__1369\ : Span4Mux_h
    port map (
            O => \N__10916\,
            I => \N__10913\
        );

    \I__1368\ : Odrv4
    port map (
            O => \N__10913\,
            I => \transmit_module.video_signal_controller.n2975\
        );

    \I__1367\ : InMux
    port map (
            O => \N__10910\,
            I => \N__10907\
        );

    \I__1366\ : LocalMux
    port map (
            O => \N__10907\,
            I => \receive_module.rx_counter.n10\
        );

    \I__1365\ : CascadeMux
    port map (
            O => \N__10904\,
            I => \receive_module.rx_counter.n14_cascade_\
        );

    \I__1364\ : InMux
    port map (
            O => \N__10901\,
            I => \N__10898\
        );

    \I__1363\ : LocalMux
    port map (
            O => \N__10898\,
            I => \N__10895\
        );

    \I__1362\ : Span4Mux_v
    port map (
            O => \N__10895\,
            I => \N__10892\
        );

    \I__1361\ : Span4Mux_h
    port map (
            O => \N__10892\,
            I => \N__10889\
        );

    \I__1360\ : Odrv4
    port map (
            O => \N__10889\,
            I => \line_buffer.n539\
        );

    \I__1359\ : InMux
    port map (
            O => \N__10886\,
            I => \N__10883\
        );

    \I__1358\ : LocalMux
    port map (
            O => \N__10883\,
            I => \N__10880\
        );

    \I__1357\ : Span12Mux_v
    port map (
            O => \N__10880\,
            I => \N__10877\
        );

    \I__1356\ : Span12Mux_h
    port map (
            O => \N__10877\,
            I => \N__10874\
        );

    \I__1355\ : Odrv12
    port map (
            O => \N__10874\,
            I => \line_buffer.n531\
        );

    \I__1354\ : InMux
    port map (
            O => \N__10871\,
            I => \N__10865\
        );

    \I__1353\ : InMux
    port map (
            O => \N__10870\,
            I => \N__10865\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__10865\,
            I => \N__10862\
        );

    \I__1351\ : Span4Mux_h
    port map (
            O => \N__10862\,
            I => \N__10857\
        );

    \I__1350\ : InMux
    port map (
            O => \N__10861\,
            I => \N__10852\
        );

    \I__1349\ : InMux
    port map (
            O => \N__10860\,
            I => \N__10852\
        );

    \I__1348\ : Odrv4
    port map (
            O => \N__10857\,
            I => \transmit_module.old_VGA_HS\
        );

    \I__1347\ : LocalMux
    port map (
            O => \N__10852\,
            I => \transmit_module.old_VGA_HS\
        );

    \I__1346\ : InMux
    port map (
            O => \N__10847\,
            I => \N__10844\
        );

    \I__1345\ : LocalMux
    port map (
            O => \N__10844\,
            I => \N__10841\
        );

    \I__1344\ : Odrv4
    port map (
            O => \N__10841\,
            I => \transmit_module.ADDR_Y_COMPONENT_7\
        );

    \I__1343\ : InMux
    port map (
            O => \N__10838\,
            I => \N__10835\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__10835\,
            I => \N__10832\
        );

    \I__1341\ : Odrv4
    port map (
            O => \N__10832\,
            I => \transmit_module.video_signal_controller.n7\
        );

    \I__1340\ : IoInMux
    port map (
            O => \N__10829\,
            I => \N__10826\
        );

    \I__1339\ : LocalMux
    port map (
            O => \N__10826\,
            I => \N__10823\
        );

    \I__1338\ : IoSpan4Mux
    port map (
            O => \N__10823\,
            I => \N__10820\
        );

    \I__1337\ : Sp12to4
    port map (
            O => \N__10820\,
            I => \N__10815\
        );

    \I__1336\ : InMux
    port map (
            O => \N__10819\,
            I => \N__10810\
        );

    \I__1335\ : InMux
    port map (
            O => \N__10818\,
            I => \N__10810\
        );

    \I__1334\ : Span12Mux_h
    port map (
            O => \N__10815\,
            I => \N__10804\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__10810\,
            I => \N__10801\
        );

    \I__1332\ : InMux
    port map (
            O => \N__10809\,
            I => \N__10794\
        );

    \I__1331\ : InMux
    port map (
            O => \N__10808\,
            I => \N__10794\
        );

    \I__1330\ : InMux
    port map (
            O => \N__10807\,
            I => \N__10794\
        );

    \I__1329\ : Odrv12
    port map (
            O => \N__10804\,
            I => \ADV_HSYNC_c\
        );

    \I__1328\ : Odrv4
    port map (
            O => \N__10801\,
            I => \ADV_HSYNC_c\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__10794\,
            I => \ADV_HSYNC_c\
        );

    \I__1326\ : InMux
    port map (
            O => \N__10787\,
            I => \receive_module.rx_counter.n3175\
        );

    \I__1325\ : InMux
    port map (
            O => \N__10784\,
            I => \receive_module.rx_counter.n3176\
        );

    \I__1324\ : InMux
    port map (
            O => \N__10781\,
            I => \receive_module.rx_counter.n3177\
        );

    \I__1323\ : InMux
    port map (
            O => \N__10778\,
            I => \receive_module.rx_counter.n3178\
        );

    \I__1322\ : InMux
    port map (
            O => \N__10775\,
            I => \receive_module.rx_counter.n3179\
        );

    \I__1321\ : InMux
    port map (
            O => \N__10772\,
            I => \receive_module.rx_counter.n3180\
        );

    \I__1320\ : InMux
    port map (
            O => \N__10769\,
            I => \receive_module.rx_counter.n3181\
        );

    \I__1319\ : InMux
    port map (
            O => \N__10766\,
            I => \bfn_13_12_0_\
        );

    \I__1318\ : InMux
    port map (
            O => \N__10763\,
            I => \receive_module.rx_counter.n3211\
        );

    \I__1317\ : InMux
    port map (
            O => \N__10760\,
            I => \receive_module.rx_counter.n3212\
        );

    \I__1316\ : InMux
    port map (
            O => \N__10757\,
            I => \receive_module.rx_counter.n3213\
        );

    \I__1315\ : InMux
    port map (
            O => \N__10754\,
            I => \receive_module.rx_counter.n3214\
        );

    \I__1314\ : InMux
    port map (
            O => \N__10751\,
            I => \receive_module.rx_counter.n3215\
        );

    \I__1313\ : InMux
    port map (
            O => \N__10748\,
            I => \receive_module.rx_counter.n3216\
        );

    \I__1312\ : InMux
    port map (
            O => \N__10745\,
            I => \bfn_13_10_0_\
        );

    \I__1311\ : InMux
    port map (
            O => \N__10742\,
            I => \receive_module.rx_counter.n3218\
        );

    \I__1310\ : InMux
    port map (
            O => \N__10739\,
            I => \bfn_13_11_0_\
        );

    \I__1309\ : InMux
    port map (
            O => \N__10736\,
            I => \N__10732\
        );

    \I__1308\ : InMux
    port map (
            O => \N__10735\,
            I => \N__10729\
        );

    \I__1307\ : LocalMux
    port map (
            O => \N__10732\,
            I => \N__10725\
        );

    \I__1306\ : LocalMux
    port map (
            O => \N__10729\,
            I => \N__10721\
        );

    \I__1305\ : InMux
    port map (
            O => \N__10728\,
            I => \N__10718\
        );

    \I__1304\ : Span4Mux_v
    port map (
            O => \N__10725\,
            I => \N__10712\
        );

    \I__1303\ : InMux
    port map (
            O => \N__10724\,
            I => \N__10709\
        );

    \I__1302\ : Sp12to4
    port map (
            O => \N__10721\,
            I => \N__10703\
        );

    \I__1301\ : LocalMux
    port map (
            O => \N__10718\,
            I => \N__10703\
        );

    \I__1300\ : InMux
    port map (
            O => \N__10717\,
            I => \N__10700\
        );

    \I__1299\ : InMux
    port map (
            O => \N__10716\,
            I => \N__10697\
        );

    \I__1298\ : InMux
    port map (
            O => \N__10715\,
            I => \N__10694\
        );

    \I__1297\ : Span4Mux_v
    port map (
            O => \N__10712\,
            I => \N__10689\
        );

    \I__1296\ : LocalMux
    port map (
            O => \N__10709\,
            I => \N__10689\
        );

    \I__1295\ : InMux
    port map (
            O => \N__10708\,
            I => \N__10686\
        );

    \I__1294\ : Span12Mux_s9_v
    port map (
            O => \N__10703\,
            I => \N__10679\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__10700\,
            I => \N__10679\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__10697\,
            I => \N__10679\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__10694\,
            I => \N__10676\
        );

    \I__1290\ : Span4Mux_v
    port map (
            O => \N__10689\,
            I => \N__10673\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__10686\,
            I => \N__10670\
        );

    \I__1288\ : Span12Mux_v
    port map (
            O => \N__10679\,
            I => \N__10665\
        );

    \I__1287\ : Span12Mux_s10_v
    port map (
            O => \N__10676\,
            I => \N__10665\
        );

    \I__1286\ : Span4Mux_v
    port map (
            O => \N__10673\,
            I => \N__10660\
        );

    \I__1285\ : Span4Mux_h
    port map (
            O => \N__10670\,
            I => \N__10660\
        );

    \I__1284\ : Span12Mux_h
    port map (
            O => \N__10665\,
            I => \N__10657\
        );

    \I__1283\ : Span4Mux_h
    port map (
            O => \N__10660\,
            I => \N__10654\
        );

    \I__1282\ : Odrv12
    port map (
            O => \N__10657\,
            I => \RX_DATA_0\
        );

    \I__1281\ : Odrv4
    port map (
            O => \N__10654\,
            I => \RX_DATA_0\
        );

    \I__1280\ : InMux
    port map (
            O => \N__10649\,
            I => \N__10646\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__10646\,
            I => \N__10643\
        );

    \I__1278\ : Span4Mux_h
    port map (
            O => \N__10643\,
            I => \N__10640\
        );

    \I__1277\ : Span4Mux_v
    port map (
            O => \N__10640\,
            I => \N__10637\
        );

    \I__1276\ : Odrv4
    port map (
            O => \N__10637\,
            I => \TVP_VIDEO_c_4\
        );

    \I__1275\ : InMux
    port map (
            O => \N__10634\,
            I => \N__10631\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__10631\,
            I => \tvp_video_buffer.BUFFER_0_4\
        );

    \I__1273\ : InMux
    port map (
            O => \N__10628\,
            I => \N__10625\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__10625\,
            I => \N__10622\
        );

    \I__1271\ : Span12Mux_h
    port map (
            O => \N__10622\,
            I => \N__10619\
        );

    \I__1270\ : Odrv12
    port map (
            O => \N__10619\,
            I => \TVP_VIDEO_c_8\
        );

    \I__1269\ : InMux
    port map (
            O => \N__10616\,
            I => \N__10613\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__10613\,
            I => \tvp_video_buffer.BUFFER_1_3\
        );

    \I__1267\ : InMux
    port map (
            O => \N__10610\,
            I => \N__10606\
        );

    \I__1266\ : InMux
    port map (
            O => \N__10609\,
            I => \N__10603\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__10606\,
            I => \N__10596\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__10603\,
            I => \N__10591\
        );

    \I__1263\ : InMux
    port map (
            O => \N__10602\,
            I => \N__10588\
        );

    \I__1262\ : InMux
    port map (
            O => \N__10601\,
            I => \N__10585\
        );

    \I__1261\ : InMux
    port map (
            O => \N__10600\,
            I => \N__10582\
        );

    \I__1260\ : InMux
    port map (
            O => \N__10599\,
            I => \N__10579\
        );

    \I__1259\ : Span4Mux_v
    port map (
            O => \N__10596\,
            I => \N__10576\
        );

    \I__1258\ : InMux
    port map (
            O => \N__10595\,
            I => \N__10573\
        );

    \I__1257\ : InMux
    port map (
            O => \N__10594\,
            I => \N__10570\
        );

    \I__1256\ : Sp12to4
    port map (
            O => \N__10591\,
            I => \N__10565\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__10588\,
            I => \N__10565\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__10585\,
            I => \N__10560\
        );

    \I__1253\ : LocalMux
    port map (
            O => \N__10582\,
            I => \N__10560\
        );

    \I__1252\ : LocalMux
    port map (
            O => \N__10579\,
            I => \N__10557\
        );

    \I__1251\ : Span4Mux_v
    port map (
            O => \N__10576\,
            I => \N__10552\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__10573\,
            I => \N__10552\
        );

    \I__1249\ : LocalMux
    port map (
            O => \N__10570\,
            I => \N__10549\
        );

    \I__1248\ : Span12Mux_v
    port map (
            O => \N__10565\,
            I => \N__10546\
        );

    \I__1247\ : Span12Mux_v
    port map (
            O => \N__10560\,
            I => \N__10541\
        );

    \I__1246\ : Span12Mux_s5_v
    port map (
            O => \N__10557\,
            I => \N__10541\
        );

    \I__1245\ : Span4Mux_v
    port map (
            O => \N__10552\,
            I => \N__10536\
        );

    \I__1244\ : Span4Mux_v
    port map (
            O => \N__10549\,
            I => \N__10536\
        );

    \I__1243\ : Span12Mux_h
    port map (
            O => \N__10546\,
            I => \N__10531\
        );

    \I__1242\ : Span12Mux_h
    port map (
            O => \N__10541\,
            I => \N__10531\
        );

    \I__1241\ : Span4Mux_h
    port map (
            O => \N__10536\,
            I => \N__10528\
        );

    \I__1240\ : Odrv12
    port map (
            O => \N__10531\,
            I => \RX_DATA_1\
        );

    \I__1239\ : Odrv4
    port map (
            O => \N__10528\,
            I => \RX_DATA_1\
        );

    \I__1238\ : InMux
    port map (
            O => \N__10523\,
            I => \N__10520\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__10520\,
            I => \tvp_video_buffer.BUFFER_1_4\
        );

    \I__1236\ : InMux
    port map (
            O => \N__10517\,
            I => \N__10514\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__10514\,
            I => \N__10510\
        );

    \I__1234\ : InMux
    port map (
            O => \N__10513\,
            I => \N__10507\
        );

    \I__1233\ : Span4Mux_s2_v
    port map (
            O => \N__10510\,
            I => \N__10504\
        );

    \I__1232\ : LocalMux
    port map (
            O => \N__10507\,
            I => \N__10501\
        );

    \I__1231\ : Span4Mux_v
    port map (
            O => \N__10504\,
            I => \N__10497\
        );

    \I__1230\ : Span4Mux_v
    port map (
            O => \N__10501\,
            I => \N__10493\
        );

    \I__1229\ : InMux
    port map (
            O => \N__10500\,
            I => \N__10490\
        );

    \I__1228\ : Span4Mux_v
    port map (
            O => \N__10497\,
            I => \N__10486\
        );

    \I__1227\ : InMux
    port map (
            O => \N__10496\,
            I => \N__10483\
        );

    \I__1226\ : Span4Mux_v
    port map (
            O => \N__10493\,
            I => \N__10477\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__10490\,
            I => \N__10477\
        );

    \I__1224\ : InMux
    port map (
            O => \N__10489\,
            I => \N__10472\
        );

    \I__1223\ : Span4Mux_v
    port map (
            O => \N__10486\,
            I => \N__10467\
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__10483\,
            I => \N__10467\
        );

    \I__1221\ : InMux
    port map (
            O => \N__10482\,
            I => \N__10464\
        );

    \I__1220\ : Span4Mux_v
    port map (
            O => \N__10477\,
            I => \N__10461\
        );

    \I__1219\ : InMux
    port map (
            O => \N__10476\,
            I => \N__10458\
        );

    \I__1218\ : InMux
    port map (
            O => \N__10475\,
            I => \N__10455\
        );

    \I__1217\ : LocalMux
    port map (
            O => \N__10472\,
            I => \N__10452\
        );

    \I__1216\ : Span4Mux_v
    port map (
            O => \N__10467\,
            I => \N__10449\
        );

    \I__1215\ : LocalMux
    port map (
            O => \N__10464\,
            I => \N__10446\
        );

    \I__1214\ : Sp12to4
    port map (
            O => \N__10461\,
            I => \N__10439\
        );

    \I__1213\ : LocalMux
    port map (
            O => \N__10458\,
            I => \N__10439\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__10455\,
            I => \N__10439\
        );

    \I__1211\ : Span4Mux_v
    port map (
            O => \N__10452\,
            I => \N__10436\
        );

    \I__1210\ : Span4Mux_v
    port map (
            O => \N__10449\,
            I => \N__10431\
        );

    \I__1209\ : Span4Mux_h
    port map (
            O => \N__10446\,
            I => \N__10431\
        );

    \I__1208\ : Span12Mux_v
    port map (
            O => \N__10439\,
            I => \N__10428\
        );

    \I__1207\ : Span4Mux_h
    port map (
            O => \N__10436\,
            I => \N__10423\
        );

    \I__1206\ : Span4Mux_h
    port map (
            O => \N__10431\,
            I => \N__10423\
        );

    \I__1205\ : Odrv12
    port map (
            O => \N__10428\,
            I => \RX_DATA_2\
        );

    \I__1204\ : Odrv4
    port map (
            O => \N__10423\,
            I => \RX_DATA_2\
        );

    \I__1203\ : InMux
    port map (
            O => \N__10418\,
            I => \N__10415\
        );

    \I__1202\ : LocalMux
    port map (
            O => \N__10415\,
            I => \tvp_video_buffer.BUFFER_0_8\
        );

    \I__1201\ : InMux
    port map (
            O => \N__10412\,
            I => \N__10409\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__10409\,
            I => \tvp_video_buffer.BUFFER_1_8\
        );

    \I__1199\ : InMux
    port map (
            O => \N__10406\,
            I => \bfn_13_9_0_\
        );

    \I__1198\ : InMux
    port map (
            O => \N__10403\,
            I => \receive_module.rx_counter.n3210\
        );

    \I__1197\ : CascadeMux
    port map (
            O => \N__10400\,
            I => \N__10396\
        );

    \I__1196\ : InMux
    port map (
            O => \N__10399\,
            I => \N__10391\
        );

    \I__1195\ : InMux
    port map (
            O => \N__10396\,
            I => \N__10384\
        );

    \I__1194\ : InMux
    port map (
            O => \N__10395\,
            I => \N__10384\
        );

    \I__1193\ : InMux
    port map (
            O => \N__10394\,
            I => \N__10384\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__10391\,
            I => \transmit_module.video_signal_controller.VGA_X_3\
        );

    \I__1191\ : LocalMux
    port map (
            O => \N__10384\,
            I => \transmit_module.video_signal_controller.VGA_X_3\
        );

    \I__1190\ : InMux
    port map (
            O => \N__10379\,
            I => \N__10373\
        );

    \I__1189\ : InMux
    port map (
            O => \N__10378\,
            I => \N__10366\
        );

    \I__1188\ : InMux
    port map (
            O => \N__10377\,
            I => \N__10366\
        );

    \I__1187\ : InMux
    port map (
            O => \N__10376\,
            I => \N__10366\
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__10373\,
            I => \transmit_module.video_signal_controller.VGA_X_4\
        );

    \I__1185\ : LocalMux
    port map (
            O => \N__10366\,
            I => \transmit_module.video_signal_controller.VGA_X_4\
        );

    \I__1184\ : InMux
    port map (
            O => \N__10361\,
            I => \N__10358\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__10358\,
            I => \N__10352\
        );

    \I__1182\ : InMux
    port map (
            O => \N__10357\,
            I => \N__10349\
        );

    \I__1181\ : InMux
    port map (
            O => \N__10356\,
            I => \N__10344\
        );

    \I__1180\ : InMux
    port map (
            O => \N__10355\,
            I => \N__10344\
        );

    \I__1179\ : Span4Mux_h
    port map (
            O => \N__10352\,
            I => \N__10341\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__10349\,
            I => \transmit_module.video_signal_controller.VGA_X_6\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__10344\,
            I => \transmit_module.video_signal_controller.VGA_X_6\
        );

    \I__1176\ : Odrv4
    port map (
            O => \N__10341\,
            I => \transmit_module.video_signal_controller.VGA_X_6\
        );

    \I__1175\ : CascadeMux
    port map (
            O => \N__10334\,
            I => \transmit_module.video_signal_controller.n3482_cascade_\
        );

    \I__1174\ : InMux
    port map (
            O => \N__10331\,
            I => \N__10328\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__10328\,
            I => \N__10322\
        );

    \I__1172\ : InMux
    port map (
            O => \N__10327\,
            I => \N__10319\
        );

    \I__1171\ : InMux
    port map (
            O => \N__10326\,
            I => \N__10314\
        );

    \I__1170\ : InMux
    port map (
            O => \N__10325\,
            I => \N__10314\
        );

    \I__1169\ : Span4Mux_h
    port map (
            O => \N__10322\,
            I => \N__10311\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__10319\,
            I => \transmit_module.video_signal_controller.VGA_X_5\
        );

    \I__1167\ : LocalMux
    port map (
            O => \N__10314\,
            I => \transmit_module.video_signal_controller.VGA_X_5\
        );

    \I__1166\ : Odrv4
    port map (
            O => \N__10311\,
            I => \transmit_module.video_signal_controller.VGA_X_5\
        );

    \I__1165\ : InMux
    port map (
            O => \N__10304\,
            I => \N__10301\
        );

    \I__1164\ : LocalMux
    port map (
            O => \N__10301\,
            I => \transmit_module.video_signal_controller.n55\
        );

    \I__1163\ : CascadeMux
    port map (
            O => \N__10298\,
            I => \transmit_module.video_signal_controller.n3478_cascade_\
        );

    \I__1162\ : InMux
    port map (
            O => \N__10295\,
            I => \N__10290\
        );

    \I__1161\ : InMux
    port map (
            O => \N__10294\,
            I => \N__10287\
        );

    \I__1160\ : InMux
    port map (
            O => \N__10293\,
            I => \N__10284\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__10290\,
            I => \transmit_module.video_signal_controller.VGA_X_7\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__10287\,
            I => \transmit_module.video_signal_controller.VGA_X_7\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__10284\,
            I => \transmit_module.video_signal_controller.VGA_X_7\
        );

    \I__1156\ : CascadeMux
    port map (
            O => \N__10277\,
            I => \N__10272\
        );

    \I__1155\ : InMux
    port map (
            O => \N__10276\,
            I => \N__10269\
        );

    \I__1154\ : InMux
    port map (
            O => \N__10275\,
            I => \N__10264\
        );

    \I__1153\ : InMux
    port map (
            O => \N__10272\,
            I => \N__10264\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__10269\,
            I => \transmit_module.video_signal_controller.VGA_X_0\
        );

    \I__1151\ : LocalMux
    port map (
            O => \N__10264\,
            I => \transmit_module.video_signal_controller.VGA_X_0\
        );

    \I__1150\ : InMux
    port map (
            O => \N__10259\,
            I => \N__10256\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__10256\,
            I => \N__10253\
        );

    \I__1148\ : Span4Mux_h
    port map (
            O => \N__10253\,
            I => \N__10250\
        );

    \I__1147\ : Odrv4
    port map (
            O => \N__10250\,
            I => \transmit_module.ADDR_Y_COMPONENT_13\
        );

    \I__1146\ : CEMux
    port map (
            O => \N__10247\,
            I => \N__10243\
        );

    \I__1145\ : CEMux
    port map (
            O => \N__10246\,
            I => \N__10240\
        );

    \I__1144\ : LocalMux
    port map (
            O => \N__10243\,
            I => \N__10237\
        );

    \I__1143\ : LocalMux
    port map (
            O => \N__10240\,
            I => \N__10234\
        );

    \I__1142\ : Span4Mux_v
    port map (
            O => \N__10237\,
            I => \N__10231\
        );

    \I__1141\ : Span4Mux_h
    port map (
            O => \N__10234\,
            I => \N__10228\
        );

    \I__1140\ : Span4Mux_h
    port map (
            O => \N__10231\,
            I => \N__10225\
        );

    \I__1139\ : Odrv4
    port map (
            O => \N__10228\,
            I => \transmit_module.n2073\
        );

    \I__1138\ : Odrv4
    port map (
            O => \N__10225\,
            I => \transmit_module.n2073\
        );

    \I__1137\ : CascadeMux
    port map (
            O => \N__10220\,
            I => \N__10216\
        );

    \I__1136\ : CascadeMux
    port map (
            O => \N__10219\,
            I => \N__10213\
        );

    \I__1135\ : CascadeBuf
    port map (
            O => \N__10216\,
            I => \N__10210\
        );

    \I__1134\ : CascadeBuf
    port map (
            O => \N__10213\,
            I => \N__10207\
        );

    \I__1133\ : CascadeMux
    port map (
            O => \N__10210\,
            I => \N__10204\
        );

    \I__1132\ : CascadeMux
    port map (
            O => \N__10207\,
            I => \N__10201\
        );

    \I__1131\ : CascadeBuf
    port map (
            O => \N__10204\,
            I => \N__10198\
        );

    \I__1130\ : CascadeBuf
    port map (
            O => \N__10201\,
            I => \N__10195\
        );

    \I__1129\ : CascadeMux
    port map (
            O => \N__10198\,
            I => \N__10192\
        );

    \I__1128\ : CascadeMux
    port map (
            O => \N__10195\,
            I => \N__10189\
        );

    \I__1127\ : CascadeBuf
    port map (
            O => \N__10192\,
            I => \N__10186\
        );

    \I__1126\ : CascadeBuf
    port map (
            O => \N__10189\,
            I => \N__10183\
        );

    \I__1125\ : CascadeMux
    port map (
            O => \N__10186\,
            I => \N__10180\
        );

    \I__1124\ : CascadeMux
    port map (
            O => \N__10183\,
            I => \N__10177\
        );

    \I__1123\ : CascadeBuf
    port map (
            O => \N__10180\,
            I => \N__10174\
        );

    \I__1122\ : CascadeBuf
    port map (
            O => \N__10177\,
            I => \N__10171\
        );

    \I__1121\ : CascadeMux
    port map (
            O => \N__10174\,
            I => \N__10168\
        );

    \I__1120\ : CascadeMux
    port map (
            O => \N__10171\,
            I => \N__10165\
        );

    \I__1119\ : CascadeBuf
    port map (
            O => \N__10168\,
            I => \N__10162\
        );

    \I__1118\ : CascadeBuf
    port map (
            O => \N__10165\,
            I => \N__10159\
        );

    \I__1117\ : CascadeMux
    port map (
            O => \N__10162\,
            I => \N__10156\
        );

    \I__1116\ : CascadeMux
    port map (
            O => \N__10159\,
            I => \N__10153\
        );

    \I__1115\ : CascadeBuf
    port map (
            O => \N__10156\,
            I => \N__10150\
        );

    \I__1114\ : CascadeBuf
    port map (
            O => \N__10153\,
            I => \N__10147\
        );

    \I__1113\ : CascadeMux
    port map (
            O => \N__10150\,
            I => \N__10144\
        );

    \I__1112\ : CascadeMux
    port map (
            O => \N__10147\,
            I => \N__10141\
        );

    \I__1111\ : CascadeBuf
    port map (
            O => \N__10144\,
            I => \N__10138\
        );

    \I__1110\ : CascadeBuf
    port map (
            O => \N__10141\,
            I => \N__10135\
        );

    \I__1109\ : CascadeMux
    port map (
            O => \N__10138\,
            I => \N__10132\
        );

    \I__1108\ : CascadeMux
    port map (
            O => \N__10135\,
            I => \N__10129\
        );

    \I__1107\ : CascadeBuf
    port map (
            O => \N__10132\,
            I => \N__10126\
        );

    \I__1106\ : CascadeBuf
    port map (
            O => \N__10129\,
            I => \N__10123\
        );

    \I__1105\ : CascadeMux
    port map (
            O => \N__10126\,
            I => \N__10120\
        );

    \I__1104\ : CascadeMux
    port map (
            O => \N__10123\,
            I => \N__10117\
        );

    \I__1103\ : CascadeBuf
    port map (
            O => \N__10120\,
            I => \N__10114\
        );

    \I__1102\ : CascadeBuf
    port map (
            O => \N__10117\,
            I => \N__10111\
        );

    \I__1101\ : CascadeMux
    port map (
            O => \N__10114\,
            I => \N__10108\
        );

    \I__1100\ : CascadeMux
    port map (
            O => \N__10111\,
            I => \N__10105\
        );

    \I__1099\ : CascadeBuf
    port map (
            O => \N__10108\,
            I => \N__10102\
        );

    \I__1098\ : CascadeBuf
    port map (
            O => \N__10105\,
            I => \N__10099\
        );

    \I__1097\ : CascadeMux
    port map (
            O => \N__10102\,
            I => \N__10096\
        );

    \I__1096\ : CascadeMux
    port map (
            O => \N__10099\,
            I => \N__10093\
        );

    \I__1095\ : CascadeBuf
    port map (
            O => \N__10096\,
            I => \N__10090\
        );

    \I__1094\ : CascadeBuf
    port map (
            O => \N__10093\,
            I => \N__10087\
        );

    \I__1093\ : CascadeMux
    port map (
            O => \N__10090\,
            I => \N__10084\
        );

    \I__1092\ : CascadeMux
    port map (
            O => \N__10087\,
            I => \N__10081\
        );

    \I__1091\ : CascadeBuf
    port map (
            O => \N__10084\,
            I => \N__10078\
        );

    \I__1090\ : CascadeBuf
    port map (
            O => \N__10081\,
            I => \N__10075\
        );

    \I__1089\ : CascadeMux
    port map (
            O => \N__10078\,
            I => \N__10072\
        );

    \I__1088\ : CascadeMux
    port map (
            O => \N__10075\,
            I => \N__10069\
        );

    \I__1087\ : CascadeBuf
    port map (
            O => \N__10072\,
            I => \N__10066\
        );

    \I__1086\ : CascadeBuf
    port map (
            O => \N__10069\,
            I => \N__10063\
        );

    \I__1085\ : CascadeMux
    port map (
            O => \N__10066\,
            I => \N__10060\
        );

    \I__1084\ : CascadeMux
    port map (
            O => \N__10063\,
            I => \N__10057\
        );

    \I__1083\ : CascadeBuf
    port map (
            O => \N__10060\,
            I => \N__10054\
        );

    \I__1082\ : CascadeBuf
    port map (
            O => \N__10057\,
            I => \N__10051\
        );

    \I__1081\ : CascadeMux
    port map (
            O => \N__10054\,
            I => \N__10048\
        );

    \I__1080\ : CascadeMux
    port map (
            O => \N__10051\,
            I => \N__10045\
        );

    \I__1079\ : CascadeBuf
    port map (
            O => \N__10048\,
            I => \N__10042\
        );

    \I__1078\ : CascadeBuf
    port map (
            O => \N__10045\,
            I => \N__10039\
        );

    \I__1077\ : CascadeMux
    port map (
            O => \N__10042\,
            I => \N__10036\
        );

    \I__1076\ : CascadeMux
    port map (
            O => \N__10039\,
            I => \N__10033\
        );

    \I__1075\ : InMux
    port map (
            O => \N__10036\,
            I => \N__10030\
        );

    \I__1074\ : InMux
    port map (
            O => \N__10033\,
            I => \N__10027\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__10030\,
            I => \N__10024\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__10027\,
            I => \N__10021\
        );

    \I__1071\ : Span4Mux_v
    port map (
            O => \N__10024\,
            I => \N__10018\
        );

    \I__1070\ : Span12Mux_v
    port map (
            O => \N__10021\,
            I => \N__10015\
        );

    \I__1069\ : Span4Mux_v
    port map (
            O => \N__10018\,
            I => \N__10012\
        );

    \I__1068\ : Span12Mux_h
    port map (
            O => \N__10015\,
            I => \N__10009\
        );

    \I__1067\ : Span4Mux_v
    port map (
            O => \N__10012\,
            I => \N__10006\
        );

    \I__1066\ : Odrv12
    port map (
            O => \N__10009\,
            I => n20
        );

    \I__1065\ : Odrv4
    port map (
            O => \N__10006\,
            I => n20
        );

    \I__1064\ : InMux
    port map (
            O => \N__10001\,
            I => \N__9998\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__9998\,
            I => \N__9995\
        );

    \I__1062\ : Span4Mux_h
    port map (
            O => \N__9995\,
            I => \N__9992\
        );

    \I__1061\ : Odrv4
    port map (
            O => \N__9992\,
            I => \tvp_video_buffer.BUFFER_1_2\
        );

    \I__1060\ : InMux
    port map (
            O => \N__9989\,
            I => \N__9985\
        );

    \I__1059\ : InMux
    port map (
            O => \N__9988\,
            I => \N__9981\
        );

    \I__1058\ : LocalMux
    port map (
            O => \N__9985\,
            I => \N__9978\
        );

    \I__1057\ : InMux
    port map (
            O => \N__9984\,
            I => \N__9975\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__9981\,
            I => \transmit_module.video_signal_controller.VGA_Y_5\
        );

    \I__1055\ : Odrv4
    port map (
            O => \N__9978\,
            I => \transmit_module.video_signal_controller.VGA_Y_5\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__9975\,
            I => \transmit_module.video_signal_controller.VGA_Y_5\
        );

    \I__1053\ : CascadeMux
    port map (
            O => \N__9968\,
            I => \transmit_module.video_signal_controller.n3485_cascade_\
        );

    \I__1052\ : InMux
    port map (
            O => \N__9965\,
            I => \N__9961\
        );

    \I__1051\ : InMux
    port map (
            O => \N__9964\,
            I => \N__9957\
        );

    \I__1050\ : LocalMux
    port map (
            O => \N__9961\,
            I => \N__9954\
        );

    \I__1049\ : InMux
    port map (
            O => \N__9960\,
            I => \N__9951\
        );

    \I__1048\ : LocalMux
    port map (
            O => \N__9957\,
            I => \transmit_module.video_signal_controller.VGA_Y_6\
        );

    \I__1047\ : Odrv4
    port map (
            O => \N__9954\,
            I => \transmit_module.video_signal_controller.VGA_Y_6\
        );

    \I__1046\ : LocalMux
    port map (
            O => \N__9951\,
            I => \transmit_module.video_signal_controller.VGA_Y_6\
        );

    \I__1045\ : InMux
    port map (
            O => \N__9944\,
            I => \N__9941\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__9941\,
            I => \transmit_module.video_signal_controller.n3676\
        );

    \I__1043\ : InMux
    port map (
            O => \N__9938\,
            I => \N__9933\
        );

    \I__1042\ : InMux
    port map (
            O => \N__9937\,
            I => \N__9930\
        );

    \I__1041\ : InMux
    port map (
            O => \N__9936\,
            I => \N__9927\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__9933\,
            I => \transmit_module.video_signal_controller.VGA_Y_9\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__9930\,
            I => \transmit_module.video_signal_controller.VGA_Y_9\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__9927\,
            I => \transmit_module.video_signal_controller.VGA_Y_9\
        );

    \I__1037\ : CascadeMux
    port map (
            O => \N__9920\,
            I => \transmit_module.video_signal_controller.n3464_cascade_\
        );

    \I__1036\ : InMux
    port map (
            O => \N__9917\,
            I => \N__9913\
        );

    \I__1035\ : InMux
    port map (
            O => \N__9916\,
            I => \N__9910\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__9913\,
            I => \transmit_module.video_signal_controller.n3378\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__9910\,
            I => \transmit_module.video_signal_controller.n3378\
        );

    \I__1032\ : InMux
    port map (
            O => \N__9905\,
            I => \N__9902\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__9902\,
            I => \N__9899\
        );

    \I__1030\ : Odrv4
    port map (
            O => \N__9899\,
            I => \transmit_module.ADDR_Y_COMPONENT_5\
        );

    \I__1029\ : InMux
    port map (
            O => \N__9896\,
            I => \N__9888\
        );

    \I__1028\ : InMux
    port map (
            O => \N__9895\,
            I => \N__9888\
        );

    \I__1027\ : InMux
    port map (
            O => \N__9894\,
            I => \N__9885\
        );

    \I__1026\ : InMux
    port map (
            O => \N__9893\,
            I => \N__9882\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__9888\,
            I => \N__9879\
        );

    \I__1024\ : LocalMux
    port map (
            O => \N__9885\,
            I => \transmit_module.video_signal_controller.VGA_Y_3\
        );

    \I__1023\ : LocalMux
    port map (
            O => \N__9882\,
            I => \transmit_module.video_signal_controller.VGA_Y_3\
        );

    \I__1022\ : Odrv4
    port map (
            O => \N__9879\,
            I => \transmit_module.video_signal_controller.VGA_Y_3\
        );

    \I__1021\ : InMux
    port map (
            O => \N__9872\,
            I => \N__9869\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__9869\,
            I => \transmit_module.video_signal_controller.n6_adj_622\
        );

    \I__1019\ : CascadeMux
    port map (
            O => \N__9866\,
            I => \N__9862\
        );

    \I__1018\ : InMux
    port map (
            O => \N__9865\,
            I => \N__9855\
        );

    \I__1017\ : InMux
    port map (
            O => \N__9862\,
            I => \N__9855\
        );

    \I__1016\ : InMux
    port map (
            O => \N__9861\,
            I => \N__9852\
        );

    \I__1015\ : InMux
    port map (
            O => \N__9860\,
            I => \N__9849\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__9855\,
            I => \N__9846\
        );

    \I__1013\ : LocalMux
    port map (
            O => \N__9852\,
            I => \transmit_module.video_signal_controller.VGA_Y_4\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__9849\,
            I => \transmit_module.video_signal_controller.VGA_Y_4\
        );

    \I__1011\ : Odrv4
    port map (
            O => \N__9846\,
            I => \transmit_module.video_signal_controller.VGA_Y_4\
        );

    \I__1010\ : InMux
    port map (
            O => \N__9839\,
            I => \N__9835\
        );

    \I__1009\ : InMux
    port map (
            O => \N__9838\,
            I => \N__9832\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__9835\,
            I => \N__9829\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__9832\,
            I => \transmit_module.video_signal_controller.n2019\
        );

    \I__1006\ : Odrv4
    port map (
            O => \N__9829\,
            I => \transmit_module.video_signal_controller.n2019\
        );

    \I__1005\ : CEMux
    port map (
            O => \N__9824\,
            I => \N__9819\
        );

    \I__1004\ : SRMux
    port map (
            O => \N__9823\,
            I => \N__9815\
        );

    \I__1003\ : SRMux
    port map (
            O => \N__9822\,
            I => \N__9812\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__9819\,
            I => \N__9809\
        );

    \I__1001\ : CEMux
    port map (
            O => \N__9818\,
            I => \N__9806\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__9815\,
            I => \N__9803\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__9812\,
            I => \N__9800\
        );

    \I__998\ : Span4Mux_v
    port map (
            O => \N__9809\,
            I => \N__9793\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__9806\,
            I => \N__9793\
        );

    \I__996\ : Span4Mux_h
    port map (
            O => \N__9803\,
            I => \N__9793\
        );

    \I__995\ : Sp12to4
    port map (
            O => \N__9800\,
            I => \N__9790\
        );

    \I__994\ : Odrv4
    port map (
            O => \N__9793\,
            I => \transmit_module.video_signal_controller.n2050\
        );

    \I__993\ : Odrv12
    port map (
            O => \N__9790\,
            I => \transmit_module.video_signal_controller.n2050\
        );

    \I__992\ : CascadeMux
    port map (
            O => \N__9785\,
            I => \transmit_module.video_signal_controller.n2050_cascade_\
        );

    \I__991\ : SRMux
    port map (
            O => \N__9782\,
            I => \N__9779\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__9779\,
            I => \N__9775\
        );

    \I__989\ : SRMux
    port map (
            O => \N__9778\,
            I => \N__9772\
        );

    \I__988\ : Span4Mux_v
    port map (
            O => \N__9775\,
            I => \N__9767\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__9772\,
            I => \N__9767\
        );

    \I__986\ : Odrv4
    port map (
            O => \N__9767\,
            I => \transmit_module.video_signal_controller.n2398\
        );

    \I__985\ : InMux
    port map (
            O => \N__9764\,
            I => \transmit_module.video_signal_controller.n3197\
        );

    \I__984\ : InMux
    port map (
            O => \N__9761\,
            I => \transmit_module.video_signal_controller.n3198\
        );

    \I__983\ : InMux
    port map (
            O => \N__9758\,
            I => \transmit_module.video_signal_controller.n3199\
        );

    \I__982\ : InMux
    port map (
            O => \N__9755\,
            I => \N__9751\
        );

    \I__981\ : InMux
    port map (
            O => \N__9754\,
            I => \N__9748\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__9751\,
            I => \transmit_module.video_signal_controller.VGA_Y_7\
        );

    \I__979\ : LocalMux
    port map (
            O => \N__9748\,
            I => \transmit_module.video_signal_controller.VGA_Y_7\
        );

    \I__978\ : InMux
    port map (
            O => \N__9743\,
            I => \transmit_module.video_signal_controller.n3200\
        );

    \I__977\ : InMux
    port map (
            O => \N__9740\,
            I => \N__9736\
        );

    \I__976\ : InMux
    port map (
            O => \N__9739\,
            I => \N__9733\
        );

    \I__975\ : LocalMux
    port map (
            O => \N__9736\,
            I => \transmit_module.video_signal_controller.VGA_Y_8\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__9733\,
            I => \transmit_module.video_signal_controller.VGA_Y_8\
        );

    \I__973\ : InMux
    port map (
            O => \N__9728\,
            I => \bfn_12_15_0_\
        );

    \I__972\ : InMux
    port map (
            O => \N__9725\,
            I => \transmit_module.video_signal_controller.n3202\
        );

    \I__971\ : InMux
    port map (
            O => \N__9722\,
            I => \transmit_module.video_signal_controller.n3203\
        );

    \I__970\ : InMux
    port map (
            O => \N__9719\,
            I => \transmit_module.video_signal_controller.n3204\
        );

    \I__969\ : InMux
    port map (
            O => \N__9716\,
            I => \N__9711\
        );

    \I__968\ : InMux
    port map (
            O => \N__9715\,
            I => \N__9708\
        );

    \I__967\ : InMux
    port map (
            O => \N__9714\,
            I => \N__9705\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__9711\,
            I => \transmit_module.video_signal_controller.VGA_Y_11\
        );

    \I__965\ : LocalMux
    port map (
            O => \N__9708\,
            I => \transmit_module.video_signal_controller.VGA_Y_11\
        );

    \I__964\ : LocalMux
    port map (
            O => \N__9705\,
            I => \transmit_module.video_signal_controller.VGA_Y_11\
        );

    \I__963\ : InMux
    port map (
            O => \N__9698\,
            I => \N__9693\
        );

    \I__962\ : InMux
    port map (
            O => \N__9697\,
            I => \N__9690\
        );

    \I__961\ : InMux
    port map (
            O => \N__9696\,
            I => \N__9687\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__9693\,
            I => \transmit_module.video_signal_controller.VGA_Y_10\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__9690\,
            I => \transmit_module.video_signal_controller.VGA_Y_10\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__9687\,
            I => \transmit_module.video_signal_controller.VGA_Y_10\
        );

    \I__957\ : InMux
    port map (
            O => \N__9680\,
            I => \N__9677\
        );

    \I__956\ : LocalMux
    port map (
            O => \N__9677\,
            I => \transmit_module.Y_DELTA_PATTERN_94\
        );

    \I__955\ : InMux
    port map (
            O => \N__9674\,
            I => \N__9671\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__9671\,
            I => \transmit_module.Y_DELTA_PATTERN_93\
        );

    \I__953\ : InMux
    port map (
            O => \N__9668\,
            I => \N__9665\
        );

    \I__952\ : LocalMux
    port map (
            O => \N__9665\,
            I => \transmit_module.Y_DELTA_PATTERN_92\
        );

    \I__951\ : InMux
    port map (
            O => \N__9662\,
            I => \N__9659\
        );

    \I__950\ : LocalMux
    port map (
            O => \N__9659\,
            I => \transmit_module.Y_DELTA_PATTERN_87\
        );

    \I__949\ : InMux
    port map (
            O => \N__9656\,
            I => \N__9653\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__9653\,
            I => \transmit_module.Y_DELTA_PATTERN_89\
        );

    \I__947\ : InMux
    port map (
            O => \N__9650\,
            I => \N__9647\
        );

    \I__946\ : LocalMux
    port map (
            O => \N__9647\,
            I => \transmit_module.Y_DELTA_PATTERN_88\
        );

    \I__945\ : InMux
    port map (
            O => \N__9644\,
            I => \N__9641\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__9641\,
            I => \transmit_module.Y_DELTA_PATTERN_91\
        );

    \I__943\ : InMux
    port map (
            O => \N__9638\,
            I => \N__9635\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__9635\,
            I => \transmit_module.Y_DELTA_PATTERN_90\
        );

    \I__941\ : CEMux
    port map (
            O => \N__9632\,
            I => \N__9627\
        );

    \I__940\ : CEMux
    port map (
            O => \N__9631\,
            I => \N__9624\
        );

    \I__939\ : CEMux
    port map (
            O => \N__9630\,
            I => \N__9621\
        );

    \I__938\ : LocalMux
    port map (
            O => \N__9627\,
            I => \N__9618\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__9624\,
            I => \N__9613\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__9621\,
            I => \N__9613\
        );

    \I__935\ : Span12Mux_h
    port map (
            O => \N__9618\,
            I => \N__9610\
        );

    \I__934\ : Sp12to4
    port map (
            O => \N__9613\,
            I => \N__9607\
        );

    \I__933\ : Odrv12
    port map (
            O => \N__9610\,
            I => \transmit_module.n2209\
        );

    \I__932\ : Odrv12
    port map (
            O => \N__9607\,
            I => \transmit_module.n2209\
        );

    \I__931\ : InMux
    port map (
            O => \N__9602\,
            I => \bfn_12_14_0_\
        );

    \I__930\ : InMux
    port map (
            O => \N__9599\,
            I => \transmit_module.video_signal_controller.n3194\
        );

    \I__929\ : InMux
    port map (
            O => \N__9596\,
            I => \transmit_module.video_signal_controller.n3195\
        );

    \I__928\ : InMux
    port map (
            O => \N__9593\,
            I => \transmit_module.video_signal_controller.n3196\
        );

    \I__927\ : InMux
    port map (
            O => \N__9590\,
            I => \N__9587\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__9587\,
            I => \N__9584\
        );

    \I__925\ : Span4Mux_v
    port map (
            O => \N__9584\,
            I => \N__9581\
        );

    \I__924\ : Odrv4
    port map (
            O => \N__9581\,
            I => \tvp_video_buffer.BUFFER_0_2\
        );

    \I__923\ : InMux
    port map (
            O => \N__9578\,
            I => \N__9575\
        );

    \I__922\ : LocalMux
    port map (
            O => \N__9575\,
            I => \N__9572\
        );

    \I__921\ : Span12Mux_h
    port map (
            O => \N__9572\,
            I => \N__9569\
        );

    \I__920\ : Odrv12
    port map (
            O => \N__9569\,
            I => \TVP_VIDEO_c_3\
        );

    \I__919\ : InMux
    port map (
            O => \N__9566\,
            I => \N__9563\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__9563\,
            I => \tvp_video_buffer.BUFFER_0_3\
        );

    \I__917\ : InMux
    port map (
            O => \N__9560\,
            I => \N__9557\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__9557\,
            I => \transmit_module.X_DELTA_PATTERN_15\
        );

    \I__915\ : InMux
    port map (
            O => \N__9554\,
            I => \N__9551\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__9551\,
            I => \transmit_module.X_DELTA_PATTERN_14\
        );

    \I__913\ : InMux
    port map (
            O => \N__9548\,
            I => \transmit_module.video_signal_controller.n3186\
        );

    \I__912\ : InMux
    port map (
            O => \N__9545\,
            I => \transmit_module.video_signal_controller.n3187\
        );

    \I__911\ : InMux
    port map (
            O => \N__9542\,
            I => \transmit_module.video_signal_controller.n3188\
        );

    \I__910\ : InMux
    port map (
            O => \N__9539\,
            I => \transmit_module.video_signal_controller.n3189\
        );

    \I__909\ : InMux
    port map (
            O => \N__9536\,
            I => \bfn_11_18_0_\
        );

    \I__908\ : InMux
    port map (
            O => \N__9533\,
            I => \transmit_module.video_signal_controller.n3191\
        );

    \I__907\ : InMux
    port map (
            O => \N__9530\,
            I => \transmit_module.video_signal_controller.n3192\
        );

    \I__906\ : InMux
    port map (
            O => \N__9527\,
            I => \transmit_module.video_signal_controller.n3193\
        );

    \I__905\ : CEMux
    port map (
            O => \N__9524\,
            I => \N__9520\
        );

    \I__904\ : CEMux
    port map (
            O => \N__9523\,
            I => \N__9517\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__9520\,
            I => \N__9509\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__9517\,
            I => \N__9506\
        );

    \I__901\ : CEMux
    port map (
            O => \N__9516\,
            I => \N__9503\
        );

    \I__900\ : CEMux
    port map (
            O => \N__9515\,
            I => \N__9499\
        );

    \I__899\ : CEMux
    port map (
            O => \N__9514\,
            I => \N__9492\
        );

    \I__898\ : CEMux
    port map (
            O => \N__9513\,
            I => \N__9489\
        );

    \I__897\ : CEMux
    port map (
            O => \N__9512\,
            I => \N__9486\
        );

    \I__896\ : Span4Mux_v
    port map (
            O => \N__9509\,
            I => \N__9477\
        );

    \I__895\ : Span4Mux_h
    port map (
            O => \N__9506\,
            I => \N__9477\
        );

    \I__894\ : LocalMux
    port map (
            O => \N__9503\,
            I => \N__9477\
        );

    \I__893\ : CEMux
    port map (
            O => \N__9502\,
            I => \N__9474\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__9499\,
            I => \N__9471\
        );

    \I__891\ : CEMux
    port map (
            O => \N__9498\,
            I => \N__9468\
        );

    \I__890\ : CEMux
    port map (
            O => \N__9497\,
            I => \N__9465\
        );

    \I__889\ : CEMux
    port map (
            O => \N__9496\,
            I => \N__9462\
        );

    \I__888\ : CEMux
    port map (
            O => \N__9495\,
            I => \N__9459\
        );

    \I__887\ : LocalMux
    port map (
            O => \N__9492\,
            I => \N__9456\
        );

    \I__886\ : LocalMux
    port map (
            O => \N__9489\,
            I => \N__9451\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__9486\,
            I => \N__9451\
        );

    \I__884\ : CEMux
    port map (
            O => \N__9485\,
            I => \N__9448\
        );

    \I__883\ : CEMux
    port map (
            O => \N__9484\,
            I => \N__9445\
        );

    \I__882\ : Span4Mux_v
    port map (
            O => \N__9477\,
            I => \N__9442\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__9474\,
            I => \N__9435\
        );

    \I__880\ : Span4Mux_h
    port map (
            O => \N__9471\,
            I => \N__9435\
        );

    \I__879\ : LocalMux
    port map (
            O => \N__9468\,
            I => \N__9435\
        );

    \I__878\ : LocalMux
    port map (
            O => \N__9465\,
            I => \N__9428\
        );

    \I__877\ : LocalMux
    port map (
            O => \N__9462\,
            I => \N__9428\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__9459\,
            I => \N__9428\
        );

    \I__875\ : Span4Mux_h
    port map (
            O => \N__9456\,
            I => \N__9421\
        );

    \I__874\ : Span4Mux_h
    port map (
            O => \N__9451\,
            I => \N__9421\
        );

    \I__873\ : LocalMux
    port map (
            O => \N__9448\,
            I => \N__9421\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__9445\,
            I => \N__9418\
        );

    \I__871\ : Span4Mux_h
    port map (
            O => \N__9442\,
            I => \N__9415\
        );

    \I__870\ : Span4Mux_v
    port map (
            O => \N__9435\,
            I => \N__9412\
        );

    \I__869\ : Sp12to4
    port map (
            O => \N__9428\,
            I => \N__9409\
        );

    \I__868\ : Sp12to4
    port map (
            O => \N__9421\,
            I => \N__9406\
        );

    \I__867\ : Span4Mux_h
    port map (
            O => \N__9418\,
            I => \N__9403\
        );

    \I__866\ : Odrv4
    port map (
            O => \N__9415\,
            I => \transmit_module.n3683\
        );

    \I__865\ : Odrv4
    port map (
            O => \N__9412\,
            I => \transmit_module.n3683\
        );

    \I__864\ : Odrv12
    port map (
            O => \N__9409\,
            I => \transmit_module.n3683\
        );

    \I__863\ : Odrv12
    port map (
            O => \N__9406\,
            I => \transmit_module.n3683\
        );

    \I__862\ : Odrv4
    port map (
            O => \N__9403\,
            I => \transmit_module.n3683\
        );

    \I__861\ : CascadeMux
    port map (
            O => \N__9392\,
            I => \transmit_module.video_signal_controller.n6_cascade_\
        );

    \I__860\ : InMux
    port map (
            O => \N__9389\,
            I => \N__9386\
        );

    \I__859\ : LocalMux
    port map (
            O => \N__9386\,
            I => \transmit_module.ADDR_Y_COMPONENT_11\
        );

    \I__858\ : InMux
    port map (
            O => \N__9383\,
            I => \N__9380\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__9380\,
            I => \N__9377\
        );

    \I__856\ : Odrv4
    port map (
            O => \N__9377\,
            I => \transmit_module.ADDR_Y_COMPONENT_12\
        );

    \I__855\ : InMux
    port map (
            O => \N__9374\,
            I => \bfn_11_17_0_\
        );

    \I__854\ : InMux
    port map (
            O => \N__9371\,
            I => \transmit_module.video_signal_controller.n3183\
        );

    \I__853\ : InMux
    port map (
            O => \N__9368\,
            I => \transmit_module.video_signal_controller.n3184\
        );

    \I__852\ : InMux
    port map (
            O => \N__9365\,
            I => \transmit_module.video_signal_controller.n3185\
        );

    \I__851\ : InMux
    port map (
            O => \N__9362\,
            I => \N__9359\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__9359\,
            I => \N__9356\
        );

    \I__849\ : Span4Mux_h
    port map (
            O => \N__9356\,
            I => \N__9353\
        );

    \I__848\ : Odrv4
    port map (
            O => \N__9353\,
            I => \transmit_module.Y_DELTA_PATTERN_99\
        );

    \I__847\ : InMux
    port map (
            O => \N__9350\,
            I => \N__9347\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__9347\,
            I => \transmit_module.Y_DELTA_PATTERN_98\
        );

    \I__845\ : InMux
    port map (
            O => \N__9344\,
            I => \N__9341\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__9341\,
            I => \transmit_module.Y_DELTA_PATTERN_97\
        );

    \I__843\ : InMux
    port map (
            O => \N__9338\,
            I => \N__9335\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__9335\,
            I => \transmit_module.Y_DELTA_PATTERN_95\
        );

    \I__841\ : InMux
    port map (
            O => \N__9332\,
            I => \N__9329\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__9329\,
            I => \transmit_module.Y_DELTA_PATTERN_60\
        );

    \I__839\ : InMux
    port map (
            O => \N__9326\,
            I => \N__9323\
        );

    \I__838\ : LocalMux
    port map (
            O => \N__9323\,
            I => \transmit_module.Y_DELTA_PATTERN_59\
        );

    \I__837\ : InMux
    port map (
            O => \N__9320\,
            I => \N__9317\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__9317\,
            I => \transmit_module.Y_DELTA_PATTERN_58\
        );

    \I__835\ : InMux
    port map (
            O => \N__9314\,
            I => \N__9311\
        );

    \I__834\ : LocalMux
    port map (
            O => \N__9311\,
            I => \transmit_module.Y_DELTA_PATTERN_54\
        );

    \I__833\ : InMux
    port map (
            O => \N__9308\,
            I => \N__9305\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__9305\,
            I => \transmit_module.Y_DELTA_PATTERN_55\
        );

    \I__831\ : InMux
    port map (
            O => \N__9302\,
            I => \N__9299\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__9299\,
            I => \transmit_module.Y_DELTA_PATTERN_57\
        );

    \I__829\ : InMux
    port map (
            O => \N__9296\,
            I => \N__9293\
        );

    \I__828\ : LocalMux
    port map (
            O => \N__9293\,
            I => \transmit_module.Y_DELTA_PATTERN_56\
        );

    \I__827\ : InMux
    port map (
            O => \N__9290\,
            I => \N__9287\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__9287\,
            I => \transmit_module.Y_DELTA_PATTERN_86\
        );

    \I__825\ : InMux
    port map (
            O => \N__9284\,
            I => \N__9281\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__9281\,
            I => \transmit_module.Y_DELTA_PATTERN_96\
        );

    \I__823\ : InMux
    port map (
            O => \N__9278\,
            I => \N__9275\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__9275\,
            I => \transmit_module.Y_DELTA_PATTERN_47\
        );

    \I__821\ : InMux
    port map (
            O => \N__9272\,
            I => \N__9269\
        );

    \I__820\ : LocalMux
    port map (
            O => \N__9269\,
            I => \transmit_module.Y_DELTA_PATTERN_46\
        );

    \I__819\ : InMux
    port map (
            O => \N__9266\,
            I => \N__9263\
        );

    \I__818\ : LocalMux
    port map (
            O => \N__9263\,
            I => \transmit_module.Y_DELTA_PATTERN_49\
        );

    \I__817\ : InMux
    port map (
            O => \N__9260\,
            I => \N__9257\
        );

    \I__816\ : LocalMux
    port map (
            O => \N__9257\,
            I => \transmit_module.Y_DELTA_PATTERN_48\
        );

    \I__815\ : InMux
    port map (
            O => \N__9254\,
            I => \N__9251\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__9251\,
            I => \N__9248\
        );

    \I__813\ : Odrv12
    port map (
            O => \N__9248\,
            I => \transmit_module.Y_DELTA_PATTERN_53\
        );

    \I__812\ : InMux
    port map (
            O => \N__9245\,
            I => \N__9242\
        );

    \I__811\ : LocalMux
    port map (
            O => \N__9242\,
            I => \transmit_module.Y_DELTA_PATTERN_52\
        );

    \I__810\ : InMux
    port map (
            O => \N__9239\,
            I => \N__9236\
        );

    \I__809\ : LocalMux
    port map (
            O => \N__9236\,
            I => \transmit_module.Y_DELTA_PATTERN_51\
        );

    \I__808\ : InMux
    port map (
            O => \N__9233\,
            I => \N__9230\
        );

    \I__807\ : LocalMux
    port map (
            O => \N__9230\,
            I => \transmit_module.Y_DELTA_PATTERN_50\
        );

    \I__806\ : InMux
    port map (
            O => \N__9227\,
            I => \N__9224\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__9224\,
            I => \transmit_module.Y_DELTA_PATTERN_82\
        );

    \I__804\ : InMux
    port map (
            O => \N__9221\,
            I => \N__9218\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__9218\,
            I => \transmit_module.Y_DELTA_PATTERN_81\
        );

    \I__802\ : InMux
    port map (
            O => \N__9215\,
            I => \N__9212\
        );

    \I__801\ : LocalMux
    port map (
            O => \N__9212\,
            I => \transmit_module.Y_DELTA_PATTERN_83\
        );

    \I__800\ : InMux
    port map (
            O => \N__9209\,
            I => \N__9206\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__9206\,
            I => \transmit_module.Y_DELTA_PATTERN_85\
        );

    \I__798\ : InMux
    port map (
            O => \N__9203\,
            I => \N__9200\
        );

    \I__797\ : LocalMux
    port map (
            O => \N__9200\,
            I => \transmit_module.Y_DELTA_PATTERN_84\
        );

    \I__796\ : InMux
    port map (
            O => \N__9197\,
            I => \N__9194\
        );

    \I__795\ : LocalMux
    port map (
            O => \N__9194\,
            I => \transmit_module.Y_DELTA_PATTERN_26\
        );

    \I__794\ : InMux
    port map (
            O => \N__9191\,
            I => \N__9188\
        );

    \I__793\ : LocalMux
    port map (
            O => \N__9188\,
            I => \transmit_module.Y_DELTA_PATTERN_27\
        );

    \I__792\ : InMux
    port map (
            O => \N__9185\,
            I => \N__9182\
        );

    \I__791\ : LocalMux
    port map (
            O => \N__9182\,
            I => \transmit_module.Y_DELTA_PATTERN_28\
        );

    \I__790\ : InMux
    port map (
            O => \N__9179\,
            I => \N__9176\
        );

    \I__789\ : LocalMux
    port map (
            O => \N__9176\,
            I => \N__9173\
        );

    \I__788\ : Odrv12
    port map (
            O => \N__9173\,
            I => \transmit_module.Y_DELTA_PATTERN_30\
        );

    \I__787\ : InMux
    port map (
            O => \N__9170\,
            I => \N__9167\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__9167\,
            I => \transmit_module.Y_DELTA_PATTERN_29\
        );

    \I__785\ : InMux
    port map (
            O => \N__9164\,
            I => \N__9161\
        );

    \I__784\ : LocalMux
    port map (
            O => \N__9161\,
            I => \transmit_module.Y_DELTA_PATTERN_75\
        );

    \I__783\ : InMux
    port map (
            O => \N__9158\,
            I => \N__9155\
        );

    \I__782\ : LocalMux
    port map (
            O => \N__9155\,
            I => \transmit_module.Y_DELTA_PATTERN_78\
        );

    \I__781\ : InMux
    port map (
            O => \N__9152\,
            I => \N__9149\
        );

    \I__780\ : LocalMux
    port map (
            O => \N__9149\,
            I => \transmit_module.Y_DELTA_PATTERN_79\
        );

    \I__779\ : InMux
    port map (
            O => \N__9146\,
            I => \N__9143\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__9143\,
            I => \transmit_module.Y_DELTA_PATTERN_77\
        );

    \I__777\ : InMux
    port map (
            O => \N__9140\,
            I => \N__9137\
        );

    \I__776\ : LocalMux
    port map (
            O => \N__9137\,
            I => \transmit_module.Y_DELTA_PATTERN_76\
        );

    \I__775\ : InMux
    port map (
            O => \N__9134\,
            I => \N__9131\
        );

    \I__774\ : LocalMux
    port map (
            O => \N__9131\,
            I => \transmit_module.Y_DELTA_PATTERN_62\
        );

    \I__773\ : InMux
    port map (
            O => \N__9128\,
            I => \N__9125\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__9125\,
            I => \transmit_module.Y_DELTA_PATTERN_61\
        );

    \I__771\ : InMux
    port map (
            O => \N__9122\,
            I => \N__9119\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__9119\,
            I => \N__9116\
        );

    \I__769\ : Odrv12
    port map (
            O => \N__9116\,
            I => \transmit_module.Y_DELTA_PATTERN_80\
        );

    \I__768\ : InMux
    port map (
            O => \N__9113\,
            I => \N__9110\
        );

    \I__767\ : LocalMux
    port map (
            O => \N__9110\,
            I => \transmit_module.Y_DELTA_PATTERN_45\
        );

    \I__766\ : IoInMux
    port map (
            O => \N__9107\,
            I => \N__9104\
        );

    \I__765\ : LocalMux
    port map (
            O => \N__9104\,
            I => \N__9101\
        );

    \I__764\ : IoSpan4Mux
    port map (
            O => \N__9101\,
            I => \N__9098\
        );

    \I__763\ : Span4Mux_s3_h
    port map (
            O => \N__9098\,
            I => \N__9094\
        );

    \I__762\ : InMux
    port map (
            O => \N__9097\,
            I => \N__9091\
        );

    \I__761\ : Span4Mux_h
    port map (
            O => \N__9094\,
            I => \N__9086\
        );

    \I__760\ : LocalMux
    port map (
            O => \N__9091\,
            I => \N__9086\
        );

    \I__759\ : Span4Mux_h
    port map (
            O => \N__9086\,
            I => \N__9083\
        );

    \I__758\ : Sp12to4
    port map (
            O => \N__9083\,
            I => \N__9080\
        );

    \I__757\ : Span12Mux_v
    port map (
            O => \N__9080\,
            I => \N__9077\
        );

    \I__756\ : Odrv12
    port map (
            O => \N__9077\,
            I => \DEBUG_c_5_c\
        );

    \I__755\ : InMux
    port map (
            O => \N__9074\,
            I => \N__9071\
        );

    \I__754\ : LocalMux
    port map (
            O => \N__9071\,
            I => \N__9065\
        );

    \I__753\ : InMux
    port map (
            O => \N__9070\,
            I => \N__9062\
        );

    \I__752\ : InMux
    port map (
            O => \N__9069\,
            I => \N__9059\
        );

    \I__751\ : InMux
    port map (
            O => \N__9068\,
            I => \N__9054\
        );

    \I__750\ : Span4Mux_h
    port map (
            O => \N__9065\,
            I => \N__9051\
        );

    \I__749\ : LocalMux
    port map (
            O => \N__9062\,
            I => \N__9048\
        );

    \I__748\ : LocalMux
    port map (
            O => \N__9059\,
            I => \N__9045\
        );

    \I__747\ : InMux
    port map (
            O => \N__9058\,
            I => \N__9042\
        );

    \I__746\ : InMux
    port map (
            O => \N__9057\,
            I => \N__9039\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__9054\,
            I => \N__9035\
        );

    \I__744\ : Span4Mux_v
    port map (
            O => \N__9051\,
            I => \N__9032\
        );

    \I__743\ : Span4Mux_v
    port map (
            O => \N__9048\,
            I => \N__9027\
        );

    \I__742\ : Span4Mux_v
    port map (
            O => \N__9045\,
            I => \N__9027\
        );

    \I__741\ : LocalMux
    port map (
            O => \N__9042\,
            I => \N__9024\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__9039\,
            I => \N__9021\
        );

    \I__739\ : InMux
    port map (
            O => \N__9038\,
            I => \N__9018\
        );

    \I__738\ : Span12Mux_h
    port map (
            O => \N__9035\,
            I => \N__9015\
        );

    \I__737\ : Span4Mux_v
    port map (
            O => \N__9032\,
            I => \N__9010\
        );

    \I__736\ : Span4Mux_h
    port map (
            O => \N__9027\,
            I => \N__9010\
        );

    \I__735\ : Span12Mux_s3_v
    port map (
            O => \N__9024\,
            I => \N__9007\
        );

    \I__734\ : Span12Mux_s4_v
    port map (
            O => \N__9021\,
            I => \N__9002\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__9018\,
            I => \N__9002\
        );

    \I__732\ : Span12Mux_v
    port map (
            O => \N__9015\,
            I => \N__8992\
        );

    \I__731\ : Sp12to4
    port map (
            O => \N__9010\,
            I => \N__8992\
        );

    \I__730\ : Span12Mux_v
    port map (
            O => \N__9007\,
            I => \N__8992\
        );

    \I__729\ : Span12Mux_v
    port map (
            O => \N__9002\,
            I => \N__8992\
        );

    \I__728\ : InMux
    port map (
            O => \N__9001\,
            I => \N__8989\
        );

    \I__727\ : Odrv12
    port map (
            O => \N__8992\,
            I => \RX_DATA_3\
        );

    \I__726\ : LocalMux
    port map (
            O => \N__8989\,
            I => \RX_DATA_3\
        );

    \I__725\ : InMux
    port map (
            O => \N__8984\,
            I => \N__8981\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__8981\,
            I => \tvp_video_buffer.BUFFER_0_5\
        );

    \I__723\ : InMux
    port map (
            O => \N__8978\,
            I => \N__8975\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__8975\,
            I => \tvp_video_buffer.BUFFER_1_5\
        );

    \I__721\ : CascadeMux
    port map (
            O => \N__8972\,
            I => \N__8969\
        );

    \I__720\ : CascadeBuf
    port map (
            O => \N__8969\,
            I => \N__8965\
        );

    \I__719\ : CascadeMux
    port map (
            O => \N__8968\,
            I => \N__8962\
        );

    \I__718\ : CascadeMux
    port map (
            O => \N__8965\,
            I => \N__8959\
        );

    \I__717\ : CascadeBuf
    port map (
            O => \N__8962\,
            I => \N__8956\
        );

    \I__716\ : CascadeBuf
    port map (
            O => \N__8959\,
            I => \N__8953\
        );

    \I__715\ : CascadeMux
    port map (
            O => \N__8956\,
            I => \N__8950\
        );

    \I__714\ : CascadeMux
    port map (
            O => \N__8953\,
            I => \N__8947\
        );

    \I__713\ : CascadeBuf
    port map (
            O => \N__8950\,
            I => \N__8944\
        );

    \I__712\ : CascadeBuf
    port map (
            O => \N__8947\,
            I => \N__8941\
        );

    \I__711\ : CascadeMux
    port map (
            O => \N__8944\,
            I => \N__8938\
        );

    \I__710\ : CascadeMux
    port map (
            O => \N__8941\,
            I => \N__8935\
        );

    \I__709\ : CascadeBuf
    port map (
            O => \N__8938\,
            I => \N__8932\
        );

    \I__708\ : CascadeBuf
    port map (
            O => \N__8935\,
            I => \N__8929\
        );

    \I__707\ : CascadeMux
    port map (
            O => \N__8932\,
            I => \N__8926\
        );

    \I__706\ : CascadeMux
    port map (
            O => \N__8929\,
            I => \N__8923\
        );

    \I__705\ : CascadeBuf
    port map (
            O => \N__8926\,
            I => \N__8920\
        );

    \I__704\ : CascadeBuf
    port map (
            O => \N__8923\,
            I => \N__8917\
        );

    \I__703\ : CascadeMux
    port map (
            O => \N__8920\,
            I => \N__8914\
        );

    \I__702\ : CascadeMux
    port map (
            O => \N__8917\,
            I => \N__8911\
        );

    \I__701\ : CascadeBuf
    port map (
            O => \N__8914\,
            I => \N__8908\
        );

    \I__700\ : CascadeBuf
    port map (
            O => \N__8911\,
            I => \N__8905\
        );

    \I__699\ : CascadeMux
    port map (
            O => \N__8908\,
            I => \N__8902\
        );

    \I__698\ : CascadeMux
    port map (
            O => \N__8905\,
            I => \N__8899\
        );

    \I__697\ : CascadeBuf
    port map (
            O => \N__8902\,
            I => \N__8896\
        );

    \I__696\ : CascadeBuf
    port map (
            O => \N__8899\,
            I => \N__8893\
        );

    \I__695\ : CascadeMux
    port map (
            O => \N__8896\,
            I => \N__8890\
        );

    \I__694\ : CascadeMux
    port map (
            O => \N__8893\,
            I => \N__8887\
        );

    \I__693\ : CascadeBuf
    port map (
            O => \N__8890\,
            I => \N__8884\
        );

    \I__692\ : CascadeBuf
    port map (
            O => \N__8887\,
            I => \N__8881\
        );

    \I__691\ : CascadeMux
    port map (
            O => \N__8884\,
            I => \N__8878\
        );

    \I__690\ : CascadeMux
    port map (
            O => \N__8881\,
            I => \N__8875\
        );

    \I__689\ : CascadeBuf
    port map (
            O => \N__8878\,
            I => \N__8872\
        );

    \I__688\ : CascadeBuf
    port map (
            O => \N__8875\,
            I => \N__8869\
        );

    \I__687\ : CascadeMux
    port map (
            O => \N__8872\,
            I => \N__8866\
        );

    \I__686\ : CascadeMux
    port map (
            O => \N__8869\,
            I => \N__8863\
        );

    \I__685\ : CascadeBuf
    port map (
            O => \N__8866\,
            I => \N__8860\
        );

    \I__684\ : CascadeBuf
    port map (
            O => \N__8863\,
            I => \N__8857\
        );

    \I__683\ : CascadeMux
    port map (
            O => \N__8860\,
            I => \N__8854\
        );

    \I__682\ : CascadeMux
    port map (
            O => \N__8857\,
            I => \N__8851\
        );

    \I__681\ : CascadeBuf
    port map (
            O => \N__8854\,
            I => \N__8848\
        );

    \I__680\ : CascadeBuf
    port map (
            O => \N__8851\,
            I => \N__8845\
        );

    \I__679\ : CascadeMux
    port map (
            O => \N__8848\,
            I => \N__8842\
        );

    \I__678\ : CascadeMux
    port map (
            O => \N__8845\,
            I => \N__8839\
        );

    \I__677\ : CascadeBuf
    port map (
            O => \N__8842\,
            I => \N__8836\
        );

    \I__676\ : CascadeBuf
    port map (
            O => \N__8839\,
            I => \N__8833\
        );

    \I__675\ : CascadeMux
    port map (
            O => \N__8836\,
            I => \N__8830\
        );

    \I__674\ : CascadeMux
    port map (
            O => \N__8833\,
            I => \N__8827\
        );

    \I__673\ : CascadeBuf
    port map (
            O => \N__8830\,
            I => \N__8824\
        );

    \I__672\ : CascadeBuf
    port map (
            O => \N__8827\,
            I => \N__8821\
        );

    \I__671\ : CascadeMux
    port map (
            O => \N__8824\,
            I => \N__8818\
        );

    \I__670\ : CascadeMux
    port map (
            O => \N__8821\,
            I => \N__8815\
        );

    \I__669\ : CascadeBuf
    port map (
            O => \N__8818\,
            I => \N__8812\
        );

    \I__668\ : CascadeBuf
    port map (
            O => \N__8815\,
            I => \N__8809\
        );

    \I__667\ : CascadeMux
    port map (
            O => \N__8812\,
            I => \N__8806\
        );

    \I__666\ : CascadeMux
    port map (
            O => \N__8809\,
            I => \N__8803\
        );

    \I__665\ : CascadeBuf
    port map (
            O => \N__8806\,
            I => \N__8800\
        );

    \I__664\ : CascadeBuf
    port map (
            O => \N__8803\,
            I => \N__8797\
        );

    \I__663\ : CascadeMux
    port map (
            O => \N__8800\,
            I => \N__8794\
        );

    \I__662\ : CascadeMux
    port map (
            O => \N__8797\,
            I => \N__8791\
        );

    \I__661\ : CascadeBuf
    port map (
            O => \N__8794\,
            I => \N__8788\
        );

    \I__660\ : InMux
    port map (
            O => \N__8791\,
            I => \N__8785\
        );

    \I__659\ : CascadeMux
    port map (
            O => \N__8788\,
            I => \N__8782\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__8785\,
            I => \N__8779\
        );

    \I__657\ : InMux
    port map (
            O => \N__8782\,
            I => \N__8776\
        );

    \I__656\ : Span4Mux_h
    port map (
            O => \N__8779\,
            I => \N__8773\
        );

    \I__655\ : LocalMux
    port map (
            O => \N__8776\,
            I => \N__8770\
        );

    \I__654\ : Span4Mux_v
    port map (
            O => \N__8773\,
            I => \N__8767\
        );

    \I__653\ : Sp12to4
    port map (
            O => \N__8770\,
            I => \N__8764\
        );

    \I__652\ : Sp12to4
    port map (
            O => \N__8767\,
            I => \N__8761\
        );

    \I__651\ : Span12Mux_s5_v
    port map (
            O => \N__8764\,
            I => \N__8756\
        );

    \I__650\ : Span12Mux_h
    port map (
            O => \N__8761\,
            I => \N__8756\
        );

    \I__649\ : Odrv12
    port map (
            O => \N__8756\,
            I => n27
        );

    \I__648\ : InMux
    port map (
            O => \N__8753\,
            I => \N__8750\
        );

    \I__647\ : LocalMux
    port map (
            O => \N__8750\,
            I => \N__8747\
        );

    \I__646\ : Span4Mux_v
    port map (
            O => \N__8747\,
            I => \N__8744\
        );

    \I__645\ : Odrv4
    port map (
            O => \N__8744\,
            I => \line_buffer.n603\
        );

    \I__644\ : InMux
    port map (
            O => \N__8741\,
            I => \N__8738\
        );

    \I__643\ : LocalMux
    port map (
            O => \N__8738\,
            I => \N__8735\
        );

    \I__642\ : Span4Mux_v
    port map (
            O => \N__8735\,
            I => \N__8732\
        );

    \I__641\ : Odrv4
    port map (
            O => \N__8732\,
            I => \line_buffer.n595\
        );

    \I__640\ : InMux
    port map (
            O => \N__8729\,
            I => \N__8726\
        );

    \I__639\ : LocalMux
    port map (
            O => \N__8726\,
            I => \N__8723\
        );

    \I__638\ : Span4Mux_v
    port map (
            O => \N__8723\,
            I => \N__8720\
        );

    \I__637\ : Odrv4
    port map (
            O => \N__8720\,
            I => \line_buffer.n602\
        );

    \I__636\ : InMux
    port map (
            O => \N__8717\,
            I => \N__8714\
        );

    \I__635\ : LocalMux
    port map (
            O => \N__8714\,
            I => \N__8711\
        );

    \I__634\ : Span4Mux_v
    port map (
            O => \N__8711\,
            I => \N__8708\
        );

    \I__633\ : Odrv4
    port map (
            O => \N__8708\,
            I => \line_buffer.n594\
        );

    \I__632\ : InMux
    port map (
            O => \N__8705\,
            I => \N__8702\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__8702\,
            I => \N__8699\
        );

    \I__630\ : IoSpan4Mux
    port map (
            O => \N__8699\,
            I => \N__8696\
        );

    \I__629\ : Odrv4
    port map (
            O => \N__8696\,
            I => \TVP_VIDEO_c_2\
        );

    \I__628\ : InMux
    port map (
            O => \N__8693\,
            I => \N__8690\
        );

    \I__627\ : LocalMux
    port map (
            O => \N__8690\,
            I => \transmit_module.Y_DELTA_PATTERN_74\
        );

    \I__626\ : InMux
    port map (
            O => \N__8687\,
            I => \N__8684\
        );

    \I__625\ : LocalMux
    port map (
            O => \N__8684\,
            I => \transmit_module.Y_DELTA_PATTERN_67\
        );

    \I__624\ : InMux
    port map (
            O => \N__8681\,
            I => \N__8678\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__8678\,
            I => \transmit_module.Y_DELTA_PATTERN_65\
        );

    \I__622\ : InMux
    port map (
            O => \N__8675\,
            I => \N__8672\
        );

    \I__621\ : LocalMux
    port map (
            O => \N__8672\,
            I => \transmit_module.Y_DELTA_PATTERN_64\
        );

    \I__620\ : InMux
    port map (
            O => \N__8669\,
            I => \N__8666\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__8666\,
            I => \transmit_module.Y_DELTA_PATTERN_69\
        );

    \I__618\ : InMux
    port map (
            O => \N__8663\,
            I => \N__8660\
        );

    \I__617\ : LocalMux
    port map (
            O => \N__8660\,
            I => \transmit_module.Y_DELTA_PATTERN_68\
        );

    \I__616\ : InMux
    port map (
            O => \N__8657\,
            I => \N__8654\
        );

    \I__615\ : LocalMux
    port map (
            O => \N__8654\,
            I => \N__8651\
        );

    \I__614\ : Odrv4
    port map (
            O => \N__8651\,
            I => \transmit_module.Y_DELTA_PATTERN_24\
        );

    \I__613\ : InMux
    port map (
            O => \N__8648\,
            I => \N__8645\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__8645\,
            I => \transmit_module.Y_DELTA_PATTERN_25\
        );

    \I__611\ : InMux
    port map (
            O => \N__8642\,
            I => \N__8639\
        );

    \I__610\ : LocalMux
    port map (
            O => \N__8639\,
            I => \transmit_module.Y_DELTA_PATTERN_43\
        );

    \I__609\ : InMux
    port map (
            O => \N__8636\,
            I => \N__8633\
        );

    \I__608\ : LocalMux
    port map (
            O => \N__8633\,
            I => \N__8630\
        );

    \I__607\ : Odrv4
    port map (
            O => \N__8630\,
            I => \transmit_module.Y_DELTA_PATTERN_42\
        );

    \I__606\ : InMux
    port map (
            O => \N__8627\,
            I => \N__8624\
        );

    \I__605\ : LocalMux
    port map (
            O => \N__8624\,
            I => \transmit_module.Y_DELTA_PATTERN_44\
        );

    \I__604\ : InMux
    port map (
            O => \N__8621\,
            I => \N__8618\
        );

    \I__603\ : LocalMux
    port map (
            O => \N__8618\,
            I => \transmit_module.Y_DELTA_PATTERN_73\
        );

    \I__602\ : InMux
    port map (
            O => \N__8615\,
            I => \N__8612\
        );

    \I__601\ : LocalMux
    port map (
            O => \N__8612\,
            I => \transmit_module.Y_DELTA_PATTERN_72\
        );

    \I__600\ : InMux
    port map (
            O => \N__8609\,
            I => \N__8606\
        );

    \I__599\ : LocalMux
    port map (
            O => \N__8606\,
            I => \transmit_module.Y_DELTA_PATTERN_63\
        );

    \I__598\ : InMux
    port map (
            O => \N__8603\,
            I => \N__8600\
        );

    \I__597\ : LocalMux
    port map (
            O => \N__8600\,
            I => \N__8597\
        );

    \I__596\ : Odrv4
    port map (
            O => \N__8597\,
            I => \transmit_module.Y_DELTA_PATTERN_71\
        );

    \I__595\ : InMux
    port map (
            O => \N__8594\,
            I => \N__8591\
        );

    \I__594\ : LocalMux
    port map (
            O => \N__8591\,
            I => \transmit_module.Y_DELTA_PATTERN_70\
        );

    \I__593\ : InMux
    port map (
            O => \N__8588\,
            I => \N__8585\
        );

    \I__592\ : LocalMux
    port map (
            O => \N__8585\,
            I => \transmit_module.Y_DELTA_PATTERN_66\
        );

    \I__591\ : InMux
    port map (
            O => \N__8582\,
            I => \N__8579\
        );

    \I__590\ : LocalMux
    port map (
            O => \N__8579\,
            I => \transmit_module.Y_DELTA_PATTERN_14\
        );

    \I__589\ : InMux
    port map (
            O => \N__8576\,
            I => \N__8573\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__8573\,
            I => \transmit_module.Y_DELTA_PATTERN_39\
        );

    \I__587\ : InMux
    port map (
            O => \N__8570\,
            I => \N__8567\
        );

    \I__586\ : LocalMux
    port map (
            O => \N__8567\,
            I => \transmit_module.Y_DELTA_PATTERN_41\
        );

    \I__585\ : InMux
    port map (
            O => \N__8564\,
            I => \N__8561\
        );

    \I__584\ : LocalMux
    port map (
            O => \N__8561\,
            I => \transmit_module.Y_DELTA_PATTERN_40\
        );

    \I__583\ : InMux
    port map (
            O => \N__8558\,
            I => \N__8555\
        );

    \I__582\ : LocalMux
    port map (
            O => \N__8555\,
            I => \N__8552\
        );

    \I__581\ : Odrv4
    port map (
            O => \N__8552\,
            I => \transmit_module.Y_DELTA_PATTERN_13\
        );

    \I__580\ : InMux
    port map (
            O => \N__8549\,
            I => \N__8546\
        );

    \I__579\ : LocalMux
    port map (
            O => \N__8546\,
            I => \transmit_module.Y_DELTA_PATTERN_12\
        );

    \I__578\ : InMux
    port map (
            O => \N__8543\,
            I => \N__8540\
        );

    \I__577\ : LocalMux
    port map (
            O => \N__8540\,
            I => \transmit_module.Y_DELTA_PATTERN_7\
        );

    \I__576\ : InMux
    port map (
            O => \N__8537\,
            I => \N__8534\
        );

    \I__575\ : LocalMux
    port map (
            O => \N__8534\,
            I => \transmit_module.Y_DELTA_PATTERN_6\
        );

    \I__574\ : InMux
    port map (
            O => \N__8531\,
            I => \N__8528\
        );

    \I__573\ : LocalMux
    port map (
            O => \N__8528\,
            I => \transmit_module.Y_DELTA_PATTERN_11\
        );

    \I__572\ : InMux
    port map (
            O => \N__8525\,
            I => \N__8522\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__8522\,
            I => \transmit_module.Y_DELTA_PATTERN_10\
        );

    \I__570\ : InMux
    port map (
            O => \N__8519\,
            I => \N__8516\
        );

    \I__569\ : LocalMux
    port map (
            O => \N__8516\,
            I => \transmit_module.Y_DELTA_PATTERN_22\
        );

    \I__568\ : InMux
    port map (
            O => \N__8513\,
            I => \N__8510\
        );

    \I__567\ : LocalMux
    port map (
            O => \N__8510\,
            I => \transmit_module.Y_DELTA_PATTERN_21\
        );

    \I__566\ : InMux
    port map (
            O => \N__8507\,
            I => \N__8504\
        );

    \I__565\ : LocalMux
    port map (
            O => \N__8504\,
            I => \transmit_module.Y_DELTA_PATTERN_20\
        );

    \I__564\ : InMux
    port map (
            O => \N__8501\,
            I => \N__8498\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__8498\,
            I => \transmit_module.Y_DELTA_PATTERN_19\
        );

    \I__562\ : InMux
    port map (
            O => \N__8495\,
            I => \N__8492\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__8492\,
            I => \transmit_module.Y_DELTA_PATTERN_18\
        );

    \I__560\ : InMux
    port map (
            O => \N__8489\,
            I => \N__8486\
        );

    \I__559\ : LocalMux
    port map (
            O => \N__8486\,
            I => \transmit_module.Y_DELTA_PATTERN_15\
        );

    \I__558\ : InMux
    port map (
            O => \N__8483\,
            I => \N__8480\
        );

    \I__557\ : LocalMux
    port map (
            O => \N__8480\,
            I => \N__8477\
        );

    \I__556\ : Odrv4
    port map (
            O => \N__8477\,
            I => \transmit_module.Y_DELTA_PATTERN_23\
        );

    \I__555\ : InMux
    port map (
            O => \N__8474\,
            I => \N__8471\
        );

    \I__554\ : LocalMux
    port map (
            O => \N__8471\,
            I => \transmit_module.Y_DELTA_PATTERN_17\
        );

    \I__553\ : InMux
    port map (
            O => \N__8468\,
            I => \N__8465\
        );

    \I__552\ : LocalMux
    port map (
            O => \N__8465\,
            I => \transmit_module.Y_DELTA_PATTERN_16\
        );

    \I__551\ : InMux
    port map (
            O => \N__8462\,
            I => \N__8459\
        );

    \I__550\ : LocalMux
    port map (
            O => \N__8459\,
            I => \transmit_module.Y_DELTA_PATTERN_31\
        );

    \I__549\ : InMux
    port map (
            O => \N__8456\,
            I => \N__8453\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__8453\,
            I => \transmit_module.Y_DELTA_PATTERN_32\
        );

    \I__547\ : InMux
    port map (
            O => \N__8450\,
            I => \N__8447\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__8447\,
            I => \transmit_module.Y_DELTA_PATTERN_33\
        );

    \I__545\ : InMux
    port map (
            O => \N__8444\,
            I => \N__8441\
        );

    \I__544\ : LocalMux
    port map (
            O => \N__8441\,
            I => \transmit_module.Y_DELTA_PATTERN_38\
        );

    \I__543\ : InMux
    port map (
            O => \N__8438\,
            I => \N__8435\
        );

    \I__542\ : LocalMux
    port map (
            O => \N__8435\,
            I => \transmit_module.Y_DELTA_PATTERN_35\
        );

    \I__541\ : InMux
    port map (
            O => \N__8432\,
            I => \N__8429\
        );

    \I__540\ : LocalMux
    port map (
            O => \N__8429\,
            I => \transmit_module.Y_DELTA_PATTERN_34\
        );

    \I__539\ : InMux
    port map (
            O => \N__8426\,
            I => \N__8423\
        );

    \I__538\ : LocalMux
    port map (
            O => \N__8423\,
            I => \transmit_module.Y_DELTA_PATTERN_9\
        );

    \I__537\ : InMux
    port map (
            O => \N__8420\,
            I => \N__8417\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__8417\,
            I => \transmit_module.Y_DELTA_PATTERN_8\
        );

    \I__535\ : InMux
    port map (
            O => \N__8414\,
            I => \N__8411\
        );

    \I__534\ : LocalMux
    port map (
            O => \N__8411\,
            I => \transmit_module.Y_DELTA_PATTERN_37\
        );

    \I__533\ : InMux
    port map (
            O => \N__8408\,
            I => \N__8405\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__8405\,
            I => \transmit_module.Y_DELTA_PATTERN_36\
        );

    \IN_MUX_bfv_12_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_14_0_\
        );

    \IN_MUX_bfv_12_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \transmit_module.video_signal_controller.n3201\,
            carryinitout => \bfn_12_15_0_\
        );

    \IN_MUX_bfv_11_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_17_0_\
        );

    \IN_MUX_bfv_11_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \transmit_module.video_signal_controller.n3190\,
            carryinitout => \bfn_11_18_0_\
        );

    \IN_MUX_bfv_14_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_15_0_\
        );

    \IN_MUX_bfv_14_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \transmit_module.n3169\,
            carryinitout => \bfn_14_16_0_\
        );

    \IN_MUX_bfv_13_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_11_0_\
        );

    \IN_MUX_bfv_13_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \receive_module.rx_counter.n3182\,
            carryinitout => \bfn_13_12_0_\
        );

    \IN_MUX_bfv_13_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_9_0_\
        );

    \IN_MUX_bfv_13_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \receive_module.rx_counter.n3217\,
            carryinitout => \bfn_13_10_0_\
        );

    \IN_MUX_bfv_16_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_10_0_\
        );

    \IN_MUX_bfv_15_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_11_0_\
        );

    \IN_MUX_bfv_15_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \receive_module.n3156\,
            carryinitout => \bfn_15_12_0_\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \transmit_module.Y_DELTA_PATTERN_i35_LC_5_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8408\,
            lcout => \transmit_module.Y_DELTA_PATTERN_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23598\,
            ce => \N__9513\,
            sr => \N__20061\
        );

    \transmit_module.Y_DELTA_PATTERN_i37_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8444\,
            lcout => \transmit_module.Y_DELTA_PATTERN_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23598\,
            ce => \N__9513\,
            sr => \N__20061\
        );

    \transmit_module.Y_DELTA_PATTERN_i36_LC_5_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8414\,
            lcout => \transmit_module.Y_DELTA_PATTERN_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23598\,
            ce => \N__9513\,
            sr => \N__20061\
        );

    \transmit_module.Y_DELTA_PATTERN_i31_LC_6_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8456\,
            lcout => \transmit_module.Y_DELTA_PATTERN_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23729\,
            ce => \N__21426\,
            sr => \N__20012\
        );

    \transmit_module.Y_DELTA_PATTERN_i30_LC_6_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8462\,
            lcout => \transmit_module.Y_DELTA_PATTERN_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23729\,
            ce => \N__21426\,
            sr => \N__20012\
        );

    \transmit_module.Y_DELTA_PATTERN_i32_LC_6_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8450\,
            lcout => \transmit_module.Y_DELTA_PATTERN_32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23729\,
            ce => \N__21426\,
            sr => \N__20012\
        );

    \transmit_module.Y_DELTA_PATTERN_i33_LC_6_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8432\,
            lcout => \transmit_module.Y_DELTA_PATTERN_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23686\,
            ce => \N__9514\,
            sr => \N__20065\
        );

    \transmit_module.Y_DELTA_PATTERN_i38_LC_6_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8576\,
            lcout => \transmit_module.Y_DELTA_PATTERN_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23686\,
            ce => \N__9514\,
            sr => \N__20065\
        );

    \transmit_module.Y_DELTA_PATTERN_i34_LC_6_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8438\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.Y_DELTA_PATTERN_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23686\,
            ce => \N__9514\,
            sr => \N__20065\
        );

    \transmit_module.Y_DELTA_PATTERN_i9_LC_6_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8525\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.Y_DELTA_PATTERN_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23708\,
            ce => \N__21429\,
            sr => \N__20056\
        );

    \transmit_module.Y_DELTA_PATTERN_i7_LC_6_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8420\,
            lcout => \transmit_module.Y_DELTA_PATTERN_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23708\,
            ce => \N__21429\,
            sr => \N__20056\
        );

    \transmit_module.Y_DELTA_PATTERN_i8_LC_6_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8426\,
            lcout => \transmit_module.Y_DELTA_PATTERN_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23708\,
            ce => \N__21429\,
            sr => \N__20056\
        );

    \transmit_module.Y_DELTA_PATTERN_i22_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8483\,
            lcout => \transmit_module.Y_DELTA_PATTERN_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23599\,
            ce => \N__21382\,
            sr => \N__20036\
        );

    \transmit_module.Y_DELTA_PATTERN_i20_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8513\,
            lcout => \transmit_module.Y_DELTA_PATTERN_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23601\,
            ce => \N__21430\,
            sr => \N__20067\
        );

    \transmit_module.Y_DELTA_PATTERN_i21_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8519\,
            lcout => \transmit_module.Y_DELTA_PATTERN_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23601\,
            ce => \N__21430\,
            sr => \N__20067\
        );

    \transmit_module.Y_DELTA_PATTERN_i19_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8507\,
            lcout => \transmit_module.Y_DELTA_PATTERN_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23601\,
            ce => \N__21430\,
            sr => \N__20067\
        );

    \transmit_module.Y_DELTA_PATTERN_i18_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8501\,
            lcout => \transmit_module.Y_DELTA_PATTERN_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23601\,
            ce => \N__21430\,
            sr => \N__20067\
        );

    \transmit_module.Y_DELTA_PATTERN_i17_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8495\,
            lcout => \transmit_module.Y_DELTA_PATTERN_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23601\,
            ce => \N__21430\,
            sr => \N__20067\
        );

    \transmit_module.Y_DELTA_PATTERN_i15_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8468\,
            lcout => \transmit_module.Y_DELTA_PATTERN_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23703\,
            ce => \N__21407\,
            sr => \N__20007\
        );

    \transmit_module.Y_DELTA_PATTERN_i14_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8489\,
            lcout => \transmit_module.Y_DELTA_PATTERN_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23703\,
            ce => \N__21407\,
            sr => \N__20007\
        );

    \transmit_module.Y_DELTA_PATTERN_i23_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8657\,
            lcout => \transmit_module.Y_DELTA_PATTERN_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23703\,
            ce => \N__21407\,
            sr => \N__20007\
        );

    \transmit_module.Y_DELTA_PATTERN_i16_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8474\,
            lcout => \transmit_module.Y_DELTA_PATTERN_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23703\,
            ce => \N__21407\,
            sr => \N__20007\
        );

    \transmit_module.Y_DELTA_PATTERN_i13_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8582\,
            lcout => \transmit_module.Y_DELTA_PATTERN_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23703\,
            ce => \N__21407\,
            sr => \N__20007\
        );

    \transmit_module.Y_DELTA_PATTERN_i39_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8564\,
            lcout => \transmit_module.Y_DELTA_PATTERN_39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23634\,
            ce => \N__9512\,
            sr => \N__20060\
        );

    \transmit_module.Y_DELTA_PATTERN_i41_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8636\,
            lcout => \transmit_module.Y_DELTA_PATTERN_41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23634\,
            ce => \N__9512\,
            sr => \N__20060\
        );

    \transmit_module.Y_DELTA_PATTERN_i40_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8570\,
            lcout => \transmit_module.Y_DELTA_PATTERN_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23634\,
            ce => \N__9512\,
            sr => \N__20060\
        );

    \transmit_module.Y_DELTA_PATTERN_i12_LC_7_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8558\,
            lcout => \transmit_module.Y_DELTA_PATTERN_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23709\,
            ce => \N__21427\,
            sr => \N__20045\
        );

    \transmit_module.Y_DELTA_PATTERN_i11_LC_7_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8549\,
            lcout => \transmit_module.Y_DELTA_PATTERN_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23486\,
            ce => \N__21431\,
            sr => \N__20069\
        );

    \transmit_module.Y_DELTA_PATTERN_i5_LC_7_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8537\,
            lcout => \transmit_module.Y_DELTA_PATTERN_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23486\,
            ce => \N__21431\,
            sr => \N__20069\
        );

    \transmit_module.Y_DELTA_PATTERN_i6_LC_7_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8543\,
            lcout => \transmit_module.Y_DELTA_PATTERN_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23486\,
            ce => \N__21431\,
            sr => \N__20069\
        );

    \transmit_module.Y_DELTA_PATTERN_i10_LC_7_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8531\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.Y_DELTA_PATTERN_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23648\,
            ce => \N__21428\,
            sr => \N__20049\
        );

    \transmit_module.Y_DELTA_PATTERN_i71_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8615\,
            lcout => \transmit_module.Y_DELTA_PATTERN_71\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23715\,
            ce => \N__9524\,
            sr => \N__20057\
        );

    \transmit_module.Y_DELTA_PATTERN_i73_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8693\,
            lcout => \transmit_module.Y_DELTA_PATTERN_73\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23715\,
            ce => \N__9524\,
            sr => \N__20057\
        );

    \transmit_module.Y_DELTA_PATTERN_i72_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8621\,
            lcout => \transmit_module.Y_DELTA_PATTERN_72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23715\,
            ce => \N__9524\,
            sr => \N__20057\
        );

    \transmit_module.Y_DELTA_PATTERN_i78_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9152\,
            lcout => \transmit_module.Y_DELTA_PATTERN_78\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23715\,
            ce => \N__9524\,
            sr => \N__20057\
        );

    \transmit_module.Y_DELTA_PATTERN_i62_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8609\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.Y_DELTA_PATTERN_62\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23600\,
            ce => \N__9523\,
            sr => \N__20044\
        );

    \transmit_module.Y_DELTA_PATTERN_i63_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8675\,
            lcout => \transmit_module.Y_DELTA_PATTERN_63\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23687\,
            ce => \N__9516\,
            sr => \N__20011\
        );

    \transmit_module.Y_DELTA_PATTERN_i69_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8594\,
            lcout => \transmit_module.Y_DELTA_PATTERN_69\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23687\,
            ce => \N__9516\,
            sr => \N__20011\
        );

    \transmit_module.Y_DELTA_PATTERN_i70_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8603\,
            lcout => \transmit_module.Y_DELTA_PATTERN_70\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23687\,
            ce => \N__9516\,
            sr => \N__20011\
        );

    \transmit_module.Y_DELTA_PATTERN_i66_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8687\,
            lcout => \transmit_module.Y_DELTA_PATTERN_66\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23646\,
            ce => \N__9515\,
            sr => \N__19994\
        );

    \transmit_module.Y_DELTA_PATTERN_i65_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8588\,
            lcout => \transmit_module.Y_DELTA_PATTERN_65\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23646\,
            ce => \N__9515\,
            sr => \N__19994\
        );

    \transmit_module.Y_DELTA_PATTERN_i67_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8663\,
            lcout => \transmit_module.Y_DELTA_PATTERN_67\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23646\,
            ce => \N__9515\,
            sr => \N__19994\
        );

    \transmit_module.Y_DELTA_PATTERN_i64_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8681\,
            lcout => \transmit_module.Y_DELTA_PATTERN_64\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23646\,
            ce => \N__9515\,
            sr => \N__19994\
        );

    \transmit_module.Y_DELTA_PATTERN_i68_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8669\,
            lcout => \transmit_module.Y_DELTA_PATTERN_68\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23646\,
            ce => \N__9515\,
            sr => \N__19994\
        );

    \transmit_module.Y_DELTA_PATTERN_i99_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20684\,
            lcout => \transmit_module.Y_DELTA_PATTERN_99\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23714\,
            ce => \N__21381\,
            sr => \N__20006\
        );

    \transmit_module.Y_DELTA_PATTERN_i24_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8648\,
            lcout => \transmit_module.Y_DELTA_PATTERN_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23714\,
            ce => \N__21381\,
            sr => \N__20006\
        );

    \transmit_module.Y_DELTA_PATTERN_i25_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9197\,
            lcout => \transmit_module.Y_DELTA_PATTERN_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23714\,
            ce => \N__21381\,
            sr => \N__20006\
        );

    \transmit_module.Y_DELTA_PATTERN_i43_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8627\,
            lcout => \transmit_module.Y_DELTA_PATTERN_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23467\,
            ce => \N__9485\,
            sr => \N__20019\
        );

    \transmit_module.Y_DELTA_PATTERN_i42_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8642\,
            lcout => \transmit_module.Y_DELTA_PATTERN_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23467\,
            ce => \N__9485\,
            sr => \N__20019\
        );

    \transmit_module.Y_DELTA_PATTERN_i44_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9113\,
            lcout => \transmit_module.Y_DELTA_PATTERN_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23467\,
            ce => \N__9485\,
            sr => \N__20019\
        );

    \transmit_module.Y_DELTA_PATTERN_i45_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9272\,
            lcout => \transmit_module.Y_DELTA_PATTERN_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23467\,
            ce => \N__9485\,
            sr => \N__20019\
        );

    \tvp_video_buffer.BUFFER_0__i4_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__9097\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \tvp_video_buffer.BUFFER_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24148\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.WIRE_OUT_i3_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8978\,
            lcout => \RX_DATA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24148\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.BUFFER_0__i12_LC_9_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8984\,
            lcout => \tvp_video_buffer.BUFFER_1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24148\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1646_4_lut_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__20259\,
            in1 => \N__14165\,
            in2 => \N__20059\,
            in3 => \N__13604\,
            lcout => n27,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2194_3_lut_LC_9_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__24733\,
            in1 => \N__8753\,
            in2 => \_gnd_net_\,
            in3 => \N__8741\,
            lcout => \line_buffer.n3531\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2206_3_lut_LC_9_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__24779\,
            in1 => \N__8729\,
            in2 => \_gnd_net_\,
            in3 => \N__8717\,
            lcout => \line_buffer.n3543\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.BUFFER_0__i1_LC_10_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8705\,
            lcout => \tvp_video_buffer.BUFFER_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24098\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.Y_DELTA_PATTERN_i74_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9164\,
            lcout => \transmit_module.Y_DELTA_PATTERN_74\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23728\,
            ce => \N__9497\,
            sr => \N__20068\
        );

    \transmit_module.Y_DELTA_PATTERN_i75_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9140\,
            lcout => \transmit_module.Y_DELTA_PATTERN_75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23728\,
            ce => \N__9497\,
            sr => \N__20068\
        );

    \transmit_module.Y_DELTA_PATTERN_i77_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9158\,
            lcout => \transmit_module.Y_DELTA_PATTERN_77\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23728\,
            ce => \N__9497\,
            sr => \N__20068\
        );

    \transmit_module.Y_DELTA_PATTERN_i79_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9122\,
            lcout => \transmit_module.Y_DELTA_PATTERN_79\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23728\,
            ce => \N__9497\,
            sr => \N__20068\
        );

    \transmit_module.Y_DELTA_PATTERN_i76_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9146\,
            lcout => \transmit_module.Y_DELTA_PATTERN_76\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23728\,
            ce => \N__9497\,
            sr => \N__20068\
        );

    \transmit_module.Y_DELTA_PATTERN_i61_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__9134\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.Y_DELTA_PATTERN_61\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23677\,
            ce => \N__9502\,
            sr => \N__20002\
        );

    \transmit_module.Y_DELTA_PATTERN_i60_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9128\,
            lcout => \transmit_module.Y_DELTA_PATTERN_60\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23677\,
            ce => \N__9502\,
            sr => \N__20002\
        );

    \transmit_module.Y_DELTA_PATTERN_i53_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9314\,
            lcout => \transmit_module.Y_DELTA_PATTERN_53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23677\,
            ce => \N__9502\,
            sr => \N__20002\
        );

    \transmit_module.Y_DELTA_PATTERN_i80_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9221\,
            lcout => \transmit_module.Y_DELTA_PATTERN_80\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23677\,
            ce => \N__9502\,
            sr => \N__20002\
        );

    \transmit_module.Y_DELTA_PATTERN_i82_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9215\,
            lcout => \transmit_module.Y_DELTA_PATTERN_82\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23704\,
            ce => \N__9496\,
            sr => \N__20050\
        );

    \transmit_module.Y_DELTA_PATTERN_i81_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9227\,
            lcout => \transmit_module.Y_DELTA_PATTERN_81\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23704\,
            ce => \N__9496\,
            sr => \N__20050\
        );

    \transmit_module.Y_DELTA_PATTERN_i83_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9203\,
            lcout => \transmit_module.Y_DELTA_PATTERN_83\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23635\,
            ce => \N__9631\,
            sr => \N__20001\
        );

    \transmit_module.Y_DELTA_PATTERN_i85_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9290\,
            lcout => \transmit_module.Y_DELTA_PATTERN_85\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23635\,
            ce => \N__9631\,
            sr => \N__20001\
        );

    \transmit_module.Y_DELTA_PATTERN_i84_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9209\,
            lcout => \transmit_module.Y_DELTA_PATTERN_84\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23635\,
            ce => \N__9631\,
            sr => \N__20001\
        );

    \transmit_module.Y_DELTA_PATTERN_i26_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9191\,
            lcout => \transmit_module.Y_DELTA_PATTERN_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23710\,
            ce => \N__21331\,
            sr => \N__19876\
        );

    \transmit_module.Y_DELTA_PATTERN_i27_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9185\,
            lcout => \transmit_module.Y_DELTA_PATTERN_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23710\,
            ce => \N__21331\,
            sr => \N__19876\
        );

    \transmit_module.Y_DELTA_PATTERN_i28_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9170\,
            lcout => \transmit_module.Y_DELTA_PATTERN_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23710\,
            ce => \N__21331\,
            sr => \N__19876\
        );

    \transmit_module.Y_DELTA_PATTERN_i29_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9179\,
            lcout => \transmit_module.Y_DELTA_PATTERN_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23710\,
            ce => \N__21331\,
            sr => \N__19876\
        );

    \transmit_module.Y_DELTA_PATTERN_i49_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9233\,
            lcout => \transmit_module.Y_DELTA_PATTERN_49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23613\,
            ce => \N__9484\,
            sr => \N__19971\
        );

    \transmit_module.Y_DELTA_PATTERN_i47_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9260\,
            lcout => \transmit_module.Y_DELTA_PATTERN_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23613\,
            ce => \N__9484\,
            sr => \N__19971\
        );

    \transmit_module.Y_DELTA_PATTERN_i51_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9245\,
            lcout => \transmit_module.Y_DELTA_PATTERN_51\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23613\,
            ce => \N__9484\,
            sr => \N__19971\
        );

    \transmit_module.Y_DELTA_PATTERN_i46_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9278\,
            lcout => \transmit_module.Y_DELTA_PATTERN_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23613\,
            ce => \N__9484\,
            sr => \N__19971\
        );

    \transmit_module.Y_DELTA_PATTERN_i48_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9266\,
            lcout => \transmit_module.Y_DELTA_PATTERN_48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23613\,
            ce => \N__9484\,
            sr => \N__19971\
        );

    \transmit_module.Y_DELTA_PATTERN_i52_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9254\,
            lcout => \transmit_module.Y_DELTA_PATTERN_52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23613\,
            ce => \N__9484\,
            sr => \N__19971\
        );

    \transmit_module.Y_DELTA_PATTERN_i50_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9239\,
            lcout => \transmit_module.Y_DELTA_PATTERN_50\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23613\,
            ce => \N__9484\,
            sr => \N__19971\
        );

    \transmit_module.ADDR_Y_COMPONENT__i11_LC_10_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24641\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23649\,
            ce => \N__20764\,
            sr => \N__19997\
        );

    \transmit_module.ADDR_Y_COMPONENT__i5_LC_10_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13538\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23649\,
            ce => \N__20764\,
            sr => \N__19997\
        );

    \transmit_module.ADDR_Y_COMPONENT__i9_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14216\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23324\,
            ce => \N__20772\,
            sr => \N__20054\
        );

    \transmit_module.ADDR_Y_COMPONENT__i13_LC_10_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23918\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23553\,
            ce => \N__20774\,
            sr => \N__20055\
        );

    \transmit_module.Y_DELTA_PATTERN_i58_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9326\,
            lcout => \transmit_module.Y_DELTA_PATTERN_58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23637\,
            ce => \N__9498\,
            sr => \N__20043\
        );

    \transmit_module.Y_DELTA_PATTERN_i59_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9332\,
            lcout => \transmit_module.Y_DELTA_PATTERN_59\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23637\,
            ce => \N__9498\,
            sr => \N__20043\
        );

    \transmit_module.Y_DELTA_PATTERN_i57_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9320\,
            lcout => \transmit_module.Y_DELTA_PATTERN_57\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23474\,
            ce => \N__9495\,
            sr => \N__19964\
        );

    \transmit_module.Y_DELTA_PATTERN_i54_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9308\,
            lcout => \transmit_module.Y_DELTA_PATTERN_54\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23474\,
            ce => \N__9495\,
            sr => \N__19964\
        );

    \transmit_module.Y_DELTA_PATTERN_i55_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9296\,
            lcout => \transmit_module.Y_DELTA_PATTERN_55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23474\,
            ce => \N__9495\,
            sr => \N__19964\
        );

    \transmit_module.Y_DELTA_PATTERN_i56_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9302\,
            lcout => \transmit_module.Y_DELTA_PATTERN_56\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23474\,
            ce => \N__9495\,
            sr => \N__19964\
        );

    \transmit_module.Y_DELTA_PATTERN_i95_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9284\,
            lcout => \transmit_module.Y_DELTA_PATTERN_95\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23602\,
            ce => \N__9630\,
            sr => \N__20018\
        );

    \transmit_module.Y_DELTA_PATTERN_i86_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9662\,
            lcout => \transmit_module.Y_DELTA_PATTERN_86\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23602\,
            ce => \N__9630\,
            sr => \N__20018\
        );

    \transmit_module.Y_DELTA_PATTERN_i96_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9344\,
            lcout => \transmit_module.Y_DELTA_PATTERN_96\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23602\,
            ce => \N__9630\,
            sr => \N__20018\
        );

    \transmit_module.Y_DELTA_PATTERN_i98_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9362\,
            lcout => \transmit_module.Y_DELTA_PATTERN_98\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23602\,
            ce => \N__9630\,
            sr => \N__20018\
        );

    \transmit_module.Y_DELTA_PATTERN_i97_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9350\,
            lcout => \transmit_module.Y_DELTA_PATTERN_97\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23602\,
            ce => \N__9630\,
            sr => \N__20018\
        );

    \transmit_module.Y_DELTA_PATTERN_i94_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9338\,
            lcout => \transmit_module.Y_DELTA_PATTERN_94\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23602\,
            ce => \N__9630\,
            sr => \N__20018\
        );

    \transmit_module.ADDR_Y_COMPONENT__i6_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15179\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23550\,
            ce => \N__20738\,
            sr => \N__19963\
        );

    \transmit_module.ADDR_Y_COMPONENT__i7_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13490\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23550\,
            ce => \N__20738\,
            sr => \N__19963\
        );

    \transmit_module.ADDR_Y_COMPONENT__i12_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22269\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23550\,
            ce => \N__20738\,
            sr => \N__19963\
        );

    \transmit_module.video_signal_controller.i2183_3_lut_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__9861\,
            in1 => \N__9894\,
            in2 => \_gnd_net_\,
            in3 => \N__9838\,
            lcout => \transmit_module.video_signal_controller.n3520\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i127_2_lut_4_lut_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__11284\,
            in1 => \N__10870\,
            in2 => \N__20034\,
            in3 => \N__10818\,
            lcout => \transmit_module.n2209\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i483_2_lut_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10958\,
            in2 => \_gnd_net_\,
            in3 => \N__11009\,
            lcout => \transmit_module.video_signal_controller.n6_adj_622\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i127_2_lut_4_lut_rep_24_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__11285\,
            in1 => \N__10871\,
            in2 => \N__20035\,
            in3 => \N__10819\,
            lcout => \transmit_module.n3683\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_2_lut_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9754\,
            in2 => \_gnd_net_\,
            in3 => \N__9739\,
            lcout => \transmit_module.video_signal_controller.n3378\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_2_lut_3_lut_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__9714\,
            in1 => \N__9696\,
            in2 => \_gnd_net_\,
            in3 => \N__9960\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i4_4_lut_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__9984\,
            in1 => \N__9936\,
            in2 => \N__9392\,
            in3 => \N__9916\,
            lcout => \transmit_module.video_signal_controller.n2019\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__rep_1_i0_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__9389\,
            in1 => \N__20252\,
            in2 => \_gnd_net_\,
            in3 => \N__13655\,
            lcout => \TX_ADDR_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23335\,
            ce => \N__10246\,
            sr => \N__19981\
        );

    \transmit_module.BRAM_ADDR__i12_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__9383\,
            in1 => \N__20251\,
            in2 => \_gnd_net_\,
            in3 => \N__13643\,
            lcout => \TX_ADDR_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23335\,
            ce => \N__10246\,
            sr => \N__19981\
        );

    \transmit_module.video_signal_controller.VGA_X_i0_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10276\,
            in2 => \_gnd_net_\,
            in3 => \N__9374\,
            lcout => \transmit_module.video_signal_controller.VGA_X_0\,
            ltout => OPEN,
            carryin => \bfn_11_17_0_\,
            carryout => \transmit_module.video_signal_controller.n3183\,
            clk => \N__23482\,
            ce => 'H',
            sr => \N__9822\
        );

    \transmit_module.video_signal_controller.VGA_X_i1_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12458\,
            in2 => \_gnd_net_\,
            in3 => \N__9371\,
            lcout => \transmit_module.video_signal_controller.VGA_X_1\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3183\,
            carryout => \transmit_module.video_signal_controller.n3184\,
            clk => \N__23482\,
            ce => 'H',
            sr => \N__9822\
        );

    \transmit_module.video_signal_controller.VGA_X_i2_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12485\,
            in2 => \_gnd_net_\,
            in3 => \N__9368\,
            lcout => \transmit_module.video_signal_controller.VGA_X_2\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3184\,
            carryout => \transmit_module.video_signal_controller.n3185\,
            clk => \N__23482\,
            ce => 'H',
            sr => \N__9822\
        );

    \transmit_module.video_signal_controller.VGA_X_i3_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10399\,
            in2 => \_gnd_net_\,
            in3 => \N__9365\,
            lcout => \transmit_module.video_signal_controller.VGA_X_3\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3185\,
            carryout => \transmit_module.video_signal_controller.n3186\,
            clk => \N__23482\,
            ce => 'H',
            sr => \N__9822\
        );

    \transmit_module.video_signal_controller.VGA_X_i4_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10379\,
            in2 => \_gnd_net_\,
            in3 => \N__9548\,
            lcout => \transmit_module.video_signal_controller.VGA_X_4\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3186\,
            carryout => \transmit_module.video_signal_controller.n3187\,
            clk => \N__23482\,
            ce => 'H',
            sr => \N__9822\
        );

    \transmit_module.video_signal_controller.VGA_X_i5_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10327\,
            in2 => \_gnd_net_\,
            in3 => \N__9545\,
            lcout => \transmit_module.video_signal_controller.VGA_X_5\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3187\,
            carryout => \transmit_module.video_signal_controller.n3188\,
            clk => \N__23482\,
            ce => 'H',
            sr => \N__9822\
        );

    \transmit_module.video_signal_controller.VGA_X_i6_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10357\,
            in2 => \_gnd_net_\,
            in3 => \N__9542\,
            lcout => \transmit_module.video_signal_controller.VGA_X_6\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3188\,
            carryout => \transmit_module.video_signal_controller.n3189\,
            clk => \N__23482\,
            ce => 'H',
            sr => \N__9822\
        );

    \transmit_module.video_signal_controller.VGA_X_i7_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10294\,
            in2 => \_gnd_net_\,
            in3 => \N__9539\,
            lcout => \transmit_module.video_signal_controller.VGA_X_7\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3189\,
            carryout => \transmit_module.video_signal_controller.n3190\,
            clk => \N__23482\,
            ce => 'H',
            sr => \N__9822\
        );

    \transmit_module.video_signal_controller.VGA_X_i8_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11846\,
            in2 => \_gnd_net_\,
            in3 => \N__9536\,
            lcout => \transmit_module.video_signal_controller.VGA_X_8\,
            ltout => OPEN,
            carryin => \bfn_11_18_0_\,
            carryout => \transmit_module.video_signal_controller.n3191\,
            clk => \N__23647\,
            ce => 'H',
            sr => \N__9823\
        );

    \transmit_module.video_signal_controller.VGA_X_i9_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12407\,
            in2 => \_gnd_net_\,
            in3 => \N__9533\,
            lcout => \transmit_module.video_signal_controller.VGA_X_9\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3191\,
            carryout => \transmit_module.video_signal_controller.n3192\,
            clk => \N__23647\,
            ce => 'H',
            sr => \N__9823\
        );

    \transmit_module.video_signal_controller.VGA_X_i10_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11548\,
            in2 => \_gnd_net_\,
            in3 => \N__9530\,
            lcout => \transmit_module.video_signal_controller.VGA_X_10\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3192\,
            carryout => \transmit_module.video_signal_controller.n3193\,
            clk => \N__23647\,
            ce => 'H',
            sr => \N__9823\
        );

    \transmit_module.video_signal_controller.VGA_X_i11_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14277\,
            in2 => \_gnd_net_\,
            in3 => \N__9527\,
            lcout => \transmit_module.video_signal_controller.VGA_X_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23647\,
            ce => 'H',
            sr => \N__9823\
        );

    \transmit_module.i1699_4_lut_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011111110100"
        )
    port map (
            in0 => \N__20682\,
            in1 => \N__20264\,
            in2 => \N__20033\,
            in3 => \N__15146\,
            lcout => \transmit_module.n2073\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.BUFFER_0__i9_LC_12_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9590\,
            lcout => \tvp_video_buffer.BUFFER_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24099\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.BUFFER_0__i10_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9566\,
            lcout => \tvp_video_buffer.BUFFER_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24114\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.BUFFER_0__i2_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9578\,
            lcout => \tvp_video_buffer.BUFFER_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24114\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.WIRE_OUT_i6_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10412\,
            lcout => \RX_DATA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24121\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.X_DELTA_PATTERN_i15_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14675\,
            lcout => \transmit_module.X_DELTA_PATTERN_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23604\,
            ce => \N__21475\,
            sr => \N__21355\
        );

    \transmit_module.X_DELTA_PATTERN_i13_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9554\,
            lcout => \transmit_module.X_DELTA_PATTERN_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23604\,
            ce => \N__21475\,
            sr => \N__21355\
        );

    \transmit_module.X_DELTA_PATTERN_i14_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9560\,
            lcout => \transmit_module.X_DELTA_PATTERN_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23604\,
            ce => \N__21475\,
            sr => \N__21355\
        );

    \transmit_module.Y_DELTA_PATTERN_i89_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9638\,
            lcout => \transmit_module.Y_DELTA_PATTERN_89\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23532\,
            ce => \N__9632\,
            sr => \N__20017\
        );

    \transmit_module.Y_DELTA_PATTERN_i92_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9674\,
            lcout => \transmit_module.Y_DELTA_PATTERN_92\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23532\,
            ce => \N__9632\,
            sr => \N__20017\
        );

    \transmit_module.Y_DELTA_PATTERN_i93_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9680\,
            lcout => \transmit_module.Y_DELTA_PATTERN_93\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23532\,
            ce => \N__9632\,
            sr => \N__20017\
        );

    \transmit_module.Y_DELTA_PATTERN_i91_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9668\,
            lcout => \transmit_module.Y_DELTA_PATTERN_91\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23532\,
            ce => \N__9632\,
            sr => \N__20017\
        );

    \transmit_module.Y_DELTA_PATTERN_i87_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9650\,
            lcout => \transmit_module.Y_DELTA_PATTERN_87\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23532\,
            ce => \N__9632\,
            sr => \N__20017\
        );

    \transmit_module.Y_DELTA_PATTERN_i88_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9656\,
            lcout => \transmit_module.Y_DELTA_PATTERN_88\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23532\,
            ce => \N__9632\,
            sr => \N__20017\
        );

    \transmit_module.Y_DELTA_PATTERN_i90_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9644\,
            lcout => \transmit_module.Y_DELTA_PATTERN_90\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23532\,
            ce => \N__9632\,
            sr => \N__20017\
        );

    \transmit_module.video_signal_controller.VGA_Y_i0_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10975\,
            in2 => \_gnd_net_\,
            in3 => \N__9602\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_0\,
            ltout => OPEN,
            carryin => \bfn_12_14_0_\,
            carryout => \transmit_module.video_signal_controller.n3194\,
            clk => \N__23667\,
            ce => \N__9824\,
            sr => \N__9782\
        );

    \transmit_module.video_signal_controller.VGA_Y_i1_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11013\,
            in2 => \_gnd_net_\,
            in3 => \N__9599\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_1\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3194\,
            carryout => \transmit_module.video_signal_controller.n3195\,
            clk => \N__23667\,
            ce => \N__9824\,
            sr => \N__9782\
        );

    \transmit_module.video_signal_controller.VGA_Y_i2_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10962\,
            in2 => \_gnd_net_\,
            in3 => \N__9596\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_2\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3195\,
            carryout => \transmit_module.video_signal_controller.n3196\,
            clk => \N__23667\,
            ce => \N__9824\,
            sr => \N__9782\
        );

    \transmit_module.video_signal_controller.VGA_Y_i3_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9893\,
            in2 => \_gnd_net_\,
            in3 => \N__9593\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_3\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3196\,
            carryout => \transmit_module.video_signal_controller.n3197\,
            clk => \N__23667\,
            ce => \N__9824\,
            sr => \N__9782\
        );

    \transmit_module.video_signal_controller.VGA_Y_i4_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9860\,
            in2 => \_gnd_net_\,
            in3 => \N__9764\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_4\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3197\,
            carryout => \transmit_module.video_signal_controller.n3198\,
            clk => \N__23667\,
            ce => \N__9824\,
            sr => \N__9782\
        );

    \transmit_module.video_signal_controller.VGA_Y_i5_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9988\,
            in2 => \_gnd_net_\,
            in3 => \N__9761\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_5\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3198\,
            carryout => \transmit_module.video_signal_controller.n3199\,
            clk => \N__23667\,
            ce => \N__9824\,
            sr => \N__9782\
        );

    \transmit_module.video_signal_controller.VGA_Y_i6_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9964\,
            in2 => \_gnd_net_\,
            in3 => \N__9758\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_6\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3199\,
            carryout => \transmit_module.video_signal_controller.n3200\,
            clk => \N__23667\,
            ce => \N__9824\,
            sr => \N__9782\
        );

    \transmit_module.video_signal_controller.VGA_Y_i7_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9755\,
            in2 => \_gnd_net_\,
            in3 => \N__9743\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_7\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3200\,
            carryout => \transmit_module.video_signal_controller.n3201\,
            clk => \N__23667\,
            ce => \N__9824\,
            sr => \N__9782\
        );

    \transmit_module.video_signal_controller.VGA_Y_i8_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9740\,
            in2 => \_gnd_net_\,
            in3 => \N__9728\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_8\,
            ltout => OPEN,
            carryin => \bfn_12_15_0_\,
            carryout => \transmit_module.video_signal_controller.n3202\,
            clk => \N__23656\,
            ce => \N__9818\,
            sr => \N__9778\
        );

    \transmit_module.video_signal_controller.VGA_Y_i9_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9938\,
            in2 => \_gnd_net_\,
            in3 => \N__9725\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_9\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3202\,
            carryout => \transmit_module.video_signal_controller.n3203\,
            clk => \N__23656\,
            ce => \N__9818\,
            sr => \N__9778\
        );

    \transmit_module.video_signal_controller.VGA_Y_i10_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9698\,
            in2 => \_gnd_net_\,
            in3 => \N__9722\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_10\,
            ltout => OPEN,
            carryin => \transmit_module.video_signal_controller.n3203\,
            carryout => \transmit_module.video_signal_controller.n3204\,
            clk => \N__23656\,
            ce => \N__9818\,
            sr => \N__9778\
        );

    \transmit_module.video_signal_controller.VGA_Y_i11_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9716\,
            in2 => \_gnd_net_\,
            in3 => \N__9719\,
            lcout => \transmit_module.video_signal_controller.VGA_Y_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23656\,
            ce => \N__9818\,
            sr => \N__9778\
        );

    \transmit_module.video_signal_controller.i1_2_lut_rep_17_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9715\,
            in2 => \_gnd_net_\,
            in3 => \N__9697\,
            lcout => \transmit_module.video_signal_controller.n3676\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i2_3_lut_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__9895\,
            in1 => \N__10964\,
            in2 => \_gnd_net_\,
            in3 => \N__11015\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n3485_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i2_4_lut_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__9989\,
            in1 => \N__9865\,
            in2 => \N__9968\,
            in3 => \N__9965\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n3464_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_4_lut_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101010"
        )
    port map (
            in0 => \N__9944\,
            in1 => \N__9937\,
            in2 => \N__9920\,
            in3 => \N__9917\,
            lcout => \transmit_module.video_signal_controller.n3382\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i6_3_lut_LC_12_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__20678\,
            in1 => \N__9905\,
            in2 => \_gnd_net_\,
            in3 => \N__13533\,
            lcout => \transmit_module.n111\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i2_3_lut_adj_34_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__10361\,
            in1 => \N__10331\,
            in2 => \_gnd_net_\,
            in3 => \N__10293\,
            lcout => \transmit_module.video_signal_controller.n2017\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_4_lut_adj_28_LC_12_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111100000"
        )
    port map (
            in0 => \N__9896\,
            in1 => \N__9872\,
            in2 => \N__9866\,
            in3 => \N__9839\,
            lcout => \transmit_module.video_signal_controller.VGA_VISIBLE_N_588\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_2_lut_adj_33_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10376\,
            in2 => \_gnd_net_\,
            in3 => \N__10394\,
            lcout => \transmit_module.video_signal_controller.n3366\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1738_4_lut_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101100"
        )
    port map (
            in0 => \N__11543\,
            in1 => \N__14269\,
            in2 => \N__10925\,
            in3 => \N__12406\,
            lcout => \transmit_module.video_signal_controller.n2050\,
            ltout => \transmit_module.video_signal_controller.n2050_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1163_2_lut_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9785\,
            in3 => \N__13577\,
            lcout => \transmit_module.video_signal_controller.n2398\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1_4_lut_adj_31_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011001100"
        )
    port map (
            in0 => \N__10377\,
            in1 => \N__10355\,
            in2 => \N__10400\,
            in3 => \N__10325\,
            lcout => \transmit_module.video_signal_controller.n55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i2_4_lut_adj_30_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010000000"
        )
    port map (
            in0 => \N__12456\,
            in1 => \N__10395\,
            in2 => \N__12483\,
            in3 => \N__10275\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n3482_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i3_4_lut_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__10378\,
            in1 => \N__10356\,
            in2 => \N__10334\,
            in3 => \N__10326\,
            lcout => OPEN,
            ltout => \transmit_module.video_signal_controller.n3478_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i2_4_lut_adj_32_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010101000100"
        )
    port map (
            in0 => \N__11544\,
            in1 => \N__10304\,
            in2 => \N__10298\,
            in3 => \N__10295\,
            lcout => \transmit_module.video_signal_controller.n7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1715_2_lut_3_lut_LC_12_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12455\,
            in2 => \N__10277\,
            in3 => \N__12473\,
            lcout => \transmit_module.video_signal_controller.n2958\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i13_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__10259\,
            in1 => \N__20253\,
            in2 => \_gnd_net_\,
            in3 => \N__13628\,
            lcout => \TX_ADDR_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23571\,
            ce => \N__10247\,
            sr => \N__19935\
        );

    \transmit_module.i1653_4_lut_LC_12_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__20226\,
            in1 => \N__12427\,
            in2 => \N__19995\,
            in3 => \N__12370\,
            lcout => n20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.ADDR_Y_COMPONENT__i3_LC_12_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16409\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23418\,
            ce => \N__20773\,
            sr => \N__20032\
        );

    \tvp_video_buffer.WIRE_OUT_i0_LC_13_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10001\,
            lcout => \RX_DATA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24102\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.BUFFER_0__i3_LC_13_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__10649\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \tvp_video_buffer.BUFFER_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24105\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.BUFFER_0__i11_LC_13_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10634\,
            lcout => \tvp_video_buffer.BUFFER_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24105\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.BUFFER_0__i7_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10628\,
            lcout => \tvp_video_buffer.BUFFER_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24110\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.WIRE_OUT_i1_LC_13_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10616\,
            lcout => \RX_DATA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24110\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.WIRE_OUT_i2_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10523\,
            lcout => \RX_DATA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24110\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.BUFFER_0__i15_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10418\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \tvp_video_buffer.BUFFER_1_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24115\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.X_246__i0_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12566\,
            in2 => \_gnd_net_\,
            in3 => \N__10406\,
            lcout => \receive_module.rx_counter.X_0\,
            ltout => OPEN,
            carryin => \bfn_13_9_0_\,
            carryout => \receive_module.rx_counter.n3210\,
            clk => \N__24118\,
            ce => 'H',
            sr => \N__12502\
        );

    \receive_module.rx_counter.X_246__i1_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12578\,
            in2 => \_gnd_net_\,
            in3 => \N__10403\,
            lcout => \receive_module.rx_counter.X_1\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3210\,
            carryout => \receive_module.rx_counter.n3211\,
            clk => \N__24118\,
            ce => 'H',
            sr => \N__12502\
        );

    \receive_module.rx_counter.X_246__i2_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12554\,
            in2 => \_gnd_net_\,
            in3 => \N__10763\,
            lcout => \receive_module.rx_counter.X_2\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3211\,
            carryout => \receive_module.rx_counter.n3212\,
            clk => \N__24118\,
            ce => 'H',
            sr => \N__12502\
        );

    \receive_module.rx_counter.X_246__i3_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12989\,
            in2 => \_gnd_net_\,
            in3 => \N__10760\,
            lcout => \receive_module.rx_counter.X_3\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3212\,
            carryout => \receive_module.rx_counter.n3213\,
            clk => \N__24118\,
            ce => 'H',
            sr => \N__12502\
        );

    \receive_module.rx_counter.X_246__i4_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12536\,
            in2 => \_gnd_net_\,
            in3 => \N__10757\,
            lcout => \receive_module.rx_counter.X_4\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3213\,
            carryout => \receive_module.rx_counter.n3214\,
            clk => \N__24118\,
            ce => 'H',
            sr => \N__12502\
        );

    \receive_module.rx_counter.X_246__i5_LC_13_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12971\,
            in2 => \_gnd_net_\,
            in3 => \N__10754\,
            lcout => \receive_module.rx_counter.X_5\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3214\,
            carryout => \receive_module.rx_counter.n3215\,
            clk => \N__24118\,
            ce => 'H',
            sr => \N__12502\
        );

    \receive_module.rx_counter.X_246__i6_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12521\,
            in2 => \_gnd_net_\,
            in3 => \N__10751\,
            lcout => \receive_module.rx_counter.X_6\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3215\,
            carryout => \receive_module.rx_counter.n3216\,
            clk => \N__24118\,
            ce => 'H',
            sr => \N__12502\
        );

    \receive_module.rx_counter.X_246__i7_LC_13_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12953\,
            in2 => \_gnd_net_\,
            in3 => \N__10748\,
            lcout => \receive_module.rx_counter.X_7\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3216\,
            carryout => \receive_module.rx_counter.n3217\,
            clk => \N__24118\,
            ce => 'H',
            sr => \N__12502\
        );

    \receive_module.rx_counter.X_246__i8_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12854\,
            in2 => \_gnd_net_\,
            in3 => \N__10745\,
            lcout => \receive_module.rx_counter.X_8\,
            ltout => OPEN,
            carryin => \bfn_13_10_0_\,
            carryout => \receive_module.rx_counter.n3218\,
            clk => \N__24122\,
            ce => 'H',
            sr => \N__12506\
        );

    \receive_module.rx_counter.X_246__i9_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12835\,
            in2 => \_gnd_net_\,
            in3 => \N__10742\,
            lcout => \receive_module.rx_counter.X_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24122\,
            ce => 'H',
            sr => \N__12506\
        );

    \receive_module.rx_counter.Y__i0_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13194\,
            in2 => \_gnd_net_\,
            in3 => \N__10739\,
            lcout => \receive_module.rx_counter.Y_0\,
            ltout => OPEN,
            carryin => \bfn_13_11_0_\,
            carryout => \receive_module.rx_counter.n3175\,
            clk => \N__24127\,
            ce => \N__12913\,
            sr => \N__17554\
        );

    \receive_module.rx_counter.Y__i1_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13219\,
            in2 => \_gnd_net_\,
            in3 => \N__10787\,
            lcout => \receive_module.rx_counter.Y_1\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3175\,
            carryout => \receive_module.rx_counter.n3176\,
            clk => \N__24127\,
            ce => \N__12913\,
            sr => \N__17554\
        );

    \receive_module.rx_counter.Y__i2_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13165\,
            in2 => \_gnd_net_\,
            in3 => \N__10784\,
            lcout => \receive_module.rx_counter.Y_2\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3176\,
            carryout => \receive_module.rx_counter.n3177\,
            clk => \N__24127\,
            ce => \N__12913\,
            sr => \N__17554\
        );

    \receive_module.rx_counter.Y__i3_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13135\,
            in2 => \_gnd_net_\,
            in3 => \N__10781\,
            lcout => \receive_module.rx_counter.Y_3\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3177\,
            carryout => \receive_module.rx_counter.n3178\,
            clk => \N__24127\,
            ce => \N__12913\,
            sr => \N__17554\
        );

    \receive_module.rx_counter.Y__i4_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13110\,
            in2 => \_gnd_net_\,
            in3 => \N__10778\,
            lcout => \receive_module.rx_counter.Y_4\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3178\,
            carryout => \receive_module.rx_counter.n3179\,
            clk => \N__24127\,
            ce => \N__12913\,
            sr => \N__17554\
        );

    \receive_module.rx_counter.Y__i5_LC_13_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12794\,
            in2 => \_gnd_net_\,
            in3 => \N__10775\,
            lcout => \receive_module.rx_counter.Y_5\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3179\,
            carryout => \receive_module.rx_counter.n3180\,
            clk => \N__24127\,
            ce => \N__12913\,
            sr => \N__17554\
        );

    \receive_module.rx_counter.Y__i6_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12812\,
            in2 => \_gnd_net_\,
            in3 => \N__10772\,
            lcout => \receive_module.rx_counter.Y_6\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3180\,
            carryout => \receive_module.rx_counter.n3181\,
            clk => \N__24127\,
            ce => \N__12913\,
            sr => \N__17554\
        );

    \receive_module.rx_counter.Y__i7_LC_13_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13309\,
            in2 => \_gnd_net_\,
            in3 => \N__10769\,
            lcout => \receive_module.rx_counter.Y_7\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3181\,
            carryout => \receive_module.rx_counter.n3182\,
            clk => \N__24127\,
            ce => \N__12913\,
            sr => \N__17554\
        );

    \receive_module.rx_counter.Y__i8_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13264\,
            in2 => \_gnd_net_\,
            in3 => \N__10766\,
            lcout => \receive_module.rx_counter.Y_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24131\,
            ce => \N__12914\,
            sr => \N__17541\
        );

    \receive_module.rx_counter.i2_2_lut_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13115\,
            in2 => \_gnd_net_\,
            in3 => \N__13310\,
            lcout => \receive_module.rx_counter.n10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i6_4_lut_LC_13_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__13223\,
            in1 => \N__13139\,
            in2 => \N__13268\,
            in3 => \N__13169\,
            lcout => OPEN,
            ltout => \receive_module.rx_counter.n14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.SYNC_46_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__10910\,
            in1 => \N__13199\,
            in2 => \N__10904\,
            in3 => \N__13283\,
            lcout => \RX_TX_SYNC\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24135\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i127_2_lut_4_lut_rep_23_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110011001100"
        )
    port map (
            in0 => \N__10808\,
            in1 => \N__19692\,
            in2 => \N__11283\,
            in3 => \N__10861\,
            lcout => \transmit_module.n3682\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2193_3_lut_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__24714\,
            in1 => \N__10901\,
            in2 => \_gnd_net_\,
            in3 => \N__10886\,
            lcout => \line_buffer.n3530\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.old_VGA_HS_40_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__10809\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.old_VGA_HS\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23603\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i2_3_lut_rep_19_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__10860\,
            in1 => \N__10807\,
            in2 => \_gnd_net_\,
            in3 => \N__11274\,
            lcout => \transmit_module.n3678\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i8_3_lut_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__20683\,
            in1 => \N__10847\,
            in2 => \N__13486\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.n109\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.VGA_HS_66_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__11860\,
            in1 => \N__12416\,
            in2 => \N__14288\,
            in3 => \N__10838\,
            lcout => \ADV_HSYNC_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23302\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i7_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101100001000"
        )
    port map (
            in0 => \N__11252\,
            in1 => \N__20129\,
            in2 => \N__19721\,
            in3 => \N__11261\,
            lcout => \transmit_module.TX_ADDR_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23302\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_14_i7_3_lut_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__15141\,
            in1 => \N__15175\,
            in2 => \_gnd_net_\,
            in3 => \N__13499\,
            lcout => \transmit_module.n141\,
            ltout => \transmit_module.n141_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1651_4_lut_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__19607\,
            in1 => \N__20127\,
            in2 => \N__11516\,
            in3 => \N__15199\,
            lcout => n22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.VGA_VISIBLE_Y_64_LC_13_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14305\,
            in2 => \_gnd_net_\,
            in3 => \N__11801\,
            lcout => \transmit_module.VGA_VISIBLE_Y\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23302\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_14_i8_3_lut_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__15144\,
            in1 => \N__13482\,
            in2 => \_gnd_net_\,
            in3 => \N__13457\,
            lcout => \transmit_module.n140\,
            ltout => \transmit_module.n140_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1652_4_lut_LC_13_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__20128\,
            in1 => \N__19608\,
            in2 => \N__11255\,
            in3 => \N__11251\,
            lcout => n21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.VGA_VS_67_LC_13_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000110010"
        )
    port map (
            in0 => \N__11014\,
            in1 => \N__10988\,
            in2 => \N__10979\,
            in3 => \N__10963\,
            lcout => \ADV_VSYNC_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23302\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1732_4_lut_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100010001000"
        )
    port map (
            in0 => \N__11819\,
            in1 => \N__11856\,
            in2 => \N__10937\,
            in3 => \N__11872\,
            lcout => \transmit_module.video_signal_controller.n2975\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_14_i2_3_lut_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__14503\,
            in1 => \N__15126\,
            in2 => \_gnd_net_\,
            in3 => \N__13322\,
            lcout => \transmit_module.n146\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i4_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__20180\,
            in1 => \N__13616\,
            in2 => \N__19837\,
            in3 => \N__11789\,
            lcout => \transmit_module.TX_ADDR_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23488\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i5_LC_13_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__20193\,
            in1 => \N__12104\,
            in2 => \N__19722\,
            in3 => \N__12113\,
            lcout => \transmit_module.TX_ADDR_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23488\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_14_i6_3_lut_LC_13_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__15127\,
            in1 => \N__13534\,
            in2 => \N__13511\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.n142\,
            ltout => \transmit_module.n142_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1650_4_lut_LC_13_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__19612\,
            in1 => \N__20179\,
            in2 => \N__12107\,
            in3 => \N__12103\,
            lcout => n23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1764_4_lut_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010000000"
        )
    port map (
            in0 => \N__12434\,
            in1 => \N__11873\,
            in2 => \N__11861\,
            in3 => \N__11818\,
            lcout => \transmit_module.video_signal_controller.n3007\,
            ltout => \transmit_module.video_signal_controller.n3007_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i2_4_lut_adj_35_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__11555\,
            in1 => \N__12377\,
            in2 => \N__11804\,
            in3 => \N__11800\,
            lcout => \transmit_module.video_signal_controller.n7_adj_624\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i8_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__20195\,
            in1 => \N__12428\,
            in2 => \N__19866\,
            in3 => \N__12371\,
            lcout => \transmit_module.TX_ADDR_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23405\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_14_i5_3_lut_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__15119\,
            in1 => \_gnd_net_\,
            in2 => \N__13553\,
            in3 => \N__20806\,
            lcout => \transmit_module.n143\,
            ltout => \transmit_module.n143_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1649_4_lut_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__19723\,
            in1 => \N__20181\,
            in2 => \N__11783\,
            in3 => \N__13615\,
            lcout => n24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1774_3_lut_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__11554\,
            in1 => \N__12415\,
            in2 => \_gnd_net_\,
            in3 => \N__11522\,
            lcout => \transmit_module.video_signal_controller.n3017\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i509_2_lut_rep_20_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12484\,
            in2 => \_gnd_net_\,
            in3 => \N__12457\,
            lcout => \transmit_module.video_signal_controller.n3679\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i9_3_lut_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__14513\,
            in1 => \N__20661\,
            in2 => \_gnd_net_\,
            in3 => \N__14535\,
            lcout => \transmit_module.n108\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i2_2_lut_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14273\,
            in2 => \_gnd_net_\,
            in3 => \N__12408\,
            lcout => \transmit_module.video_signal_controller.n6_adj_623\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_14_i9_3_lut_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__15115\,
            in1 => \N__14534\,
            in2 => \_gnd_net_\,
            in3 => \N__13448\,
            lcout => \transmit_module.n139\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_14_i10_3_lut_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__14211\,
            in1 => \_gnd_net_\,
            in2 => \N__15143\,
            in3 => \N__13436\,
            lcout => \transmit_module.n138\,
            ltout => \transmit_module.n138_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1654_4_lut_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__19727\,
            in1 => \N__20194\,
            in2 => \N__12359\,
            in3 => \N__14176\,
            lcout => n19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_12__bdd_4_lut_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__22306\,
            in1 => \N__12140\,
            in2 => \N__23919\,
            in3 => \N__12131\,
            lcout => \line_buffer.n3620\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.i1144_1_lut_LC_13_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__15142\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.n2388\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i7_LC_13_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101000001100"
        )
    port map (
            in0 => \N__12743\,
            in1 => \N__12650\,
            in2 => \N__23933\,
            in3 => \N__12119\,
            lcout => \TX_DATA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23228\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2197_3_lut_LC_13_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__12776\,
            in1 => \N__12761\,
            in2 => \_gnd_net_\,
            in3 => \N__24780\,
            lcout => \line_buffer.n3534\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.VGA_R__i8_LC_13_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12737\,
            lcout => \ADV_B_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23257\,
            ce => 'H',
            sr => \N__22670\
        );

    \line_buffer.i2196_3_lut_LC_13_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__12677\,
            in1 => \N__12665\,
            in2 => \_gnd_net_\,
            in3 => \N__24798\,
            lcout => \line_buffer.n3533\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1_2_lut_3_lut_4_lut_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__14927\,
            in1 => \N__14828\,
            in2 => \N__14882\,
            in3 => \N__18682\,
            lcout => \line_buffer.n542\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i2_3_lut_adj_23_LC_14_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__12577\,
            in1 => \N__12565\,
            in2 => \_gnd_net_\,
            in3 => \N__12553\,
            lcout => \receive_module.rx_counter.n3225\,
            ltout => \receive_module.rx_counter.n3225_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i3_4_lut_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__12534\,
            in1 => \N__12988\,
            in2 => \N__12542\,
            in3 => \N__12969\,
            lcout => OPEN,
            ltout => \receive_module.rx_counter.n3458_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1_4_lut_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__12520\,
            in1 => \N__12951\,
            in2 => \N__12539\,
            in3 => \N__12852\,
            lcout => \receive_module.rx_counter.n39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1_2_lut_adj_24_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__12535\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12519\,
            lcout => \receive_module.rx_counter.n6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i5_1_lut_LC_14_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14335\,
            lcout => \receive_module.rx_counter.n3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i2_2_lut_adj_25_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12987\,
            in2 => \_gnd_net_\,
            in3 => \N__12970\,
            lcout => OPEN,
            ltout => \receive_module.rx_counter.n7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i2092_4_lut_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101000"
        )
    port map (
            in0 => \N__12952\,
            in1 => \N__12935\,
            in2 => \N__12929\,
            in3 => \N__12926\,
            lcout => \receive_module.rx_counter.n3429\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.old_HS_51_LC_14_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14344\,
            lcout => \receive_module.rx_counter.old_HS\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24123\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i252_3_lut_LC_14_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111101010101"
        )
    port map (
            in0 => \N__18862\,
            in1 => \_gnd_net_\,
            in2 => \N__14345\,
            in3 => \N__12920\,
            lcout => \receive_module.rx_counter.n2081\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1_2_lut_3_lut_4_lut_adj_19_LC_14_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__14867\,
            in1 => \N__18662\,
            in2 => \N__14827\,
            in3 => \N__14923\,
            lcout => \line_buffer.n573\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i609_2_lut_rep_21_LC_14_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12811\,
            in2 => \_gnd_net_\,
            in3 => \N__12792\,
            lcout => \receive_module.rx_counter.n3680\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i58_4_lut_LC_14_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000100000001"
        )
    port map (
            in0 => \N__12860\,
            in1 => \N__12853\,
            in2 => \N__12836\,
            in3 => \N__12821\,
            lcout => \receive_module.rx_counter.n54\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1_2_lut_3_lut_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__13304\,
            in1 => \N__12810\,
            in2 => \_gnd_net_\,
            in3 => \N__12793\,
            lcout => OPEN,
            ltout => \receive_module.rx_counter.n5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i3_4_lut_adj_21_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__13262\,
            in1 => \N__13088\,
            in2 => \N__13313\,
            in3 => \N__13145\,
            lcout => \receive_module.rx_counter.n3481\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i2_4_lut_LC_14_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101100"
        )
    port map (
            in0 => \N__13218\,
            in1 => \N__13133\,
            in2 => \N__13198\,
            in3 => \N__13163\,
            lcout => OPEN,
            ltout => \receive_module.rx_counter.n3455_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1_4_lut_adj_22_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010000000"
        )
    port map (
            in0 => \N__13114\,
            in1 => \N__13305\,
            in2 => \N__13286\,
            in3 => \N__13279\,
            lcout => OPEN,
            ltout => \receive_module.rx_counter.n4_adj_612_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.O_VISIBLE_53_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001001100"
        )
    port map (
            in0 => \N__13263\,
            in1 => \N__13238\,
            in2 => \N__13232\,
            in3 => \N__13229\,
            lcout => \DEBUG_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24128\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i2_3_lut_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__13217\,
            in1 => \N__13193\,
            in2 => \_gnd_net_\,
            in3 => \N__13164\,
            lcout => \receive_module.rx_counter.n3453\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1_2_lut_adj_27_LC_14_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__13134\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13109\,
            lcout => \receive_module.rx_counter.n4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sync_buffer.BUFFER_0__i1_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__13082\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \sync_buffer.BUFFER_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23531\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1_2_lut_3_lut_4_lut_adj_18_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__14922\,
            in1 => \N__14879\,
            in2 => \N__14821\,
            in3 => \N__18661\,
            lcout => \line_buffer.n477\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1_2_lut_3_lut_4_lut_adj_14_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__14880\,
            in1 => \N__18659\,
            in2 => \N__14825\,
            in3 => \N__14920\,
            lcout => \line_buffer.n541\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1_2_lut_3_lut_4_lut_adj_15_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__14921\,
            in1 => \N__14881\,
            in2 => \N__14822\,
            in3 => \N__18660\,
            lcout => \line_buffer.n605\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i2_3_lut_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__20162\,
            in1 => \N__19694\,
            in2 => \_gnd_net_\,
            in3 => \N__15145\,
            lcout => \transmit_module.n2087\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2215_3_lut_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__13370\,
            in1 => \N__13352\,
            in2 => \_gnd_net_\,
            in3 => \N__24715\,
            lcout => \line_buffer.n3552\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sync_buffer.BUFFER_0__i2_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13337\,
            lcout => \sync_buffer.BUFFER_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23666\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i0_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101100001000"
        )
    port map (
            in0 => \N__14144\,
            in1 => \N__20163\,
            in2 => \N__19836\,
            in3 => \N__14129\,
            lcout => \transmit_module.TX_ADDR_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23666\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i7_3_lut_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__20676\,
            in1 => \N__13331\,
            in2 => \_gnd_net_\,
            in3 => \N__15173\,
            lcout => \transmit_module.n110\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1_3_lut_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__19693\,
            in1 => \N__20677\,
            in2 => \_gnd_net_\,
            in3 => \N__20161\,
            lcout => \transmit_module.n2313\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_2_lut_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14450\,
            in2 => \N__14671\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.n132\,
            ltout => OPEN,
            carryin => \bfn_14_15_0_\,
            carryout => \transmit_module.n3162\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_3_lut_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14492\,
            in2 => \_gnd_net_\,
            in3 => \N__13316\,
            lcout => \transmit_module.n131\,
            ltout => OPEN,
            carryin => \transmit_module.n3162\,
            carryout => \transmit_module.n3163\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_4_lut_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20573\,
            in2 => \_gnd_net_\,
            in3 => \N__13559\,
            lcout => \transmit_module.n130\,
            ltout => OPEN,
            carryin => \transmit_module.n3163\,
            carryout => \transmit_module.n3164\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_5_lut_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16404\,
            in3 => \N__13556\,
            lcout => \transmit_module.n129\,
            ltout => OPEN,
            carryin => \transmit_module.n3164\,
            carryout => \transmit_module.n3165\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_6_lut_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20804\,
            in2 => \_gnd_net_\,
            in3 => \N__13541\,
            lcout => \transmit_module.n128\,
            ltout => OPEN,
            carryin => \transmit_module.n3165\,
            carryout => \transmit_module.n3166\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_7_lut_LC_14_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13532\,
            in2 => \_gnd_net_\,
            in3 => \N__13502\,
            lcout => \transmit_module.n127\,
            ltout => OPEN,
            carryin => \transmit_module.n3166\,
            carryout => \transmit_module.n3167\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_8_lut_LC_14_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15174\,
            in3 => \N__13493\,
            lcout => \transmit_module.n126\,
            ltout => OPEN,
            carryin => \transmit_module.n3167\,
            carryout => \transmit_module.n3168\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_9_lut_LC_14_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13478\,
            in2 => \_gnd_net_\,
            in3 => \N__13451\,
            lcout => \transmit_module.n125\,
            ltout => OPEN,
            carryin => \transmit_module.n3168\,
            carryout => \transmit_module.n3169\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_10_lut_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14539\,
            in3 => \N__13439\,
            lcout => \transmit_module.n124\,
            ltout => OPEN,
            carryin => \bfn_14_16_0_\,
            carryout => \transmit_module.n3170\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_11_lut_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14210\,
            in3 => \N__13424\,
            lcout => \transmit_module.n123\,
            ltout => OPEN,
            carryin => \transmit_module.n3170\,
            carryout => \transmit_module.n3171\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_12_lut_LC_14_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14578\,
            in3 => \N__13421\,
            lcout => \transmit_module.n122\,
            ltout => OPEN,
            carryin => \transmit_module.n3171\,
            carryout => \transmit_module.n3172\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_13_lut_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24732\,
            in2 => \_gnd_net_\,
            in3 => \N__13646\,
            lcout => \transmit_module.n121\,
            ltout => OPEN,
            carryin => \transmit_module.n3172\,
            carryout => \transmit_module.n3173\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_14_lut_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22305\,
            in2 => \_gnd_net_\,
            in3 => \N__13634\,
            lcout => \transmit_module.n120\,
            ltout => OPEN,
            carryin => \transmit_module.n3173\,
            carryout => \transmit_module.n3174\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.add_13_15_lut_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23917\,
            in2 => \_gnd_net_\,
            in3 => \N__13631\,
            lcout => \transmit_module.n119\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i5_3_lut_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__20672\,
            in1 => \N__20783\,
            in2 => \_gnd_net_\,
            in3 => \N__20805\,
            lcout => \transmit_module.n112\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i1_LC_14_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__20261\,
            in1 => \N__14164\,
            in2 => \N__19838\,
            in3 => \N__13600\,
            lcout => \transmit_module.TX_ADDR_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23560\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sync_buffer.WIRE_OUT_0__9_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13586\,
            lcout => \RX_TX_SYNC_BUFF\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23376\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_14_i11_3_lut_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__15096\,
            in1 => \N__14573\,
            in2 => \_gnd_net_\,
            in3 => \N__13568\,
            lcout => \transmit_module.n137\,
            ltout => \transmit_module.n137_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i10_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000110000"
        )
    port map (
            in0 => \N__13895\,
            in1 => \N__19739\,
            in2 => \N__13562\,
            in3 => \N__20262\,
            lcout => \transmit_module.TX_ADDR_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23376\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i9_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__20263\,
            in1 => \N__14180\,
            in2 => \N__19875\,
            in3 => \N__14324\,
            lcout => \transmit_module.TX_ADDR_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23376\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.video_signal_controller.VGA_VISIBLE_65_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__14312\,
            in1 => \N__14294\,
            in2 => \N__14287\,
            in3 => \N__14240\,
            lcout => \transmit_module.VGA_VISIBLE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23376\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_14_i1_3_lut_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__15097\,
            in1 => \N__14234\,
            in2 => \_gnd_net_\,
            in3 => \N__14460\,
            lcout => \transmit_module.n147\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i11_3_lut_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__20625\,
            in1 => \N__14549\,
            in2 => \_gnd_net_\,
            in3 => \N__14574\,
            lcout => \transmit_module.n106\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i10_3_lut_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__20671\,
            in1 => \N__14225\,
            in2 => \_gnd_net_\,
            in3 => \N__14212\,
            lcout => \transmit_module.n107\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i2_3_lut_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__20647\,
            in1 => \N__14471\,
            in2 => \_gnd_net_\,
            in3 => \N__14502\,
            lcout => \transmit_module.n115\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_12_i1_3_lut_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__14435\,
            in1 => \N__20648\,
            in2 => \_gnd_net_\,
            in3 => \N__14461\,
            lcout => \transmit_module.n116\,
            ltout => \transmit_module.n116_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1640_4_lut_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000101000000"
        )
    port map (
            in0 => \N__19873\,
            in1 => \N__20236\,
            in2 => \N__14132\,
            in3 => \N__14125\,
            lcout => n28,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1655_4_lut_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001100100000"
        )
    port map (
            in0 => \N__13894\,
            in1 => \N__19874\,
            in2 => \N__20260\,
            in3 => \N__13883\,
            lcout => n18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.ADDR_Y_COMPONENT__i10_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14579\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23417\,
            ce => \N__20748\,
            sr => \N__20058\
        );

    \transmit_module.ADDR_Y_COMPONENT__i8_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14540\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23417\,
            ce => \N__20748\,
            sr => \N__20058\
        );

    \transmit_module.ADDR_Y_COMPONENT__i1_LC_14_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14504\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23417\,
            ce => \N__20748\,
            sr => \N__20058\
        );

    \transmit_module.ADDR_Y_COMPONENT__i0_LC_14_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14465\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23417\,
            ce => \N__20748\,
            sr => \N__20058\
        );

    \tvp_vs_buffer.BUFFER_0__i1_LC_15_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14413\,
            lcout => \tvp_vs_buffer.BUFFER_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24100\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.BUFFER_0__i5_LC_15_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14389\,
            lcout => \tvp_video_buffer.BUFFER_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24106\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_vs_buffer.BUFFER_0__i2_LC_15_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14360\,
            lcout => \tvp_vs_buffer.BUFFER_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24106\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.BUFFER_0__i13_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14351\,
            lcout => \tvp_video_buffer.BUFFER_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24111\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_hs_buffer.WIRE_OUT_0__9_LC_15_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20849\,
            lcout => \TVP_HSYNC_buff\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24111\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.X_DELTA_PATTERN_i10_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14615\,
            lcout => \transmit_module.X_DELTA_PATTERN_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23551\,
            ce => \N__21476\,
            sr => \N__21362\
        );

    \transmit_module.X_DELTA_PATTERN_i9_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14627\,
            lcout => \transmit_module.X_DELTA_PATTERN_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23551\,
            ce => \N__21476\,
            sr => \N__21362\
        );

    \transmit_module.X_DELTA_PATTERN_i8_LC_15_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14621\,
            lcout => \transmit_module.X_DELTA_PATTERN_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23551\,
            ce => \N__21476\,
            sr => \N__21362\
        );

    \transmit_module.X_DELTA_PATTERN_i11_LC_15_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14597\,
            lcout => \transmit_module.X_DELTA_PATTERN_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23551\,
            ce => \N__21476\,
            sr => \N__21362\
        );

    \transmit_module.X_DELTA_PATTERN_i12_LC_15_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14609\,
            lcout => \transmit_module.X_DELTA_PATTERN_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23551\,
            ce => \N__21476\,
            sr => \N__21362\
        );

    \receive_module.add_12_2_lut_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18099\,
            in2 => \_gnd_net_\,
            in3 => \N__14591\,
            lcout => \receive_module.n137\,
            ltout => OPEN,
            carryin => \bfn_15_11_0_\,
            carryout => \receive_module.n3149\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_3_lut_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15540\,
            in2 => \_gnd_net_\,
            in3 => \N__14588\,
            lcout => \receive_module.n136\,
            ltout => OPEN,
            carryin => \receive_module.n3149\,
            carryout => \receive_module.n3150\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_4_lut_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15288\,
            in2 => \_gnd_net_\,
            in3 => \N__14585\,
            lcout => \receive_module.n135\,
            ltout => OPEN,
            carryin => \receive_module.n3150\,
            carryout => \receive_module.n3151\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_5_lut_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17862\,
            in2 => \_gnd_net_\,
            in3 => \N__14582\,
            lcout => \receive_module.n134\,
            ltout => OPEN,
            carryin => \receive_module.n3151\,
            carryout => \receive_module.n3152\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_6_lut_LC_15_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17244\,
            in2 => \_gnd_net_\,
            in3 => \N__14654\,
            lcout => \receive_module.n133\,
            ltout => OPEN,
            carryin => \receive_module.n3152\,
            carryout => \receive_module.n3153\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_7_lut_LC_15_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16992\,
            in2 => \_gnd_net_\,
            in3 => \N__14651\,
            lcout => \receive_module.n132\,
            ltout => OPEN,
            carryin => \receive_module.n3153\,
            carryout => \receive_module.n3154\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_8_lut_LC_15_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16725\,
            in2 => \_gnd_net_\,
            in3 => \N__14648\,
            lcout => \receive_module.n131\,
            ltout => OPEN,
            carryin => \receive_module.n3154\,
            carryout => \receive_module.n3155\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_9_lut_LC_15_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16464\,
            in2 => \_gnd_net_\,
            in3 => \N__14645\,
            lcout => \receive_module.n130\,
            ltout => OPEN,
            carryin => \receive_module.n3155\,
            carryout => \receive_module.n3156\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_10_lut_LC_15_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15828\,
            in2 => \_gnd_net_\,
            in3 => \N__14642\,
            lcout => \receive_module.n129\,
            ltout => OPEN,
            carryin => \bfn_15_12_0_\,
            carryout => \receive_module.n3157\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_11_lut_LC_15_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16173\,
            in2 => \_gnd_net_\,
            in3 => \N__14639\,
            lcout => \receive_module.n128\,
            ltout => OPEN,
            carryin => \receive_module.n3157\,
            carryout => \receive_module.n3158\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.add_12_12_lut_LC_15_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17625\,
            in2 => \_gnd_net_\,
            in3 => \N__14636\,
            lcout => \receive_module.n127\,
            ltout => OPEN,
            carryin => \receive_module.n3158\,
            carryout => \receive_module.n3159\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.BRAM_ADDR__i11_LC_15_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14916\,
            in2 => \_gnd_net_\,
            in3 => \N__14633\,
            lcout => \RX_ADDR_11\,
            ltout => OPEN,
            carryin => \receive_module.n3159\,
            carryout => \receive_module.n3160\,
            clk => \N__24124\,
            ce => \N__14939\,
            sr => \N__17513\
        );

    \receive_module.BRAM_ADDR__i12_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14868\,
            in2 => \_gnd_net_\,
            in3 => \N__14630\,
            lcout => \RX_ADDR_12\,
            ltout => OPEN,
            carryin => \receive_module.n3160\,
            carryout => \receive_module.n3161\,
            clk => \N__24124\,
            ce => \N__14939\,
            sr => \N__17513\
        );

    \receive_module.BRAM_ADDR__i13_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14817\,
            in2 => \_gnd_net_\,
            in3 => \N__15038\,
            lcout => \RX_ADDR_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24124\,
            ce => \N__14939\,
            sr => \N__17513\
        );

    \tvp_vs_buffer.WIRE_OUT_0__9_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14681\,
            lcout => \TVP_VSYNC_buff\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24129\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1_2_lut_3_lut_4_lut_adj_16_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__14918\,
            in1 => \N__14865\,
            in2 => \N__14823\,
            in3 => \N__18663\,
            lcout => \line_buffer.n606\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1_2_lut_3_lut_4_lut_adj_17_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__18665\,
            in1 => \N__14864\,
            in2 => \N__14826\,
            in3 => \N__14917\,
            lcout => \line_buffer.n476\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.O_VS_I_0_1_lut_rep_18_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18843\,
            lcout => \receive_module.n3677\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i249_2_lut_rep_15_2_lut_LC_15_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__18844\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18669\,
            lcout => \receive_module.n3674\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i1_2_lut_3_lut_4_lut_adj_20_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__14919\,
            in1 => \N__14866\,
            in2 => \N__14824\,
            in3 => \N__18664\,
            lcout => \line_buffer.n574\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_vs_buffer.BUFFER_0__i3_LC_15_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14693\,
            lcout => \tvp_vs_buffer.BUFFER_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24129\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.X_DELTA_PATTERN_i0_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15245\,
            lcout => \transmit_module.X_DELTA_PATTERN_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23409\,
            ce => \N__21464\,
            sr => \N__21327\
        );

    \transmit_module.X_DELTA_PATTERN_i1_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15230\,
            lcout => \transmit_module.X_DELTA_PATTERN_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23409\,
            ce => \N__21464\,
            sr => \N__21327\
        );

    \transmit_module.X_DELTA_PATTERN_i7_LC_15_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15239\,
            lcout => \transmit_module.X_DELTA_PATTERN_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23409\,
            ce => \N__21464\,
            sr => \N__21327\
        );

    \transmit_module.X_DELTA_PATTERN_i2_LC_15_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15224\,
            lcout => \transmit_module.X_DELTA_PATTERN_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23409\,
            ce => \N__21464\,
            sr => \N__21327\
        );

    \transmit_module.X_DELTA_PATTERN_i3_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15212\,
            lcout => \transmit_module.X_DELTA_PATTERN_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23409\,
            ce => \N__21464\,
            sr => \N__21327\
        );

    \transmit_module.X_DELTA_PATTERN_i6_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15218\,
            lcout => \transmit_module.X_DELTA_PATTERN_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23409\,
            ce => \N__21464\,
            sr => \N__21327\
        );

    \transmit_module.X_DELTA_PATTERN_i4_LC_15_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21485\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \transmit_module.X_DELTA_PATTERN_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23409\,
            ce => \N__21464\,
            sr => \N__21327\
        );

    \transmit_module.mux_14_i4_3_lut_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__15206\,
            in1 => \N__15140\,
            in2 => \_gnd_net_\,
            in3 => \N__16397\,
            lcout => \transmit_module.n144\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i6_LC_15_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__20254\,
            in1 => \N__15200\,
            in2 => \N__19951\,
            in3 => \N__15188\,
            lcout => \transmit_module.TX_ADDR_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23383\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.mux_14_i3_3_lut_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__20577\,
            in1 => \N__15114\,
            in2 => \_gnd_net_\,
            in3 => \N__15044\,
            lcout => \transmit_module.n145\,
            ltout => \transmit_module.n145_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i2_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010000010000"
        )
    port map (
            in0 => \N__20037\,
            in1 => \N__20255\,
            in2 => \N__15785\,
            in3 => \N__20552\,
            lcout => \transmit_module.TX_ADDR_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23133\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.BRAM_ADDR__i3_LC_15_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__20256\,
            in1 => \N__19517\,
            in2 => \N__20066\,
            in3 => \N__19495\,
            lcout => \transmit_module.TX_ADDR_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23133\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.Y_DELTA_PATTERN_i1_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15782\,
            lcout => \transmit_module.Y_DELTA_PATTERN_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23404\,
            ce => \N__21406\,
            sr => \N__20041\
        );

    \transmit_module.Y_DELTA_PATTERN_i2_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15761\,
            lcout => \transmit_module.Y_DELTA_PATTERN_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23404\,
            ce => \N__21406\,
            sr => \N__20041\
        );

    \transmit_module.Y_DELTA_PATTERN_i4_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15776\,
            lcout => \transmit_module.Y_DELTA_PATTERN_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23404\,
            ce => \N__21406\,
            sr => \N__20041\
        );

    \transmit_module.Y_DELTA_PATTERN_i3_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15767\,
            lcout => \transmit_module.Y_DELTA_PATTERN_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23404\,
            ce => \N__21406\,
            sr => \N__20041\
        );

    \transmit_module.Y_DELTA_PATTERN_i0_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1001",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15755\,
            lcout => \transmit_module.Y_DELTA_PATTERN_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23232\,
            ce => \N__21405\,
            sr => \N__19912\
        );

    \receive_module.BRAM_ADDR__i1_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111011000100"
        )
    port map (
            in0 => \N__18892\,
            in1 => \N__15749\,
            in2 => \N__18753\,
            in3 => \N__15515\,
            lcout => \RX_ADDR_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24141\,
            ce => 'H',
            sr => \N__17542\
        );

    \receive_module.BRAM_ADDR__i2_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111010100010"
        )
    port map (
            in0 => \N__15491\,
            in1 => \N__18895\,
            in2 => \N__18754\,
            in3 => \N__15272\,
            lcout => \RX_ADDR_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24141\,
            ce => 'H',
            sr => \N__17542\
        );

    \receive_module.BRAM_ADDR__i4_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111011000100"
        )
    port map (
            in0 => \N__18893\,
            in1 => \N__17453\,
            in2 => \N__18755\,
            in3 => \N__17219\,
            lcout => \RX_ADDR_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24141\,
            ce => 'H',
            sr => \N__17542\
        );

    \receive_module.BRAM_ADDR__i5_LC_15_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__18896\,
            in1 => \N__17189\,
            in2 => \N__16976\,
            in3 => \N__18733\,
            lcout => \RX_ADDR_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24141\,
            ce => 'H',
            sr => \N__17542\
        );

    \receive_module.BRAM_ADDR__i6_LC_15_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100001000"
        )
    port map (
            in0 => \N__18894\,
            in1 => \N__16700\,
            in2 => \N__18756\,
            in3 => \N__16934\,
            lcout => \RX_ADDR_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24141\,
            ce => 'H',
            sr => \N__17542\
        );

    \receive_module.BRAM_ADDR__i7_LC_15_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100100000"
        )
    port map (
            in0 => \N__18897\,
            in1 => \N__18737\,
            in2 => \N__16457\,
            in3 => \N__16673\,
            lcout => \RX_ADDR_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24141\,
            ce => 'H',
            sr => \N__17542\
        );

    \transmit_module.mux_12_i4_3_lut_LC_15_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__20655\,
            in1 => \N__16418\,
            in2 => \_gnd_net_\,
            in3 => \N__16405\,
            lcout => \transmit_module.n113\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.BRAM_ADDR__i9_LC_15_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100001000"
        )
    port map (
            in0 => \N__18908\,
            in1 => \N__16145\,
            in2 => \N__18768\,
            in3 => \N__16373\,
            lcout => \RX_ADDR_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24146\,
            ce => 'H',
            sr => \N__17555\
        );

    \GB_BUFFER_DEBUG_c_3_c_THRU_LUT4_0_LC_15_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__24173\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \GB_BUFFER_DEBUG_c_3_c_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.VGA_R__i1_LC_15_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22070\,
            lcout => n1821,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22876\,
            ce => 'H',
            sr => \N__22688\
        );

    \receive_module.BRAM_ADDR__i8_LC_15_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100001000"
        )
    port map (
            in0 => \N__18918\,
            in1 => \N__15812\,
            in2 => \N__18777\,
            in3 => \N__16034\,
            lcout => \RX_ADDR_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24155\,
            ce => 'H',
            sr => \N__17565\
        );

    \receive_module.BRAM_ADDR__i0_LC_15_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111011000100"
        )
    port map (
            in0 => \N__18919\,
            in1 => \N__18302\,
            in2 => \N__18766\,
            in3 => \N__18080\,
            lcout => \RX_ADDR_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24157\,
            ce => 'H',
            sr => \N__17566\
        );

    \receive_module.BRAM_ADDR__i3_LC_15_31_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111011000100"
        )
    port map (
            in0 => \N__18926\,
            in1 => \N__18056\,
            in2 => \N__18785\,
            in3 => \N__17846\,
            lcout => \RX_ADDR_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24161\,
            ce => 'H',
            sr => \N__17570\
        );

    \receive_module.BRAM_ADDR__i10_LC_15_31_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110100001000"
        )
    port map (
            in0 => \N__18925\,
            in1 => \N__17597\,
            in2 => \N__18784\,
            in3 => \N__17822\,
            lcout => \RX_ADDR_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24161\,
            ce => 'H',
            sr => \N__17570\
        );

    \PULSE_1HZ_I_0_2_lut_LC_16_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__18805\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17477\,
            lcout => \LED_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.PULSE_1HZ_49_LC_16_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17473\,
            in2 => \_gnd_net_\,
            in3 => \N__18428\,
            lcout => \PULSE_1HZ\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24103\,
            ce => \N__18326\,
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1_2_lut_adj_26_LC_16_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18355\,
            in2 => \_gnd_net_\,
            in3 => \N__18385\,
            lcout => \receive_module.rx_counter.n7_adj_619\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i134_2_lut_rep_16_2_lut_LC_16_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__18871\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17462\,
            lcout => \receive_module.rx_counter.n3675\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i1307_2_lut_3_lut_3_lut_LC_16_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__17461\,
            in1 => \N__18870\,
            in2 => \_gnd_net_\,
            in3 => \N__18427\,
            lcout => \receive_module.rx_counter.n2550\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.old_VS_52_LC_16_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__18872\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \receive_module.rx_counter.old_VS\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24107\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i2185_2_lut_LC_16_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18400\,
            in2 => \_gnd_net_\,
            in3 => \N__18337\,
            lcout => OPEN,
            ltout => \receive_module.rx_counter.n3522_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.i5_4_lut_LC_16_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111111"
        )
    port map (
            in0 => \N__18415\,
            in1 => \N__18370\,
            in2 => \N__18437\,
            in3 => \N__18434\,
            lcout => \receive_module.rx_counter.n11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.rx_counter.FRAME_COUNTER_247__i0_LC_16_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18416\,
            in2 => \_gnd_net_\,
            in3 => \N__18404\,
            lcout => \receive_module.rx_counter.FRAME_COUNTER_0\,
            ltout => OPEN,
            carryin => \bfn_16_10_0_\,
            carryout => \receive_module.rx_counter.n3205\,
            clk => \N__24112\,
            ce => \N__18325\,
            sr => \N__19163\
        );

    \receive_module.rx_counter.FRAME_COUNTER_247__i1_LC_16_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18401\,
            in2 => \_gnd_net_\,
            in3 => \N__18389\,
            lcout => \receive_module.rx_counter.FRAME_COUNTER_1\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3205\,
            carryout => \receive_module.rx_counter.n3206\,
            clk => \N__24112\,
            ce => \N__18325\,
            sr => \N__19163\
        );

    \receive_module.rx_counter.FRAME_COUNTER_247__i2_LC_16_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18386\,
            in2 => \_gnd_net_\,
            in3 => \N__18374\,
            lcout => \receive_module.rx_counter.FRAME_COUNTER_2\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3206\,
            carryout => \receive_module.rx_counter.n3207\,
            clk => \N__24112\,
            ce => \N__18325\,
            sr => \N__19163\
        );

    \receive_module.rx_counter.FRAME_COUNTER_247__i3_LC_16_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18371\,
            in2 => \_gnd_net_\,
            in3 => \N__18359\,
            lcout => \receive_module.rx_counter.FRAME_COUNTER_3\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3207\,
            carryout => \receive_module.rx_counter.n3208\,
            clk => \N__24112\,
            ce => \N__18325\,
            sr => \N__19163\
        );

    \receive_module.rx_counter.FRAME_COUNTER_247__i4_LC_16_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18356\,
            in2 => \_gnd_net_\,
            in3 => \N__18344\,
            lcout => \receive_module.rx_counter.FRAME_COUNTER_4\,
            ltout => OPEN,
            carryin => \receive_module.rx_counter.n3208\,
            carryout => \receive_module.rx_counter.n3209\,
            clk => \N__24112\,
            ce => \N__18325\,
            sr => \N__19163\
        );

    \receive_module.rx_counter.FRAME_COUNTER_247__i5_LC_16_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18338\,
            in2 => \_gnd_net_\,
            in3 => \N__18341\,
            lcout => \receive_module.rx_counter.FRAME_COUNTER_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24112\,
            ce => \N__18325\,
            sr => \N__19163\
        );

    \tvp_video_buffer.WIRE_OUT_i4_LC_16_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19157\,
            lcout => \RX_DATA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24116\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.sync_wd.i2_2_lut_LC_16_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19081\,
            in2 => \_gnd_net_\,
            in3 => \N__18525\,
            lcout => OPEN,
            ltout => \receive_module.sync_wd.n6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.sync_wd.i1_4_lut_LC_16_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000001"
        )
    port map (
            in0 => \N__18959\,
            in1 => \N__22456\,
            in2 => \N__18932\,
            in3 => \N__18680\,
            lcout => OPEN,
            ltout => \receive_module.sync_wd.n4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.sync_wd.SYNC_BAD_16_LC_16_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100111000000000"
        )
    port map (
            in0 => \N__18602\,
            in1 => \N__18798\,
            in2 => \N__18929\,
            in3 => \N__18854\,
            lcout => \DEBUG_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24119\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \receive_module.sync_wd.old_visible_17_LC_16_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18681\,
            lcout => \receive_module.sync_wd.old_visible\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24119\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.WIRE_OUT_i7_LC_16_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22532\,
            lcout => \RX_DATA_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24125\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_LC_16_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__24764\,
            in1 => \N__18500\,
            in2 => \N__22376\,
            in3 => \N__18482\,
            lcout => \line_buffer.n3656\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_2260_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__24772\,
            in1 => \N__18467\,
            in2 => \N__22377\,
            in3 => \N__18449\,
            lcout => \line_buffer.n3590\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i1_LC_16_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__23940\,
            in1 => \N__21242\,
            in2 => \_gnd_net_\,
            in3 => \N__21209\,
            lcout => \TX_DATA_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22908\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.ADDR_Y_COMPONENT__i4_LC_16_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20810\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23132\,
            ce => \N__20757\,
            sr => \N__19911\
        );

    \transmit_module.ADDR_Y_COMPONENT__i2_LC_16_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20578\,
            lcout => \transmit_module.ADDR_Y_COMPONENT_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23375\,
            ce => \N__20771\,
            sr => \N__20042\
        );

    \transmit_module.mux_12_i3_3_lut_LC_16_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__20690\,
            in1 => \N__20626\,
            in2 => \_gnd_net_\,
            in3 => \N__20579\,
            lcout => \transmit_module.n114\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1647_4_lut_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110100001000"
        )
    port map (
            in0 => \N__20257\,
            in1 => \N__20548\,
            in2 => \N__20013\,
            in3 => \N__20537\,
            lcout => n26,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n3626_bdd_4_lut_LC_16_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__20306\,
            in1 => \N__22339\,
            in2 => \N__20285\,
            in3 => \N__21779\,
            lcout => \line_buffer.n3629\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.i1648_4_lut_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100100000"
        )
    port map (
            in0 => \N__20258\,
            in1 => \N__19910\,
            in2 => \N__19516\,
            in3 => \N__19499\,
            lcout => n25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.VGA_R__i4_LC_16_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21074\,
            lcout => n1818,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22987\,
            ce => 'H',
            sr => \N__22649\
        );

    \line_buffer.n3590_bdd_4_lut_LC_16_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__22375\,
            in1 => \N__19205\,
            in2 => \N__19193\,
            in3 => \N__19172\,
            lcout => OPEN,
            ltout => \line_buffer.n3593_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i3_LC_16_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23932\,
            in2 => \N__21086\,
            in3 => \N__21083\,
            lcout => \TX_DATA_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23201\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2214_3_lut_LC_16_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21068\,
            in1 => \N__21053\,
            in2 => \_gnd_net_\,
            in3 => \N__24797\,
            lcout => OPEN,
            ltout => \line_buffer.n3551_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i4_LC_16_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__23938\,
            in1 => \N__21035\,
            in2 => \N__21020\,
            in3 => \N__21692\,
            lcout => \TX_DATA_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23039\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2200_3_lut_LC_16_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__24796\,
            in1 => \N__21017\,
            in2 => \_gnd_net_\,
            in3 => \N__20996\,
            lcout => \line_buffer.n3537\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.VGA_R__i5_LC_16_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20978\,
            lcout => n1817,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23125\,
            ce => 'H',
            sr => \N__22680\
        );

    \transmit_module.VGA_R__i2_LC_16_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20906\,
            lcout => n1820,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__22869\,
            ce => 'H',
            sr => \N__22692\
        );

    \tvp_hs_buffer.BUFFER_0__i2_LC_17_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21608\,
            lcout => \tvp_hs_buffer.BUFFER_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24101\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2199_3_lut_LC_17_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__24794\,
            in1 => \N__20840\,
            in2 => \_gnd_net_\,
            in3 => \N__20822\,
            lcout => \line_buffer.n3536\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2235_3_lut_LC_17_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__24795\,
            in1 => \N__21521\,
            in2 => \_gnd_net_\,
            in3 => \N__21503\,
            lcout => \line_buffer.n3572\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.X_DELTA_PATTERN_i5_LC_17_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21494\,
            lcout => \transmit_module.X_DELTA_PATTERN_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23487\,
            ce => \N__21474\,
            sr => \N__21354\
        );

    \line_buffer.n3650_bdd_4_lut_LC_17_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__21278\,
            in1 => \N__22346\,
            in2 => \N__21260\,
            in3 => \N__21878\,
            lcout => \line_buffer.n3653\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n3632_bdd_4_lut_LC_17_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__21236\,
            in1 => \N__21149\,
            in2 => \N__21224\,
            in3 => \N__22350\,
            lcout => \line_buffer.n3635\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2233_3_lut_LC_17_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21203\,
            in1 => \N__21185\,
            in2 => \_gnd_net_\,
            in3 => \N__24686\,
            lcout => \line_buffer.n3570\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_2294_LC_17_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__24745\,
            in1 => \N__21176\,
            in2 => \N__22372\,
            in3 => \N__21167\,
            lcout => \line_buffer.n3632\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_12__bdd_4_lut_2269_LC_17_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__22337\,
            in1 => \N__21566\,
            in2 => \N__23950\,
            in3 => \N__21143\,
            lcout => OPEN,
            ltout => \line_buffer.n3602_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i2_LC_17_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__23944\,
            in1 => \N__21656\,
            in2 => \N__21131\,
            in3 => \N__21128\,
            lcout => \TX_DATA_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23336\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n3656_bdd_4_lut_LC_17_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__21122\,
            in1 => \N__22338\,
            in2 => \N__21107\,
            in3 => \N__21818\,
            lcout => \line_buffer.n3659\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_2289_LC_17_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__24765\,
            in1 => \N__21806\,
            in2 => \N__22373\,
            in3 => \N__21791\,
            lcout => \line_buffer.n3626\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.VGA_R__i3_LC_17_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21773\,
            lcout => n1819,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23227\,
            ce => 'H',
            sr => \N__22687\
        );

    \line_buffer.TX_ADDR_12__bdd_4_lut_2279_LC_17_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__22374\,
            in1 => \N__21710\,
            in2 => \N__23949\,
            in3 => \N__21704\,
            lcout => \line_buffer.n3614\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2232_3_lut_LC_17_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21686\,
            in1 => \N__21674\,
            in2 => \_gnd_net_\,
            in3 => \N__24743\,
            lcout => \line_buffer.n3569\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_hs_buffer.BUFFER_0__i1_LC_18_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21628\,
            lcout => \tvp_hs_buffer.BUFFER_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24108\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2236_3_lut_LC_18_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__24763\,
            in1 => \N__21602\,
            in2 => \_gnd_net_\,
            in3 => \N__21587\,
            lcout => \line_buffer.n3573\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i5_LC_18_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__23939\,
            in1 => \N__21908\,
            in2 => \_gnd_net_\,
            in3 => \N__21560\,
            lcout => \TX_DATA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23570\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_2299_LC_18_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__24784\,
            in1 => \N__21554\,
            in2 => \N__22381\,
            in3 => \N__21536\,
            lcout => \line_buffer.n3638\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n3638_bdd_4_lut_LC_18_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__22124\,
            in1 => \N__22389\,
            in2 => \N__22109\,
            in3 => \N__22085\,
            lcout => \line_buffer.n3641\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i0_LC_18_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__23937\,
            in1 => \N__22076\,
            in2 => \_gnd_net_\,
            in3 => \N__22010\,
            lcout => \TX_DATA_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23439\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.n3644_bdd_4_lut_LC_18_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__22390\,
            in1 => \N__22058\,
            in2 => \N__22034\,
            in3 => \N__22577\,
            lcout => \line_buffer.n3647\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.VGA_R__i6_LC_18_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22004\,
            lcout => n1816,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23038\,
            ce => 'H',
            sr => \N__22694\
        );

    \line_buffer.n3596_bdd_4_lut_LC_19_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000110000"
        )
    port map (
            in0 => \N__21950\,
            in1 => \N__22391\,
            in2 => \N__21932\,
            in3 => \N__22175\,
            lcout => \line_buffer.n3599\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_2309_LC_19_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__24785\,
            in1 => \N__21902\,
            in2 => \N__22393\,
            in3 => \N__21893\,
            lcout => \line_buffer.n3650\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2239_3_lut_LC_19_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__24786\,
            in1 => \N__21866\,
            in2 => \_gnd_net_\,
            in3 => \N__21848\,
            lcout => \line_buffer.n3576\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_12__bdd_4_lut_2274_LC_19_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__22388\,
            in1 => \N__21827\,
            in2 => \N__23951\,
            in3 => \N__24530\,
            lcout => OPEN,
            ltout => \line_buffer.n3608_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.dout_i6_LC_19_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__23948\,
            in1 => \N__22541\,
            in2 => \N__23813\,
            in3 => \N__23810\,
            lcout => \TX_DATA_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23248\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \transmit_module.VGA_R__i7_LC_19_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23801\,
            lcout => n1815,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__23440\,
            ce => 'H',
            sr => \N__22693\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_2304_LC_19_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__24799\,
            in1 => \N__22613\,
            in2 => \N__22394\,
            in3 => \N__22598\,
            lcout => \line_buffer.n3644\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2238_3_lut_LC_19_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__22571\,
            in1 => \N__22556\,
            in2 => \_gnd_net_\,
            in3 => \N__24744\,
            lcout => \line_buffer.n3575\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.BUFFER_0__i16_LC_20_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__24185\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \tvp_video_buffer.BUFFER_1_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24132\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.WIRE_OUT_i5_LC_20_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24806\,
            lcout => \RX_DATA_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24139\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.TX_ADDR_11__bdd_4_lut_2284_LC_20_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__24793\,
            in1 => \N__22406\,
            in2 => \N__22392\,
            in3 => \N__22193\,
            lcout => \line_buffer.n3596\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.BUFFER_0__i6_LC_20_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22165\,
            lcout => \tvp_video_buffer.BUFFER_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24139\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.BUFFER_0__i14_LC_20_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24812\,
            lcout => \tvp_video_buffer.BUFFER_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24139\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \line_buffer.i2205_3_lut_LC_20_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__24800\,
            in1 => \N__24566\,
            in2 => \_gnd_net_\,
            in3 => \N__24551\,
            lcout => \line_buffer.n3542\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_22_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tvp_video_buffer.BUFFER_0__i8_LC_24_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__24194\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \tvp_video_buffer.BUFFER_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__24133\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
