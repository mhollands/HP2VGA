-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2017.08.27940

-- Build Date:         Sep 11 2017 17:29:57

-- File Generated:     Sep 9 2018 04:44:37

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "RAM" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of RAM
entity RAM is
port (
    raddr : in std_logic_vector(13 downto 0);
    waddr : in std_logic_vector(13 downto 0);
    dout : out std_logic_vector(7 downto 0);
    din : in std_logic_vector(7 downto 0);
    rclk : in std_logic;
    wclk : in std_logic;
    write_en : in std_logic);
end RAM;

-- Architecture of RAM
-- View name is \INTERFACE\
architecture \INTERFACE\ of RAM is

signal \N__13191\ : std_logic;
signal \N__13190\ : std_logic;
signal \N__13189\ : std_logic;
signal \N__13181\ : std_logic;
signal \N__13180\ : std_logic;
signal \N__13179\ : std_logic;
signal \N__13170\ : std_logic;
signal \N__13169\ : std_logic;
signal \N__13168\ : std_logic;
signal \N__13161\ : std_logic;
signal \N__13160\ : std_logic;
signal \N__13159\ : std_logic;
signal \N__13152\ : std_logic;
signal \N__13151\ : std_logic;
signal \N__13150\ : std_logic;
signal \N__13143\ : std_logic;
signal \N__13142\ : std_logic;
signal \N__13141\ : std_logic;
signal \N__13134\ : std_logic;
signal \N__13133\ : std_logic;
signal \N__13132\ : std_logic;
signal \N__13125\ : std_logic;
signal \N__13124\ : std_logic;
signal \N__13123\ : std_logic;
signal \N__13116\ : std_logic;
signal \N__13115\ : std_logic;
signal \N__13114\ : std_logic;
signal \N__13107\ : std_logic;
signal \N__13106\ : std_logic;
signal \N__13105\ : std_logic;
signal \N__13098\ : std_logic;
signal \N__13097\ : std_logic;
signal \N__13096\ : std_logic;
signal \N__13089\ : std_logic;
signal \N__13088\ : std_logic;
signal \N__13087\ : std_logic;
signal \N__13080\ : std_logic;
signal \N__13079\ : std_logic;
signal \N__13078\ : std_logic;
signal \N__13071\ : std_logic;
signal \N__13070\ : std_logic;
signal \N__13069\ : std_logic;
signal \N__13062\ : std_logic;
signal \N__13061\ : std_logic;
signal \N__13060\ : std_logic;
signal \N__13053\ : std_logic;
signal \N__13052\ : std_logic;
signal \N__13051\ : std_logic;
signal \N__13044\ : std_logic;
signal \N__13043\ : std_logic;
signal \N__13042\ : std_logic;
signal \N__13035\ : std_logic;
signal \N__13034\ : std_logic;
signal \N__13033\ : std_logic;
signal \N__13026\ : std_logic;
signal \N__13025\ : std_logic;
signal \N__13024\ : std_logic;
signal \N__13017\ : std_logic;
signal \N__13016\ : std_logic;
signal \N__13015\ : std_logic;
signal \N__13008\ : std_logic;
signal \N__13007\ : std_logic;
signal \N__13006\ : std_logic;
signal \N__12999\ : std_logic;
signal \N__12998\ : std_logic;
signal \N__12997\ : std_logic;
signal \N__12990\ : std_logic;
signal \N__12989\ : std_logic;
signal \N__12988\ : std_logic;
signal \N__12981\ : std_logic;
signal \N__12980\ : std_logic;
signal \N__12979\ : std_logic;
signal \N__12972\ : std_logic;
signal \N__12971\ : std_logic;
signal \N__12970\ : std_logic;
signal \N__12963\ : std_logic;
signal \N__12962\ : std_logic;
signal \N__12961\ : std_logic;
signal \N__12954\ : std_logic;
signal \N__12953\ : std_logic;
signal \N__12952\ : std_logic;
signal \N__12945\ : std_logic;
signal \N__12944\ : std_logic;
signal \N__12943\ : std_logic;
signal \N__12936\ : std_logic;
signal \N__12935\ : std_logic;
signal \N__12934\ : std_logic;
signal \N__12927\ : std_logic;
signal \N__12926\ : std_logic;
signal \N__12925\ : std_logic;
signal \N__12918\ : std_logic;
signal \N__12917\ : std_logic;
signal \N__12916\ : std_logic;
signal \N__12909\ : std_logic;
signal \N__12908\ : std_logic;
signal \N__12907\ : std_logic;
signal \N__12900\ : std_logic;
signal \N__12899\ : std_logic;
signal \N__12898\ : std_logic;
signal \N__12891\ : std_logic;
signal \N__12890\ : std_logic;
signal \N__12889\ : std_logic;
signal \N__12882\ : std_logic;
signal \N__12881\ : std_logic;
signal \N__12880\ : std_logic;
signal \N__12873\ : std_logic;
signal \N__12872\ : std_logic;
signal \N__12871\ : std_logic;
signal \N__12864\ : std_logic;
signal \N__12863\ : std_logic;
signal \N__12862\ : std_logic;
signal \N__12855\ : std_logic;
signal \N__12854\ : std_logic;
signal \N__12853\ : std_logic;
signal \N__12846\ : std_logic;
signal \N__12845\ : std_logic;
signal \N__12844\ : std_logic;
signal \N__12837\ : std_logic;
signal \N__12836\ : std_logic;
signal \N__12835\ : std_logic;
signal \N__12828\ : std_logic;
signal \N__12827\ : std_logic;
signal \N__12826\ : std_logic;
signal \N__12819\ : std_logic;
signal \N__12818\ : std_logic;
signal \N__12817\ : std_logic;
signal \N__12810\ : std_logic;
signal \N__12809\ : std_logic;
signal \N__12808\ : std_logic;
signal \N__12801\ : std_logic;
signal \N__12800\ : std_logic;
signal \N__12799\ : std_logic;
signal \N__12792\ : std_logic;
signal \N__12791\ : std_logic;
signal \N__12790\ : std_logic;
signal \N__12783\ : std_logic;
signal \N__12782\ : std_logic;
signal \N__12781\ : std_logic;
signal \N__12774\ : std_logic;
signal \N__12773\ : std_logic;
signal \N__12772\ : std_logic;
signal \N__12755\ : std_logic;
signal \N__12752\ : std_logic;
signal \N__12751\ : std_logic;
signal \N__12750\ : std_logic;
signal \N__12749\ : std_logic;
signal \N__12748\ : std_logic;
signal \N__12747\ : std_logic;
signal \N__12744\ : std_logic;
signal \N__12739\ : std_logic;
signal \N__12736\ : std_logic;
signal \N__12731\ : std_logic;
signal \N__12730\ : std_logic;
signal \N__12729\ : std_logic;
signal \N__12728\ : std_logic;
signal \N__12719\ : std_logic;
signal \N__12716\ : std_logic;
signal \N__12715\ : std_logic;
signal \N__12714\ : std_logic;
signal \N__12713\ : std_logic;
signal \N__12712\ : std_logic;
signal \N__12711\ : std_logic;
signal \N__12708\ : std_logic;
signal \N__12705\ : std_logic;
signal \N__12700\ : std_logic;
signal \N__12697\ : std_logic;
signal \N__12694\ : std_logic;
signal \N__12691\ : std_logic;
signal \N__12688\ : std_logic;
signal \N__12685\ : std_logic;
signal \N__12684\ : std_logic;
signal \N__12683\ : std_logic;
signal \N__12680\ : std_logic;
signal \N__12677\ : std_logic;
signal \N__12674\ : std_logic;
signal \N__12667\ : std_logic;
signal \N__12662\ : std_logic;
signal \N__12659\ : std_logic;
signal \N__12656\ : std_logic;
signal \N__12651\ : std_logic;
signal \N__12648\ : std_logic;
signal \N__12645\ : std_logic;
signal \N__12638\ : std_logic;
signal \N__12635\ : std_logic;
signal \N__12632\ : std_logic;
signal \N__12629\ : std_logic;
signal \N__12626\ : std_logic;
signal \N__12623\ : std_logic;
signal \N__12620\ : std_logic;
signal \N__12615\ : std_logic;
signal \N__12612\ : std_logic;
signal \N__12609\ : std_logic;
signal \N__12606\ : std_logic;
signal \N__12603\ : std_logic;
signal \N__12598\ : std_logic;
signal \N__12593\ : std_logic;
signal \N__12590\ : std_logic;
signal \N__12587\ : std_logic;
signal \N__12584\ : std_logic;
signal \N__12581\ : std_logic;
signal \N__12580\ : std_logic;
signal \N__12579\ : std_logic;
signal \N__12578\ : std_logic;
signal \N__12575\ : std_logic;
signal \N__12572\ : std_logic;
signal \N__12567\ : std_logic;
signal \N__12566\ : std_logic;
signal \N__12561\ : std_logic;
signal \N__12560\ : std_logic;
signal \N__12559\ : std_logic;
signal \N__12558\ : std_logic;
signal \N__12555\ : std_logic;
signal \N__12552\ : std_logic;
signal \N__12549\ : std_logic;
signal \N__12546\ : std_logic;
signal \N__12543\ : std_logic;
signal \N__12540\ : std_logic;
signal \N__12535\ : std_logic;
signal \N__12532\ : std_logic;
signal \N__12529\ : std_logic;
signal \N__12524\ : std_logic;
signal \N__12521\ : std_logic;
signal \N__12516\ : std_logic;
signal \N__12513\ : std_logic;
signal \N__12510\ : std_logic;
signal \N__12507\ : std_logic;
signal \N__12504\ : std_logic;
signal \N__12501\ : std_logic;
signal \N__12498\ : std_logic;
signal \N__12493\ : std_logic;
signal \N__12488\ : std_logic;
signal \N__12485\ : std_logic;
signal \N__12482\ : std_logic;
signal \N__12479\ : std_logic;
signal \N__12476\ : std_logic;
signal \N__12473\ : std_logic;
signal \N__12470\ : std_logic;
signal \N__12467\ : std_logic;
signal \N__12464\ : std_logic;
signal \N__12461\ : std_logic;
signal \N__12458\ : std_logic;
signal \N__12455\ : std_logic;
signal \N__12452\ : std_logic;
signal \N__12449\ : std_logic;
signal \N__12446\ : std_logic;
signal \N__12443\ : std_logic;
signal \N__12440\ : std_logic;
signal \N__12437\ : std_logic;
signal \N__12434\ : std_logic;
signal \N__12431\ : std_logic;
signal \N__12430\ : std_logic;
signal \N__12425\ : std_logic;
signal \N__12424\ : std_logic;
signal \N__12423\ : std_logic;
signal \N__12420\ : std_logic;
signal \N__12415\ : std_logic;
signal \N__12414\ : std_logic;
signal \N__12413\ : std_logic;
signal \N__12408\ : std_logic;
signal \N__12403\ : std_logic;
signal \N__12402\ : std_logic;
signal \N__12401\ : std_logic;
signal \N__12400\ : std_logic;
signal \N__12399\ : std_logic;
signal \N__12394\ : std_logic;
signal \N__12391\ : std_logic;
signal \N__12388\ : std_logic;
signal \N__12385\ : std_logic;
signal \N__12384\ : std_logic;
signal \N__12381\ : std_logic;
signal \N__12376\ : std_logic;
signal \N__12369\ : std_logic;
signal \N__12366\ : std_logic;
signal \N__12365\ : std_logic;
signal \N__12364\ : std_logic;
signal \N__12359\ : std_logic;
signal \N__12358\ : std_logic;
signal \N__12357\ : std_logic;
signal \N__12354\ : std_logic;
signal \N__12351\ : std_logic;
signal \N__12350\ : std_logic;
signal \N__12349\ : std_logic;
signal \N__12346\ : std_logic;
signal \N__12345\ : std_logic;
signal \N__12342\ : std_logic;
signal \N__12339\ : std_logic;
signal \N__12336\ : std_logic;
signal \N__12335\ : std_logic;
signal \N__12330\ : std_logic;
signal \N__12329\ : std_logic;
signal \N__12328\ : std_logic;
signal \N__12327\ : std_logic;
signal \N__12322\ : std_logic;
signal \N__12321\ : std_logic;
signal \N__12320\ : std_logic;
signal \N__12315\ : std_logic;
signal \N__12314\ : std_logic;
signal \N__12313\ : std_logic;
signal \N__12306\ : std_logic;
signal \N__12303\ : std_logic;
signal \N__12300\ : std_logic;
signal \N__12297\ : std_logic;
signal \N__12294\ : std_logic;
signal \N__12291\ : std_logic;
signal \N__12290\ : std_logic;
signal \N__12289\ : std_logic;
signal \N__12286\ : std_logic;
signal \N__12283\ : std_logic;
signal \N__12280\ : std_logic;
signal \N__12279\ : std_logic;
signal \N__12278\ : std_logic;
signal \N__12275\ : std_logic;
signal \N__12270\ : std_logic;
signal \N__12265\ : std_logic;
signal \N__12264\ : std_logic;
signal \N__12263\ : std_logic;
signal \N__12258\ : std_logic;
signal \N__12253\ : std_logic;
signal \N__12248\ : std_logic;
signal \N__12245\ : std_logic;
signal \N__12240\ : std_logic;
signal \N__12235\ : std_logic;
signal \N__12232\ : std_logic;
signal \N__12229\ : std_logic;
signal \N__12226\ : std_logic;
signal \N__12221\ : std_logic;
signal \N__12218\ : std_logic;
signal \N__12215\ : std_logic;
signal \N__12212\ : std_logic;
signal \N__12209\ : std_logic;
signal \N__12206\ : std_logic;
signal \N__12203\ : std_logic;
signal \N__12200\ : std_logic;
signal \N__12197\ : std_logic;
signal \N__12192\ : std_logic;
signal \N__12189\ : std_logic;
signal \N__12186\ : std_logic;
signal \N__12183\ : std_logic;
signal \N__12178\ : std_logic;
signal \N__12175\ : std_logic;
signal \N__12170\ : std_logic;
signal \N__12165\ : std_logic;
signal \N__12160\ : std_logic;
signal \N__12155\ : std_logic;
signal \N__12150\ : std_logic;
signal \N__12143\ : std_logic;
signal \N__12140\ : std_logic;
signal \N__12137\ : std_logic;
signal \N__12134\ : std_logic;
signal \N__12131\ : std_logic;
signal \N__12128\ : std_logic;
signal \N__12125\ : std_logic;
signal \N__12122\ : std_logic;
signal \N__12119\ : std_logic;
signal \N__12116\ : std_logic;
signal \N__12113\ : std_logic;
signal \N__12110\ : std_logic;
signal \N__12107\ : std_logic;
signal \N__12104\ : std_logic;
signal \N__12101\ : std_logic;
signal \N__12098\ : std_logic;
signal \N__12095\ : std_logic;
signal \N__12092\ : std_logic;
signal \N__12089\ : std_logic;
signal \N__12086\ : std_logic;
signal \N__12083\ : std_logic;
signal \N__12080\ : std_logic;
signal \N__12077\ : std_logic;
signal \N__12074\ : std_logic;
signal \N__12071\ : std_logic;
signal \N__12068\ : std_logic;
signal \N__12065\ : std_logic;
signal \N__12062\ : std_logic;
signal \N__12059\ : std_logic;
signal \N__12056\ : std_logic;
signal \N__12053\ : std_logic;
signal \N__12050\ : std_logic;
signal \N__12047\ : std_logic;
signal \N__12044\ : std_logic;
signal \N__12041\ : std_logic;
signal \N__12038\ : std_logic;
signal \N__12035\ : std_logic;
signal \N__12032\ : std_logic;
signal \N__12029\ : std_logic;
signal \N__12026\ : std_logic;
signal \N__12023\ : std_logic;
signal \N__12020\ : std_logic;
signal \N__12017\ : std_logic;
signal \N__12014\ : std_logic;
signal \N__12011\ : std_logic;
signal \N__12008\ : std_logic;
signal \N__12005\ : std_logic;
signal \N__12002\ : std_logic;
signal \N__11999\ : std_logic;
signal \N__11996\ : std_logic;
signal \N__11993\ : std_logic;
signal \N__11990\ : std_logic;
signal \N__11987\ : std_logic;
signal \N__11984\ : std_logic;
signal \N__11981\ : std_logic;
signal \N__11978\ : std_logic;
signal \N__11975\ : std_logic;
signal \N__11972\ : std_logic;
signal \N__11969\ : std_logic;
signal \N__11966\ : std_logic;
signal \N__11963\ : std_logic;
signal \N__11960\ : std_logic;
signal \N__11957\ : std_logic;
signal \N__11954\ : std_logic;
signal \N__11951\ : std_logic;
signal \N__11948\ : std_logic;
signal \N__11945\ : std_logic;
signal \N__11942\ : std_logic;
signal \N__11939\ : std_logic;
signal \N__11936\ : std_logic;
signal \N__11933\ : std_logic;
signal \N__11930\ : std_logic;
signal \N__11927\ : std_logic;
signal \N__11924\ : std_logic;
signal \N__11921\ : std_logic;
signal \N__11918\ : std_logic;
signal \N__11915\ : std_logic;
signal \N__11912\ : std_logic;
signal \N__11909\ : std_logic;
signal \N__11906\ : std_logic;
signal \N__11903\ : std_logic;
signal \N__11900\ : std_logic;
signal \N__11897\ : std_logic;
signal \N__11894\ : std_logic;
signal \N__11891\ : std_logic;
signal \N__11888\ : std_logic;
signal \N__11885\ : std_logic;
signal \N__11882\ : std_logic;
signal \N__11879\ : std_logic;
signal \N__11876\ : std_logic;
signal \N__11873\ : std_logic;
signal \N__11870\ : std_logic;
signal \N__11867\ : std_logic;
signal \N__11864\ : std_logic;
signal \N__11861\ : std_logic;
signal \N__11858\ : std_logic;
signal \N__11855\ : std_logic;
signal \N__11852\ : std_logic;
signal \N__11849\ : std_logic;
signal \N__11846\ : std_logic;
signal \N__11843\ : std_logic;
signal \N__11840\ : std_logic;
signal \N__11837\ : std_logic;
signal \N__11834\ : std_logic;
signal \N__11831\ : std_logic;
signal \N__11828\ : std_logic;
signal \N__11825\ : std_logic;
signal \N__11822\ : std_logic;
signal \N__11819\ : std_logic;
signal \N__11816\ : std_logic;
signal \N__11813\ : std_logic;
signal \N__11810\ : std_logic;
signal \N__11807\ : std_logic;
signal \N__11804\ : std_logic;
signal \N__11801\ : std_logic;
signal \N__11798\ : std_logic;
signal \N__11795\ : std_logic;
signal \N__11792\ : std_logic;
signal \N__11789\ : std_logic;
signal \N__11786\ : std_logic;
signal \N__11783\ : std_logic;
signal \N__11780\ : std_logic;
signal \N__11777\ : std_logic;
signal \N__11774\ : std_logic;
signal \N__11771\ : std_logic;
signal \N__11768\ : std_logic;
signal \N__11765\ : std_logic;
signal \N__11762\ : std_logic;
signal \N__11759\ : std_logic;
signal \N__11756\ : std_logic;
signal \N__11753\ : std_logic;
signal \N__11750\ : std_logic;
signal \N__11747\ : std_logic;
signal \N__11744\ : std_logic;
signal \N__11741\ : std_logic;
signal \N__11738\ : std_logic;
signal \N__11735\ : std_logic;
signal \N__11732\ : std_logic;
signal \N__11729\ : std_logic;
signal \N__11726\ : std_logic;
signal \N__11723\ : std_logic;
signal \N__11720\ : std_logic;
signal \N__11717\ : std_logic;
signal \N__11714\ : std_logic;
signal \N__11711\ : std_logic;
signal \N__11708\ : std_logic;
signal \N__11705\ : std_logic;
signal \N__11702\ : std_logic;
signal \N__11699\ : std_logic;
signal \N__11696\ : std_logic;
signal \N__11693\ : std_logic;
signal \N__11690\ : std_logic;
signal \N__11687\ : std_logic;
signal \N__11684\ : std_logic;
signal \N__11681\ : std_logic;
signal \N__11678\ : std_logic;
signal \N__11675\ : std_logic;
signal \N__11672\ : std_logic;
signal \N__11669\ : std_logic;
signal \N__11666\ : std_logic;
signal \N__11663\ : std_logic;
signal \N__11660\ : std_logic;
signal \N__11657\ : std_logic;
signal \N__11654\ : std_logic;
signal \N__11651\ : std_logic;
signal \N__11648\ : std_logic;
signal \N__11645\ : std_logic;
signal \N__11642\ : std_logic;
signal \N__11639\ : std_logic;
signal \N__11636\ : std_logic;
signal \N__11633\ : std_logic;
signal \N__11630\ : std_logic;
signal \N__11627\ : std_logic;
signal \N__11624\ : std_logic;
signal \N__11621\ : std_logic;
signal \N__11618\ : std_logic;
signal \N__11615\ : std_logic;
signal \N__11612\ : std_logic;
signal \N__11609\ : std_logic;
signal \N__11606\ : std_logic;
signal \N__11603\ : std_logic;
signal \N__11600\ : std_logic;
signal \N__11597\ : std_logic;
signal \N__11594\ : std_logic;
signal \N__11591\ : std_logic;
signal \N__11588\ : std_logic;
signal \N__11585\ : std_logic;
signal \N__11582\ : std_logic;
signal \N__11579\ : std_logic;
signal \N__11576\ : std_logic;
signal \N__11573\ : std_logic;
signal \N__11570\ : std_logic;
signal \N__11567\ : std_logic;
signal \N__11564\ : std_logic;
signal \N__11561\ : std_logic;
signal \N__11558\ : std_logic;
signal \N__11555\ : std_logic;
signal \N__11552\ : std_logic;
signal \N__11549\ : std_logic;
signal \N__11546\ : std_logic;
signal \N__11543\ : std_logic;
signal \N__11540\ : std_logic;
signal \N__11537\ : std_logic;
signal \N__11534\ : std_logic;
signal \N__11531\ : std_logic;
signal \N__11528\ : std_logic;
signal \N__11525\ : std_logic;
signal \N__11522\ : std_logic;
signal \N__11519\ : std_logic;
signal \N__11516\ : std_logic;
signal \N__11513\ : std_logic;
signal \N__11510\ : std_logic;
signal \N__11507\ : std_logic;
signal \N__11504\ : std_logic;
signal \N__11501\ : std_logic;
signal \N__11498\ : std_logic;
signal \N__11495\ : std_logic;
signal \N__11492\ : std_logic;
signal \N__11489\ : std_logic;
signal \N__11486\ : std_logic;
signal \N__11483\ : std_logic;
signal \N__11480\ : std_logic;
signal \N__11477\ : std_logic;
signal \N__11474\ : std_logic;
signal \N__11471\ : std_logic;
signal \N__11468\ : std_logic;
signal \N__11465\ : std_logic;
signal \N__11462\ : std_logic;
signal \N__11459\ : std_logic;
signal \N__11456\ : std_logic;
signal \N__11453\ : std_logic;
signal \N__11450\ : std_logic;
signal \N__11447\ : std_logic;
signal \N__11444\ : std_logic;
signal \N__11441\ : std_logic;
signal \N__11438\ : std_logic;
signal \N__11435\ : std_logic;
signal \N__11432\ : std_logic;
signal \N__11429\ : std_logic;
signal \N__11426\ : std_logic;
signal \N__11423\ : std_logic;
signal \N__11420\ : std_logic;
signal \N__11417\ : std_logic;
signal \N__11414\ : std_logic;
signal \N__11411\ : std_logic;
signal \N__11408\ : std_logic;
signal \N__11405\ : std_logic;
signal \N__11402\ : std_logic;
signal \N__11399\ : std_logic;
signal \N__11396\ : std_logic;
signal \N__11393\ : std_logic;
signal \N__11390\ : std_logic;
signal \N__11387\ : std_logic;
signal \N__11384\ : std_logic;
signal \N__11381\ : std_logic;
signal \N__11378\ : std_logic;
signal \N__11375\ : std_logic;
signal \N__11372\ : std_logic;
signal \N__11369\ : std_logic;
signal \N__11366\ : std_logic;
signal \N__11363\ : std_logic;
signal \N__11360\ : std_logic;
signal \N__11357\ : std_logic;
signal \N__11354\ : std_logic;
signal \N__11351\ : std_logic;
signal \N__11348\ : std_logic;
signal \N__11345\ : std_logic;
signal \N__11342\ : std_logic;
signal \N__11339\ : std_logic;
signal \N__11336\ : std_logic;
signal \N__11333\ : std_logic;
signal \N__11330\ : std_logic;
signal \N__11327\ : std_logic;
signal \N__11324\ : std_logic;
signal \N__11321\ : std_logic;
signal \N__11318\ : std_logic;
signal \N__11315\ : std_logic;
signal \N__11312\ : std_logic;
signal \N__11309\ : std_logic;
signal \N__11306\ : std_logic;
signal \N__11303\ : std_logic;
signal \N__11300\ : std_logic;
signal \N__11297\ : std_logic;
signal \N__11294\ : std_logic;
signal \N__11291\ : std_logic;
signal \N__11288\ : std_logic;
signal \N__11285\ : std_logic;
signal \N__11282\ : std_logic;
signal \N__11279\ : std_logic;
signal \N__11276\ : std_logic;
signal \N__11273\ : std_logic;
signal \N__11270\ : std_logic;
signal \N__11267\ : std_logic;
signal \N__11264\ : std_logic;
signal \N__11261\ : std_logic;
signal \N__11258\ : std_logic;
signal \N__11255\ : std_logic;
signal \N__11252\ : std_logic;
signal \N__11249\ : std_logic;
signal \N__11246\ : std_logic;
signal \N__11243\ : std_logic;
signal \N__11240\ : std_logic;
signal \N__11237\ : std_logic;
signal \N__11234\ : std_logic;
signal \N__11231\ : std_logic;
signal \N__11228\ : std_logic;
signal \N__11225\ : std_logic;
signal \N__11222\ : std_logic;
signal \N__11219\ : std_logic;
signal \N__11216\ : std_logic;
signal \N__11213\ : std_logic;
signal \N__11210\ : std_logic;
signal \N__11207\ : std_logic;
signal \N__11204\ : std_logic;
signal \N__11201\ : std_logic;
signal \N__11198\ : std_logic;
signal \N__11195\ : std_logic;
signal \N__11192\ : std_logic;
signal \N__11189\ : std_logic;
signal \N__11186\ : std_logic;
signal \N__11183\ : std_logic;
signal \N__11180\ : std_logic;
signal \N__11177\ : std_logic;
signal \N__11174\ : std_logic;
signal \N__11171\ : std_logic;
signal \N__11168\ : std_logic;
signal \N__11165\ : std_logic;
signal \N__11162\ : std_logic;
signal \N__11159\ : std_logic;
signal \N__11156\ : std_logic;
signal \N__11153\ : std_logic;
signal \N__11150\ : std_logic;
signal \N__11147\ : std_logic;
signal \N__11144\ : std_logic;
signal \N__11141\ : std_logic;
signal \N__11138\ : std_logic;
signal \N__11135\ : std_logic;
signal \N__11132\ : std_logic;
signal \N__11129\ : std_logic;
signal \N__11126\ : std_logic;
signal \N__11123\ : std_logic;
signal \N__11120\ : std_logic;
signal \N__11117\ : std_logic;
signal \N__11114\ : std_logic;
signal \N__11111\ : std_logic;
signal \N__11108\ : std_logic;
signal \N__11105\ : std_logic;
signal \N__11102\ : std_logic;
signal \N__11099\ : std_logic;
signal \N__11096\ : std_logic;
signal \N__11093\ : std_logic;
signal \N__11090\ : std_logic;
signal \N__11087\ : std_logic;
signal \N__11084\ : std_logic;
signal \N__11081\ : std_logic;
signal \N__11078\ : std_logic;
signal \N__11075\ : std_logic;
signal \N__11072\ : std_logic;
signal \N__11069\ : std_logic;
signal \N__11066\ : std_logic;
signal \N__11063\ : std_logic;
signal \N__11060\ : std_logic;
signal \N__11057\ : std_logic;
signal \N__11054\ : std_logic;
signal \N__11051\ : std_logic;
signal \N__11048\ : std_logic;
signal \N__11045\ : std_logic;
signal \N__11042\ : std_logic;
signal \N__11039\ : std_logic;
signal \N__11036\ : std_logic;
signal \N__11033\ : std_logic;
signal \N__11030\ : std_logic;
signal \N__11027\ : std_logic;
signal \N__11024\ : std_logic;
signal \N__11021\ : std_logic;
signal \N__11018\ : std_logic;
signal \N__11015\ : std_logic;
signal \N__11012\ : std_logic;
signal \N__11009\ : std_logic;
signal \N__11006\ : std_logic;
signal \N__11003\ : std_logic;
signal \N__11000\ : std_logic;
signal \N__10999\ : std_logic;
signal \N__10998\ : std_logic;
signal \N__10995\ : std_logic;
signal \N__10992\ : std_logic;
signal \N__10991\ : std_logic;
signal \N__10990\ : std_logic;
signal \N__10987\ : std_logic;
signal \N__10986\ : std_logic;
signal \N__10985\ : std_logic;
signal \N__10980\ : std_logic;
signal \N__10977\ : std_logic;
signal \N__10974\ : std_logic;
signal \N__10971\ : std_logic;
signal \N__10968\ : std_logic;
signal \N__10965\ : std_logic;
signal \N__10964\ : std_logic;
signal \N__10963\ : std_logic;
signal \N__10962\ : std_logic;
signal \N__10961\ : std_logic;
signal \N__10960\ : std_logic;
signal \N__10953\ : std_logic;
signal \N__10946\ : std_logic;
signal \N__10943\ : std_logic;
signal \N__10940\ : std_logic;
signal \N__10937\ : std_logic;
signal \N__10934\ : std_logic;
signal \N__10933\ : std_logic;
signal \N__10932\ : std_logic;
signal \N__10931\ : std_logic;
signal \N__10928\ : std_logic;
signal \N__10927\ : std_logic;
signal \N__10926\ : std_logic;
signal \N__10925\ : std_logic;
signal \N__10924\ : std_logic;
signal \N__10923\ : std_logic;
signal \N__10922\ : std_logic;
signal \N__10921\ : std_logic;
signal \N__10920\ : std_logic;
signal \N__10911\ : std_logic;
signal \N__10906\ : std_logic;
signal \N__10903\ : std_logic;
signal \N__10900\ : std_logic;
signal \N__10899\ : std_logic;
signal \N__10898\ : std_logic;
signal \N__10895\ : std_logic;
signal \N__10892\ : std_logic;
signal \N__10889\ : std_logic;
signal \N__10886\ : std_logic;
signal \N__10885\ : std_logic;
signal \N__10882\ : std_logic;
signal \N__10879\ : std_logic;
signal \N__10878\ : std_logic;
signal \N__10877\ : std_logic;
signal \N__10876\ : std_logic;
signal \N__10873\ : std_logic;
signal \N__10870\ : std_logic;
signal \N__10869\ : std_logic;
signal \N__10868\ : std_logic;
signal \N__10865\ : std_logic;
signal \N__10864\ : std_logic;
signal \N__10863\ : std_logic;
signal \N__10862\ : std_logic;
signal \N__10859\ : std_logic;
signal \N__10858\ : std_logic;
signal \N__10849\ : std_logic;
signal \N__10846\ : std_logic;
signal \N__10843\ : std_logic;
signal \N__10842\ : std_logic;
signal \N__10835\ : std_logic;
signal \N__10832\ : std_logic;
signal \N__10829\ : std_logic;
signal \N__10828\ : std_logic;
signal \N__10823\ : std_logic;
signal \N__10820\ : std_logic;
signal \N__10817\ : std_logic;
signal \N__10816\ : std_logic;
signal \N__10813\ : std_logic;
signal \N__10812\ : std_logic;
signal \N__10811\ : std_logic;
signal \N__10808\ : std_logic;
signal \N__10805\ : std_logic;
signal \N__10802\ : std_logic;
signal \N__10799\ : std_logic;
signal \N__10798\ : std_logic;
signal \N__10795\ : std_logic;
signal \N__10792\ : std_logic;
signal \N__10789\ : std_logic;
signal \N__10788\ : std_logic;
signal \N__10787\ : std_logic;
signal \N__10786\ : std_logic;
signal \N__10783\ : std_logic;
signal \N__10780\ : std_logic;
signal \N__10777\ : std_logic;
signal \N__10770\ : std_logic;
signal \N__10767\ : std_logic;
signal \N__10760\ : std_logic;
signal \N__10757\ : std_logic;
signal \N__10750\ : std_logic;
signal \N__10747\ : std_logic;
signal \N__10744\ : std_logic;
signal \N__10741\ : std_logic;
signal \N__10740\ : std_logic;
signal \N__10737\ : std_logic;
signal \N__10736\ : std_logic;
signal \N__10727\ : std_logic;
signal \N__10724\ : std_logic;
signal \N__10717\ : std_logic;
signal \N__10714\ : std_logic;
signal \N__10711\ : std_logic;
signal \N__10710\ : std_logic;
signal \N__10709\ : std_logic;
signal \N__10706\ : std_logic;
signal \N__10705\ : std_logic;
signal \N__10704\ : std_logic;
signal \N__10703\ : std_logic;
signal \N__10696\ : std_logic;
signal \N__10687\ : std_logic;
signal \N__10678\ : std_logic;
signal \N__10675\ : std_logic;
signal \N__10672\ : std_logic;
signal \N__10669\ : std_logic;
signal \N__10664\ : std_logic;
signal \N__10657\ : std_logic;
signal \N__10654\ : std_logic;
signal \N__10651\ : std_logic;
signal \N__10648\ : std_logic;
signal \N__10645\ : std_logic;
signal \N__10642\ : std_logic;
signal \N__10641\ : std_logic;
signal \N__10640\ : std_logic;
signal \N__10639\ : std_logic;
signal \N__10638\ : std_logic;
signal \N__10637\ : std_logic;
signal \N__10636\ : std_logic;
signal \N__10633\ : std_logic;
signal \N__10632\ : std_logic;
signal \N__10631\ : std_logic;
signal \N__10624\ : std_logic;
signal \N__10617\ : std_logic;
signal \N__10608\ : std_logic;
signal \N__10601\ : std_logic;
signal \N__10598\ : std_logic;
signal \N__10595\ : std_logic;
signal \N__10594\ : std_logic;
signal \N__10591\ : std_logic;
signal \N__10590\ : std_logic;
signal \N__10589\ : std_logic;
signal \N__10586\ : std_logic;
signal \N__10583\ : std_logic;
signal \N__10582\ : std_logic;
signal \N__10579\ : std_logic;
signal \N__10576\ : std_logic;
signal \N__10573\ : std_logic;
signal \N__10570\ : std_logic;
signal \N__10567\ : std_logic;
signal \N__10564\ : std_logic;
signal \N__10555\ : std_logic;
signal \N__10552\ : std_logic;
signal \N__10549\ : std_logic;
signal \N__10546\ : std_logic;
signal \N__10543\ : std_logic;
signal \N__10540\ : std_logic;
signal \N__10537\ : std_logic;
signal \N__10534\ : std_logic;
signal \N__10531\ : std_logic;
signal \N__10530\ : std_logic;
signal \N__10527\ : std_logic;
signal \N__10524\ : std_logic;
signal \N__10521\ : std_logic;
signal \N__10518\ : std_logic;
signal \N__10513\ : std_logic;
signal \N__10510\ : std_logic;
signal \N__10507\ : std_logic;
signal \N__10504\ : std_logic;
signal \N__10501\ : std_logic;
signal \N__10496\ : std_logic;
signal \N__10493\ : std_logic;
signal \N__10490\ : std_logic;
signal \N__10487\ : std_logic;
signal \N__10480\ : std_logic;
signal \N__10475\ : std_logic;
signal \N__10472\ : std_logic;
signal \N__10465\ : std_logic;
signal \N__10460\ : std_logic;
signal \N__10455\ : std_logic;
signal \N__10452\ : std_logic;
signal \N__10439\ : std_logic;
signal \N__10436\ : std_logic;
signal \N__10433\ : std_logic;
signal \N__10430\ : std_logic;
signal \N__10427\ : std_logic;
signal \N__10424\ : std_logic;
signal \N__10421\ : std_logic;
signal \N__10418\ : std_logic;
signal \N__10415\ : std_logic;
signal \N__10412\ : std_logic;
signal \N__10409\ : std_logic;
signal \N__10406\ : std_logic;
signal \N__10403\ : std_logic;
signal \N__10400\ : std_logic;
signal \N__10397\ : std_logic;
signal \N__10394\ : std_logic;
signal \N__10391\ : std_logic;
signal \N__10388\ : std_logic;
signal \N__10385\ : std_logic;
signal \N__10382\ : std_logic;
signal \N__10379\ : std_logic;
signal \N__10376\ : std_logic;
signal \N__10373\ : std_logic;
signal \N__10370\ : std_logic;
signal \N__10367\ : std_logic;
signal \N__10364\ : std_logic;
signal \N__10361\ : std_logic;
signal \N__10358\ : std_logic;
signal \N__10355\ : std_logic;
signal \N__10352\ : std_logic;
signal \N__10349\ : std_logic;
signal \N__10346\ : std_logic;
signal \N__10343\ : std_logic;
signal \N__10340\ : std_logic;
signal \N__10337\ : std_logic;
signal \N__10334\ : std_logic;
signal \N__10331\ : std_logic;
signal \N__10328\ : std_logic;
signal \N__10325\ : std_logic;
signal \N__10324\ : std_logic;
signal \N__10321\ : std_logic;
signal \N__10318\ : std_logic;
signal \N__10317\ : std_logic;
signal \N__10314\ : std_logic;
signal \N__10311\ : std_logic;
signal \N__10308\ : std_logic;
signal \N__10301\ : std_logic;
signal \N__10300\ : std_logic;
signal \N__10297\ : std_logic;
signal \N__10294\ : std_logic;
signal \N__10289\ : std_logic;
signal \N__10288\ : std_logic;
signal \N__10285\ : std_logic;
signal \N__10282\ : std_logic;
signal \N__10281\ : std_logic;
signal \N__10276\ : std_logic;
signal \N__10273\ : std_logic;
signal \N__10272\ : std_logic;
signal \N__10267\ : std_logic;
signal \N__10264\ : std_logic;
signal \N__10261\ : std_logic;
signal \N__10258\ : std_logic;
signal \N__10255\ : std_logic;
signal \N__10252\ : std_logic;
signal \N__10247\ : std_logic;
signal \N__10246\ : std_logic;
signal \N__10243\ : std_logic;
signal \N__10240\ : std_logic;
signal \N__10239\ : std_logic;
signal \N__10238\ : std_logic;
signal \N__10233\ : std_logic;
signal \N__10230\ : std_logic;
signal \N__10227\ : std_logic;
signal \N__10220\ : std_logic;
signal \N__10217\ : std_logic;
signal \N__10214\ : std_logic;
signal \N__10211\ : std_logic;
signal \N__10208\ : std_logic;
signal \N__10205\ : std_logic;
signal \N__10202\ : std_logic;
signal \N__10199\ : std_logic;
signal \N__10198\ : std_logic;
signal \N__10197\ : std_logic;
signal \N__10196\ : std_logic;
signal \N__10193\ : std_logic;
signal \N__10190\ : std_logic;
signal \N__10187\ : std_logic;
signal \N__10184\ : std_logic;
signal \N__10181\ : std_logic;
signal \N__10178\ : std_logic;
signal \N__10173\ : std_logic;
signal \N__10168\ : std_logic;
signal \N__10165\ : std_logic;
signal \N__10162\ : std_logic;
signal \N__10159\ : std_logic;
signal \N__10156\ : std_logic;
signal \N__10153\ : std_logic;
signal \N__10148\ : std_logic;
signal \N__10145\ : std_logic;
signal \N__10144\ : std_logic;
signal \N__10141\ : std_logic;
signal \N__10138\ : std_logic;
signal \N__10137\ : std_logic;
signal \N__10136\ : std_logic;
signal \N__10131\ : std_logic;
signal \N__10128\ : std_logic;
signal \N__10125\ : std_logic;
signal \N__10118\ : std_logic;
signal \N__10115\ : std_logic;
signal \N__10112\ : std_logic;
signal \N__10109\ : std_logic;
signal \N__10106\ : std_logic;
signal \N__10103\ : std_logic;
signal \N__10100\ : std_logic;
signal \N__10099\ : std_logic;
signal \N__10098\ : std_logic;
signal \N__10097\ : std_logic;
signal \N__10096\ : std_logic;
signal \N__10095\ : std_logic;
signal \N__10094\ : std_logic;
signal \N__10093\ : std_logic;
signal \N__10076\ : std_logic;
signal \N__10073\ : std_logic;
signal \N__10070\ : std_logic;
signal \N__10067\ : std_logic;
signal \N__10064\ : std_logic;
signal \N__10063\ : std_logic;
signal \N__10062\ : std_logic;
signal \N__10061\ : std_logic;
signal \N__10060\ : std_logic;
signal \N__10059\ : std_logic;
signal \N__10058\ : std_logic;
signal \N__10057\ : std_logic;
signal \N__10040\ : std_logic;
signal \N__10037\ : std_logic;
signal \N__10034\ : std_logic;
signal \N__10031\ : std_logic;
signal \N__10028\ : std_logic;
signal \N__10027\ : std_logic;
signal \N__10026\ : std_logic;
signal \N__10025\ : std_logic;
signal \N__10022\ : std_logic;
signal \N__10021\ : std_logic;
signal \N__10018\ : std_logic;
signal \N__10017\ : std_logic;
signal \N__10014\ : std_logic;
signal \N__10013\ : std_logic;
signal \N__10010\ : std_logic;
signal \N__10009\ : std_logic;
signal \N__9992\ : std_logic;
signal \N__9989\ : std_logic;
signal \N__9986\ : std_logic;
signal \N__9983\ : std_logic;
signal \N__9980\ : std_logic;
signal \N__9979\ : std_logic;
signal \N__9978\ : std_logic;
signal \N__9977\ : std_logic;
signal \N__9976\ : std_logic;
signal \N__9973\ : std_logic;
signal \N__9972\ : std_logic;
signal \N__9969\ : std_logic;
signal \N__9968\ : std_logic;
signal \N__9965\ : std_logic;
signal \N__9964\ : std_logic;
signal \N__9961\ : std_logic;
signal \N__9944\ : std_logic;
signal \N__9941\ : std_logic;
signal \N__9938\ : std_logic;
signal \N__9937\ : std_logic;
signal \N__9936\ : std_logic;
signal \N__9935\ : std_logic;
signal \N__9932\ : std_logic;
signal \N__9929\ : std_logic;
signal \N__9926\ : std_logic;
signal \N__9923\ : std_logic;
signal \N__9918\ : std_logic;
signal \N__9913\ : std_logic;
signal \N__9908\ : std_logic;
signal \N__9905\ : std_logic;
signal \N__9902\ : std_logic;
signal \N__9899\ : std_logic;
signal \N__9896\ : std_logic;
signal \N__9893\ : std_logic;
signal \N__9890\ : std_logic;
signal \N__9887\ : std_logic;
signal \N__9884\ : std_logic;
signal \N__9881\ : std_logic;
signal \N__9878\ : std_logic;
signal \N__9875\ : std_logic;
signal \N__9872\ : std_logic;
signal \N__9869\ : std_logic;
signal \N__9866\ : std_logic;
signal \N__9863\ : std_logic;
signal \N__9860\ : std_logic;
signal \N__9857\ : std_logic;
signal \N__9854\ : std_logic;
signal \N__9851\ : std_logic;
signal \N__9848\ : std_logic;
signal \N__9845\ : std_logic;
signal \N__9842\ : std_logic;
signal \N__9839\ : std_logic;
signal \N__9836\ : std_logic;
signal \N__9833\ : std_logic;
signal \N__9830\ : std_logic;
signal \N__9827\ : std_logic;
signal \N__9824\ : std_logic;
signal \N__9821\ : std_logic;
signal \N__9818\ : std_logic;
signal \N__9815\ : std_logic;
signal \N__9814\ : std_logic;
signal \N__9811\ : std_logic;
signal \N__9808\ : std_logic;
signal \N__9805\ : std_logic;
signal \N__9802\ : std_logic;
signal \N__9799\ : std_logic;
signal \N__9796\ : std_logic;
signal \N__9793\ : std_logic;
signal \N__9790\ : std_logic;
signal \N__9787\ : std_logic;
signal \N__9784\ : std_logic;
signal \N__9781\ : std_logic;
signal \N__9778\ : std_logic;
signal \N__9775\ : std_logic;
signal \N__9772\ : std_logic;
signal \N__9769\ : std_logic;
signal \N__9766\ : std_logic;
signal \N__9763\ : std_logic;
signal \N__9760\ : std_logic;
signal \N__9757\ : std_logic;
signal \N__9754\ : std_logic;
signal \N__9751\ : std_logic;
signal \N__9748\ : std_logic;
signal \N__9745\ : std_logic;
signal \N__9742\ : std_logic;
signal \N__9739\ : std_logic;
signal \N__9736\ : std_logic;
signal \N__9733\ : std_logic;
signal \N__9730\ : std_logic;
signal \N__9727\ : std_logic;
signal \N__9724\ : std_logic;
signal \N__9721\ : std_logic;
signal \N__9718\ : std_logic;
signal \N__9715\ : std_logic;
signal \N__9712\ : std_logic;
signal \N__9709\ : std_logic;
signal \N__9706\ : std_logic;
signal \N__9703\ : std_logic;
signal \N__9700\ : std_logic;
signal \N__9697\ : std_logic;
signal \N__9694\ : std_logic;
signal \N__9691\ : std_logic;
signal \N__9688\ : std_logic;
signal \N__9685\ : std_logic;
signal \N__9682\ : std_logic;
signal \N__9679\ : std_logic;
signal \N__9676\ : std_logic;
signal \N__9673\ : std_logic;
signal \N__9670\ : std_logic;
signal \N__9667\ : std_logic;
signal \N__9664\ : std_logic;
signal \N__9661\ : std_logic;
signal \N__9658\ : std_logic;
signal \N__9655\ : std_logic;
signal \N__9652\ : std_logic;
signal \N__9649\ : std_logic;
signal \N__9646\ : std_logic;
signal \N__9643\ : std_logic;
signal \N__9640\ : std_logic;
signal \N__9637\ : std_logic;
signal \N__9634\ : std_logic;
signal \N__9631\ : std_logic;
signal \N__9628\ : std_logic;
signal \N__9625\ : std_logic;
signal \N__9622\ : std_logic;
signal \N__9619\ : std_logic;
signal \N__9616\ : std_logic;
signal \N__9613\ : std_logic;
signal \N__9610\ : std_logic;
signal \N__9605\ : std_logic;
signal \N__9602\ : std_logic;
signal \N__9599\ : std_logic;
signal \N__9598\ : std_logic;
signal \N__9597\ : std_logic;
signal \N__9594\ : std_logic;
signal \N__9591\ : std_logic;
signal \N__9588\ : std_logic;
signal \N__9587\ : std_logic;
signal \N__9580\ : std_logic;
signal \N__9577\ : std_logic;
signal \N__9572\ : std_logic;
signal \N__9569\ : std_logic;
signal \N__9566\ : std_logic;
signal \N__9565\ : std_logic;
signal \N__9562\ : std_logic;
signal \N__9559\ : std_logic;
signal \N__9558\ : std_logic;
signal \N__9555\ : std_logic;
signal \N__9552\ : std_logic;
signal \N__9549\ : std_logic;
signal \N__9542\ : std_logic;
signal \N__9541\ : std_logic;
signal \N__9538\ : std_logic;
signal \N__9535\ : std_logic;
signal \N__9530\ : std_logic;
signal \N__9527\ : std_logic;
signal \N__9524\ : std_logic;
signal \N__9523\ : std_logic;
signal \N__9522\ : std_logic;
signal \N__9521\ : std_logic;
signal \N__9520\ : std_logic;
signal \N__9517\ : std_logic;
signal \N__9516\ : std_logic;
signal \N__9513\ : std_logic;
signal \N__9510\ : std_logic;
signal \N__9507\ : std_logic;
signal \N__9504\ : std_logic;
signal \N__9501\ : std_logic;
signal \N__9498\ : std_logic;
signal \N__9497\ : std_logic;
signal \N__9494\ : std_logic;
signal \N__9491\ : std_logic;
signal \N__9488\ : std_logic;
signal \N__9487\ : std_logic;
signal \N__9484\ : std_logic;
signal \N__9479\ : std_logic;
signal \N__9476\ : std_logic;
signal \N__9473\ : std_logic;
signal \N__9468\ : std_logic;
signal \N__9465\ : std_logic;
signal \N__9462\ : std_logic;
signal \N__9459\ : std_logic;
signal \N__9456\ : std_logic;
signal \N__9453\ : std_logic;
signal \N__9450\ : std_logic;
signal \N__9447\ : std_logic;
signal \N__9442\ : std_logic;
signal \N__9439\ : std_logic;
signal \N__9436\ : std_logic;
signal \N__9431\ : std_logic;
signal \N__9422\ : std_logic;
signal \N__9419\ : std_logic;
signal \N__9416\ : std_logic;
signal \N__9413\ : std_logic;
signal \N__9412\ : std_logic;
signal \N__9409\ : std_logic;
signal \N__9406\ : std_logic;
signal \N__9403\ : std_logic;
signal \N__9400\ : std_logic;
signal \N__9397\ : std_logic;
signal \N__9394\ : std_logic;
signal \N__9391\ : std_logic;
signal \N__9388\ : std_logic;
signal \N__9385\ : std_logic;
signal \N__9382\ : std_logic;
signal \N__9379\ : std_logic;
signal \N__9376\ : std_logic;
signal \N__9373\ : std_logic;
signal \N__9370\ : std_logic;
signal \N__9367\ : std_logic;
signal \N__9364\ : std_logic;
signal \N__9361\ : std_logic;
signal \N__9358\ : std_logic;
signal \N__9355\ : std_logic;
signal \N__9352\ : std_logic;
signal \N__9349\ : std_logic;
signal \N__9346\ : std_logic;
signal \N__9343\ : std_logic;
signal \N__9340\ : std_logic;
signal \N__9337\ : std_logic;
signal \N__9334\ : std_logic;
signal \N__9331\ : std_logic;
signal \N__9328\ : std_logic;
signal \N__9325\ : std_logic;
signal \N__9322\ : std_logic;
signal \N__9319\ : std_logic;
signal \N__9316\ : std_logic;
signal \N__9313\ : std_logic;
signal \N__9310\ : std_logic;
signal \N__9307\ : std_logic;
signal \N__9304\ : std_logic;
signal \N__9301\ : std_logic;
signal \N__9298\ : std_logic;
signal \N__9295\ : std_logic;
signal \N__9292\ : std_logic;
signal \N__9289\ : std_logic;
signal \N__9286\ : std_logic;
signal \N__9283\ : std_logic;
signal \N__9280\ : std_logic;
signal \N__9277\ : std_logic;
signal \N__9274\ : std_logic;
signal \N__9271\ : std_logic;
signal \N__9268\ : std_logic;
signal \N__9265\ : std_logic;
signal \N__9262\ : std_logic;
signal \N__9259\ : std_logic;
signal \N__9256\ : std_logic;
signal \N__9253\ : std_logic;
signal \N__9250\ : std_logic;
signal \N__9247\ : std_logic;
signal \N__9244\ : std_logic;
signal \N__9241\ : std_logic;
signal \N__9238\ : std_logic;
signal \N__9235\ : std_logic;
signal \N__9232\ : std_logic;
signal \N__9229\ : std_logic;
signal \N__9226\ : std_logic;
signal \N__9223\ : std_logic;
signal \N__9220\ : std_logic;
signal \N__9217\ : std_logic;
signal \N__9214\ : std_logic;
signal \N__9211\ : std_logic;
signal \N__9208\ : std_logic;
signal \N__9203\ : std_logic;
signal \N__9200\ : std_logic;
signal \N__9197\ : std_logic;
signal \N__9194\ : std_logic;
signal \N__9193\ : std_logic;
signal \N__9190\ : std_logic;
signal \N__9187\ : std_logic;
signal \N__9184\ : std_logic;
signal \N__9181\ : std_logic;
signal \N__9178\ : std_logic;
signal \N__9175\ : std_logic;
signal \N__9172\ : std_logic;
signal \N__9169\ : std_logic;
signal \N__9166\ : std_logic;
signal \N__9163\ : std_logic;
signal \N__9160\ : std_logic;
signal \N__9157\ : std_logic;
signal \N__9154\ : std_logic;
signal \N__9151\ : std_logic;
signal \N__9148\ : std_logic;
signal \N__9145\ : std_logic;
signal \N__9142\ : std_logic;
signal \N__9139\ : std_logic;
signal \N__9136\ : std_logic;
signal \N__9133\ : std_logic;
signal \N__9130\ : std_logic;
signal \N__9127\ : std_logic;
signal \N__9124\ : std_logic;
signal \N__9121\ : std_logic;
signal \N__9118\ : std_logic;
signal \N__9115\ : std_logic;
signal \N__9112\ : std_logic;
signal \N__9109\ : std_logic;
signal \N__9106\ : std_logic;
signal \N__9103\ : std_logic;
signal \N__9100\ : std_logic;
signal \N__9097\ : std_logic;
signal \N__9094\ : std_logic;
signal \N__9091\ : std_logic;
signal \N__9088\ : std_logic;
signal \N__9085\ : std_logic;
signal \N__9082\ : std_logic;
signal \N__9079\ : std_logic;
signal \N__9076\ : std_logic;
signal \N__9073\ : std_logic;
signal \N__9070\ : std_logic;
signal \N__9067\ : std_logic;
signal \N__9064\ : std_logic;
signal \N__9061\ : std_logic;
signal \N__9058\ : std_logic;
signal \N__9055\ : std_logic;
signal \N__9052\ : std_logic;
signal \N__9049\ : std_logic;
signal \N__9046\ : std_logic;
signal \N__9043\ : std_logic;
signal \N__9040\ : std_logic;
signal \N__9037\ : std_logic;
signal \N__9034\ : std_logic;
signal \N__9031\ : std_logic;
signal \N__9028\ : std_logic;
signal \N__9025\ : std_logic;
signal \N__9022\ : std_logic;
signal \N__9019\ : std_logic;
signal \N__9016\ : std_logic;
signal \N__9013\ : std_logic;
signal \N__9010\ : std_logic;
signal \N__9007\ : std_logic;
signal \N__9004\ : std_logic;
signal \N__9001\ : std_logic;
signal \N__8998\ : std_logic;
signal \N__8995\ : std_logic;
signal \N__8992\ : std_logic;
signal \N__8989\ : std_logic;
signal \N__8984\ : std_logic;
signal \N__8981\ : std_logic;
signal \N__8978\ : std_logic;
signal \N__8975\ : std_logic;
signal \N__8972\ : std_logic;
signal \N__8969\ : std_logic;
signal \N__8968\ : std_logic;
signal \N__8965\ : std_logic;
signal \N__8962\ : std_logic;
signal \N__8959\ : std_logic;
signal \N__8956\ : std_logic;
signal \N__8953\ : std_logic;
signal \N__8950\ : std_logic;
signal \N__8947\ : std_logic;
signal \N__8944\ : std_logic;
signal \N__8941\ : std_logic;
signal \N__8938\ : std_logic;
signal \N__8935\ : std_logic;
signal \N__8932\ : std_logic;
signal \N__8929\ : std_logic;
signal \N__8926\ : std_logic;
signal \N__8923\ : std_logic;
signal \N__8920\ : std_logic;
signal \N__8917\ : std_logic;
signal \N__8914\ : std_logic;
signal \N__8911\ : std_logic;
signal \N__8908\ : std_logic;
signal \N__8905\ : std_logic;
signal \N__8902\ : std_logic;
signal \N__8899\ : std_logic;
signal \N__8896\ : std_logic;
signal \N__8893\ : std_logic;
signal \N__8890\ : std_logic;
signal \N__8887\ : std_logic;
signal \N__8884\ : std_logic;
signal \N__8881\ : std_logic;
signal \N__8878\ : std_logic;
signal \N__8875\ : std_logic;
signal \N__8872\ : std_logic;
signal \N__8869\ : std_logic;
signal \N__8866\ : std_logic;
signal \N__8863\ : std_logic;
signal \N__8860\ : std_logic;
signal \N__8857\ : std_logic;
signal \N__8854\ : std_logic;
signal \N__8851\ : std_logic;
signal \N__8848\ : std_logic;
signal \N__8845\ : std_logic;
signal \N__8842\ : std_logic;
signal \N__8839\ : std_logic;
signal \N__8836\ : std_logic;
signal \N__8833\ : std_logic;
signal \N__8830\ : std_logic;
signal \N__8827\ : std_logic;
signal \N__8824\ : std_logic;
signal \N__8821\ : std_logic;
signal \N__8818\ : std_logic;
signal \N__8815\ : std_logic;
signal \N__8812\ : std_logic;
signal \N__8809\ : std_logic;
signal \N__8806\ : std_logic;
signal \N__8803\ : std_logic;
signal \N__8800\ : std_logic;
signal \N__8797\ : std_logic;
signal \N__8794\ : std_logic;
signal \N__8791\ : std_logic;
signal \N__8788\ : std_logic;
signal \N__8785\ : std_logic;
signal \N__8782\ : std_logic;
signal \N__8779\ : std_logic;
signal \N__8776\ : std_logic;
signal \N__8771\ : std_logic;
signal \N__8770\ : std_logic;
signal \N__8769\ : std_logic;
signal \N__8768\ : std_logic;
signal \N__8767\ : std_logic;
signal \N__8766\ : std_logic;
signal \N__8765\ : std_logic;
signal \N__8764\ : std_logic;
signal \N__8763\ : std_logic;
signal \N__8762\ : std_logic;
signal \N__8761\ : std_logic;
signal \N__8760\ : std_logic;
signal \N__8759\ : std_logic;
signal \N__8758\ : std_logic;
signal \N__8757\ : std_logic;
signal \N__8756\ : std_logic;
signal \N__8755\ : std_logic;
signal \N__8754\ : std_logic;
signal \N__8753\ : std_logic;
signal \N__8752\ : std_logic;
signal \N__8751\ : std_logic;
signal \N__8750\ : std_logic;
signal \N__8749\ : std_logic;
signal \N__8748\ : std_logic;
signal \N__8747\ : std_logic;
signal \N__8746\ : std_logic;
signal \N__8745\ : std_logic;
signal \N__8744\ : std_logic;
signal \N__8743\ : std_logic;
signal \N__8742\ : std_logic;
signal \N__8741\ : std_logic;
signal \N__8740\ : std_logic;
signal \N__8675\ : std_logic;
signal \N__8672\ : std_logic;
signal \N__8669\ : std_logic;
signal \N__8666\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8662\ : std_logic;
signal \N__8659\ : std_logic;
signal \N__8656\ : std_logic;
signal \N__8653\ : std_logic;
signal \N__8650\ : std_logic;
signal \N__8647\ : std_logic;
signal \N__8644\ : std_logic;
signal \N__8641\ : std_logic;
signal \N__8638\ : std_logic;
signal \N__8635\ : std_logic;
signal \N__8632\ : std_logic;
signal \N__8629\ : std_logic;
signal \N__8626\ : std_logic;
signal \N__8623\ : std_logic;
signal \N__8620\ : std_logic;
signal \N__8617\ : std_logic;
signal \N__8614\ : std_logic;
signal \N__8611\ : std_logic;
signal \N__8608\ : std_logic;
signal \N__8605\ : std_logic;
signal \N__8602\ : std_logic;
signal \N__8599\ : std_logic;
signal \N__8596\ : std_logic;
signal \N__8593\ : std_logic;
signal \N__8590\ : std_logic;
signal \N__8587\ : std_logic;
signal \N__8584\ : std_logic;
signal \N__8581\ : std_logic;
signal \N__8578\ : std_logic;
signal \N__8575\ : std_logic;
signal \N__8572\ : std_logic;
signal \N__8569\ : std_logic;
signal \N__8566\ : std_logic;
signal \N__8563\ : std_logic;
signal \N__8560\ : std_logic;
signal \N__8557\ : std_logic;
signal \N__8554\ : std_logic;
signal \N__8551\ : std_logic;
signal \N__8548\ : std_logic;
signal \N__8545\ : std_logic;
signal \N__8542\ : std_logic;
signal \N__8539\ : std_logic;
signal \N__8536\ : std_logic;
signal \N__8533\ : std_logic;
signal \N__8530\ : std_logic;
signal \N__8527\ : std_logic;
signal \N__8524\ : std_logic;
signal \N__8521\ : std_logic;
signal \N__8518\ : std_logic;
signal \N__8515\ : std_logic;
signal \N__8512\ : std_logic;
signal \N__8509\ : std_logic;
signal \N__8506\ : std_logic;
signal \N__8503\ : std_logic;
signal \N__8500\ : std_logic;
signal \N__8497\ : std_logic;
signal \N__8494\ : std_logic;
signal \N__8491\ : std_logic;
signal \N__8488\ : std_logic;
signal \N__8485\ : std_logic;
signal \N__8482\ : std_logic;
signal \N__8479\ : std_logic;
signal \N__8476\ : std_logic;
signal \N__8473\ : std_logic;
signal \N__8470\ : std_logic;
signal \N__8467\ : std_logic;
signal \N__8464\ : std_logic;
signal \N__8461\ : std_logic;
signal \N__8458\ : std_logic;
signal \N__8455\ : std_logic;
signal \N__8452\ : std_logic;
signal \N__8447\ : std_logic;
signal \N__8444\ : std_logic;
signal \N__8441\ : std_logic;
signal \N__8438\ : std_logic;
signal \N__8437\ : std_logic;
signal \N__8434\ : std_logic;
signal \N__8431\ : std_logic;
signal \N__8428\ : std_logic;
signal \N__8425\ : std_logic;
signal \N__8422\ : std_logic;
signal \N__8419\ : std_logic;
signal \N__8416\ : std_logic;
signal \N__8413\ : std_logic;
signal \N__8410\ : std_logic;
signal \N__8407\ : std_logic;
signal \N__8404\ : std_logic;
signal \N__8401\ : std_logic;
signal \N__8398\ : std_logic;
signal \N__8395\ : std_logic;
signal \N__8392\ : std_logic;
signal \N__8389\ : std_logic;
signal \N__8386\ : std_logic;
signal \N__8383\ : std_logic;
signal \N__8380\ : std_logic;
signal \N__8377\ : std_logic;
signal \N__8374\ : std_logic;
signal \N__8371\ : std_logic;
signal \N__8368\ : std_logic;
signal \N__8365\ : std_logic;
signal \N__8362\ : std_logic;
signal \N__8359\ : std_logic;
signal \N__8356\ : std_logic;
signal \N__8353\ : std_logic;
signal \N__8350\ : std_logic;
signal \N__8347\ : std_logic;
signal \N__8344\ : std_logic;
signal \N__8341\ : std_logic;
signal \N__8338\ : std_logic;
signal \N__8335\ : std_logic;
signal \N__8332\ : std_logic;
signal \N__8329\ : std_logic;
signal \N__8326\ : std_logic;
signal \N__8323\ : std_logic;
signal \N__8320\ : std_logic;
signal \N__8317\ : std_logic;
signal \N__8314\ : std_logic;
signal \N__8311\ : std_logic;
signal \N__8308\ : std_logic;
signal \N__8305\ : std_logic;
signal \N__8302\ : std_logic;
signal \N__8299\ : std_logic;
signal \N__8296\ : std_logic;
signal \N__8293\ : std_logic;
signal \N__8290\ : std_logic;
signal \N__8287\ : std_logic;
signal \N__8284\ : std_logic;
signal \N__8281\ : std_logic;
signal \N__8278\ : std_logic;
signal \N__8275\ : std_logic;
signal \N__8272\ : std_logic;
signal \N__8269\ : std_logic;
signal \N__8266\ : std_logic;
signal \N__8263\ : std_logic;
signal \N__8260\ : std_logic;
signal \N__8257\ : std_logic;
signal \N__8254\ : std_logic;
signal \N__8251\ : std_logic;
signal \N__8248\ : std_logic;
signal \N__8245\ : std_logic;
signal \N__8242\ : std_logic;
signal \N__8239\ : std_logic;
signal \N__8236\ : std_logic;
signal \N__8233\ : std_logic;
signal \N__8228\ : std_logic;
signal \N__8225\ : std_logic;
signal \N__8222\ : std_logic;
signal \N__8219\ : std_logic;
signal \N__8216\ : std_logic;
signal \N__8213\ : std_logic;
signal \N__8212\ : std_logic;
signal \N__8209\ : std_logic;
signal \N__8206\ : std_logic;
signal \N__8203\ : std_logic;
signal \N__8200\ : std_logic;
signal \N__8197\ : std_logic;
signal \N__8194\ : std_logic;
signal \N__8191\ : std_logic;
signal \N__8188\ : std_logic;
signal \N__8185\ : std_logic;
signal \N__8182\ : std_logic;
signal \N__8179\ : std_logic;
signal \N__8176\ : std_logic;
signal \N__8173\ : std_logic;
signal \N__8170\ : std_logic;
signal \N__8167\ : std_logic;
signal \N__8164\ : std_logic;
signal \N__8161\ : std_logic;
signal \N__8158\ : std_logic;
signal \N__8155\ : std_logic;
signal \N__8152\ : std_logic;
signal \N__8149\ : std_logic;
signal \N__8146\ : std_logic;
signal \N__8143\ : std_logic;
signal \N__8140\ : std_logic;
signal \N__8137\ : std_logic;
signal \N__8134\ : std_logic;
signal \N__8131\ : std_logic;
signal \N__8128\ : std_logic;
signal \N__8125\ : std_logic;
signal \N__8122\ : std_logic;
signal \N__8119\ : std_logic;
signal \N__8116\ : std_logic;
signal \N__8113\ : std_logic;
signal \N__8110\ : std_logic;
signal \N__8107\ : std_logic;
signal \N__8104\ : std_logic;
signal \N__8101\ : std_logic;
signal \N__8098\ : std_logic;
signal \N__8095\ : std_logic;
signal \N__8092\ : std_logic;
signal \N__8089\ : std_logic;
signal \N__8086\ : std_logic;
signal \N__8083\ : std_logic;
signal \N__8080\ : std_logic;
signal \N__8077\ : std_logic;
signal \N__8074\ : std_logic;
signal \N__8071\ : std_logic;
signal \N__8068\ : std_logic;
signal \N__8065\ : std_logic;
signal \N__8062\ : std_logic;
signal \N__8059\ : std_logic;
signal \N__8056\ : std_logic;
signal \N__8053\ : std_logic;
signal \N__8050\ : std_logic;
signal \N__8047\ : std_logic;
signal \N__8044\ : std_logic;
signal \N__8041\ : std_logic;
signal \N__8038\ : std_logic;
signal \N__8035\ : std_logic;
signal \N__8032\ : std_logic;
signal \N__8029\ : std_logic;
signal \N__8026\ : std_logic;
signal \N__8023\ : std_logic;
signal \N__8020\ : std_logic;
signal \N__8015\ : std_logic;
signal \N__8014\ : std_logic;
signal \N__8013\ : std_logic;
signal \N__8012\ : std_logic;
signal \N__8009\ : std_logic;
signal \N__8006\ : std_logic;
signal \N__8005\ : std_logic;
signal \N__8004\ : std_logic;
signal \N__8003\ : std_logic;
signal \N__8002\ : std_logic;
signal \N__7999\ : std_logic;
signal \N__7996\ : std_logic;
signal \N__7993\ : std_logic;
signal \N__7990\ : std_logic;
signal \N__7987\ : std_logic;
signal \N__7984\ : std_logic;
signal \N__7981\ : std_logic;
signal \N__7978\ : std_logic;
signal \N__7975\ : std_logic;
signal \N__7972\ : std_logic;
signal \N__7967\ : std_logic;
signal \N__7964\ : std_logic;
signal \N__7961\ : std_logic;
signal \N__7958\ : std_logic;
signal \N__7955\ : std_logic;
signal \N__7952\ : std_logic;
signal \N__7949\ : std_logic;
signal \N__7946\ : std_logic;
signal \N__7941\ : std_logic;
signal \N__7936\ : std_logic;
signal \N__7933\ : std_logic;
signal \N__7930\ : std_logic;
signal \N__7927\ : std_logic;
signal \N__7924\ : std_logic;
signal \N__7917\ : std_logic;
signal \N__7910\ : std_logic;
signal \N__7907\ : std_logic;
signal \N__7904\ : std_logic;
signal \N__7903\ : std_logic;
signal \N__7900\ : std_logic;
signal \N__7897\ : std_logic;
signal \N__7894\ : std_logic;
signal \N__7891\ : std_logic;
signal \N__7888\ : std_logic;
signal \N__7885\ : std_logic;
signal \N__7882\ : std_logic;
signal \N__7879\ : std_logic;
signal \N__7876\ : std_logic;
signal \N__7873\ : std_logic;
signal \N__7870\ : std_logic;
signal \N__7867\ : std_logic;
signal \N__7864\ : std_logic;
signal \N__7861\ : std_logic;
signal \N__7858\ : std_logic;
signal \N__7855\ : std_logic;
signal \N__7852\ : std_logic;
signal \N__7849\ : std_logic;
signal \N__7846\ : std_logic;
signal \N__7843\ : std_logic;
signal \N__7840\ : std_logic;
signal \N__7837\ : std_logic;
signal \N__7834\ : std_logic;
signal \N__7831\ : std_logic;
signal \N__7828\ : std_logic;
signal \N__7825\ : std_logic;
signal \N__7822\ : std_logic;
signal \N__7819\ : std_logic;
signal \N__7816\ : std_logic;
signal \N__7813\ : std_logic;
signal \N__7810\ : std_logic;
signal \N__7807\ : std_logic;
signal \N__7804\ : std_logic;
signal \N__7801\ : std_logic;
signal \N__7798\ : std_logic;
signal \N__7795\ : std_logic;
signal \N__7792\ : std_logic;
signal \N__7789\ : std_logic;
signal \N__7786\ : std_logic;
signal \N__7783\ : std_logic;
signal \N__7780\ : std_logic;
signal \N__7777\ : std_logic;
signal \N__7774\ : std_logic;
signal \N__7771\ : std_logic;
signal \N__7768\ : std_logic;
signal \N__7765\ : std_logic;
signal \N__7762\ : std_logic;
signal \N__7759\ : std_logic;
signal \N__7756\ : std_logic;
signal \N__7753\ : std_logic;
signal \N__7750\ : std_logic;
signal \N__7747\ : std_logic;
signal \N__7744\ : std_logic;
signal \N__7741\ : std_logic;
signal \N__7738\ : std_logic;
signal \N__7735\ : std_logic;
signal \N__7732\ : std_logic;
signal \N__7729\ : std_logic;
signal \N__7726\ : std_logic;
signal \N__7723\ : std_logic;
signal \N__7720\ : std_logic;
signal \N__7717\ : std_logic;
signal \N__7714\ : std_logic;
signal \N__7711\ : std_logic;
signal \N__7708\ : std_logic;
signal \N__7705\ : std_logic;
signal \N__7702\ : std_logic;
signal \N__7699\ : std_logic;
signal \N__7694\ : std_logic;
signal \N__7691\ : std_logic;
signal \N__7688\ : std_logic;
signal \N__7685\ : std_logic;
signal \N__7682\ : std_logic;
signal \N__7681\ : std_logic;
signal \N__7678\ : std_logic;
signal \N__7675\ : std_logic;
signal \N__7672\ : std_logic;
signal \N__7669\ : std_logic;
signal \N__7666\ : std_logic;
signal \N__7663\ : std_logic;
signal \N__7660\ : std_logic;
signal \N__7657\ : std_logic;
signal \N__7654\ : std_logic;
signal \N__7651\ : std_logic;
signal \N__7648\ : std_logic;
signal \N__7645\ : std_logic;
signal \N__7642\ : std_logic;
signal \N__7639\ : std_logic;
signal \N__7636\ : std_logic;
signal \N__7633\ : std_logic;
signal \N__7630\ : std_logic;
signal \N__7627\ : std_logic;
signal \N__7624\ : std_logic;
signal \N__7621\ : std_logic;
signal \N__7618\ : std_logic;
signal \N__7615\ : std_logic;
signal \N__7612\ : std_logic;
signal \N__7609\ : std_logic;
signal \N__7606\ : std_logic;
signal \N__7603\ : std_logic;
signal \N__7600\ : std_logic;
signal \N__7597\ : std_logic;
signal \N__7594\ : std_logic;
signal \N__7591\ : std_logic;
signal \N__7588\ : std_logic;
signal \N__7585\ : std_logic;
signal \N__7582\ : std_logic;
signal \N__7579\ : std_logic;
signal \N__7576\ : std_logic;
signal \N__7573\ : std_logic;
signal \N__7570\ : std_logic;
signal \N__7567\ : std_logic;
signal \N__7564\ : std_logic;
signal \N__7561\ : std_logic;
signal \N__7558\ : std_logic;
signal \N__7555\ : std_logic;
signal \N__7552\ : std_logic;
signal \N__7549\ : std_logic;
signal \N__7546\ : std_logic;
signal \N__7543\ : std_logic;
signal \N__7540\ : std_logic;
signal \N__7537\ : std_logic;
signal \N__7534\ : std_logic;
signal \N__7531\ : std_logic;
signal \N__7528\ : std_logic;
signal \N__7525\ : std_logic;
signal \N__7522\ : std_logic;
signal \N__7519\ : std_logic;
signal \N__7516\ : std_logic;
signal \N__7513\ : std_logic;
signal \N__7510\ : std_logic;
signal \N__7507\ : std_logic;
signal \N__7504\ : std_logic;
signal \N__7501\ : std_logic;
signal \N__7498\ : std_logic;
signal \N__7495\ : std_logic;
signal \N__7492\ : std_logic;
signal \N__7489\ : std_logic;
signal \N__7486\ : std_logic;
signal \N__7483\ : std_logic;
signal \N__7480\ : std_logic;
signal \N__7477\ : std_logic;
signal \N__7472\ : std_logic;
signal \N__7469\ : std_logic;
signal \N__7466\ : std_logic;
signal \N__7463\ : std_logic;
signal \N__7462\ : std_logic;
signal \N__7459\ : std_logic;
signal \N__7456\ : std_logic;
signal \N__7453\ : std_logic;
signal \N__7450\ : std_logic;
signal \N__7447\ : std_logic;
signal \N__7444\ : std_logic;
signal \N__7441\ : std_logic;
signal \N__7438\ : std_logic;
signal \N__7435\ : std_logic;
signal \N__7432\ : std_logic;
signal \N__7429\ : std_logic;
signal \N__7426\ : std_logic;
signal \N__7423\ : std_logic;
signal \N__7420\ : std_logic;
signal \N__7417\ : std_logic;
signal \N__7414\ : std_logic;
signal \N__7411\ : std_logic;
signal \N__7408\ : std_logic;
signal \N__7405\ : std_logic;
signal \N__7402\ : std_logic;
signal \N__7399\ : std_logic;
signal \N__7396\ : std_logic;
signal \N__7393\ : std_logic;
signal \N__7390\ : std_logic;
signal \N__7387\ : std_logic;
signal \N__7384\ : std_logic;
signal \N__7381\ : std_logic;
signal \N__7378\ : std_logic;
signal \N__7375\ : std_logic;
signal \N__7372\ : std_logic;
signal \N__7369\ : std_logic;
signal \N__7366\ : std_logic;
signal \N__7363\ : std_logic;
signal \N__7360\ : std_logic;
signal \N__7357\ : std_logic;
signal \N__7354\ : std_logic;
signal \N__7351\ : std_logic;
signal \N__7348\ : std_logic;
signal \N__7345\ : std_logic;
signal \N__7342\ : std_logic;
signal \N__7339\ : std_logic;
signal \N__7336\ : std_logic;
signal \N__7333\ : std_logic;
signal \N__7330\ : std_logic;
signal \N__7327\ : std_logic;
signal \N__7324\ : std_logic;
signal \N__7321\ : std_logic;
signal \N__7318\ : std_logic;
signal \N__7315\ : std_logic;
signal \N__7312\ : std_logic;
signal \N__7309\ : std_logic;
signal \N__7306\ : std_logic;
signal \N__7303\ : std_logic;
signal \N__7300\ : std_logic;
signal \N__7297\ : std_logic;
signal \N__7294\ : std_logic;
signal \N__7291\ : std_logic;
signal \N__7288\ : std_logic;
signal \N__7285\ : std_logic;
signal \N__7282\ : std_logic;
signal \N__7279\ : std_logic;
signal \N__7276\ : std_logic;
signal \N__7273\ : std_logic;
signal \N__7270\ : std_logic;
signal \N__7267\ : std_logic;
signal \N__7264\ : std_logic;
signal \N__7261\ : std_logic;
signal \N__7258\ : std_logic;
signal \N__7253\ : std_logic;
signal \N__7250\ : std_logic;
signal \N__7249\ : std_logic;
signal \N__7246\ : std_logic;
signal \N__7243\ : std_logic;
signal \N__7240\ : std_logic;
signal \N__7237\ : std_logic;
signal \N__7234\ : std_logic;
signal \N__7231\ : std_logic;
signal \N__7228\ : std_logic;
signal \N__7225\ : std_logic;
signal \N__7222\ : std_logic;
signal \N__7219\ : std_logic;
signal \N__7216\ : std_logic;
signal \N__7213\ : std_logic;
signal \N__7210\ : std_logic;
signal \N__7207\ : std_logic;
signal \N__7204\ : std_logic;
signal \N__7201\ : std_logic;
signal \N__7198\ : std_logic;
signal \N__7195\ : std_logic;
signal \N__7192\ : std_logic;
signal \N__7189\ : std_logic;
signal \N__7186\ : std_logic;
signal \N__7183\ : std_logic;
signal \N__7180\ : std_logic;
signal \N__7177\ : std_logic;
signal \N__7174\ : std_logic;
signal \N__7171\ : std_logic;
signal \N__7168\ : std_logic;
signal \N__7165\ : std_logic;
signal \N__7162\ : std_logic;
signal \N__7159\ : std_logic;
signal \N__7156\ : std_logic;
signal \N__7153\ : std_logic;
signal \N__7150\ : std_logic;
signal \N__7147\ : std_logic;
signal \N__7144\ : std_logic;
signal \N__7141\ : std_logic;
signal \N__7138\ : std_logic;
signal \N__7135\ : std_logic;
signal \N__7132\ : std_logic;
signal \N__7129\ : std_logic;
signal \N__7126\ : std_logic;
signal \N__7123\ : std_logic;
signal \N__7120\ : std_logic;
signal \N__7117\ : std_logic;
signal \N__7114\ : std_logic;
signal \N__7111\ : std_logic;
signal \N__7108\ : std_logic;
signal \N__7105\ : std_logic;
signal \N__7102\ : std_logic;
signal \N__7099\ : std_logic;
signal \N__7096\ : std_logic;
signal \N__7093\ : std_logic;
signal \N__7090\ : std_logic;
signal \N__7087\ : std_logic;
signal \N__7084\ : std_logic;
signal \N__7081\ : std_logic;
signal \N__7078\ : std_logic;
signal \N__7075\ : std_logic;
signal \N__7072\ : std_logic;
signal \N__7069\ : std_logic;
signal \N__7066\ : std_logic;
signal \N__7063\ : std_logic;
signal \N__7060\ : std_logic;
signal \N__7057\ : std_logic;
signal \N__7054\ : std_logic;
signal \N__7051\ : std_logic;
signal \N__7048\ : std_logic;
signal \N__7045\ : std_logic;
signal \N__7042\ : std_logic;
signal \N__7039\ : std_logic;
signal \N__7036\ : std_logic;
signal \N__7033\ : std_logic;
signal \N__7028\ : std_logic;
signal \N__7025\ : std_logic;
signal \N__7022\ : std_logic;
signal \N__7019\ : std_logic;
signal \N__7016\ : std_logic;
signal \N__7015\ : std_logic;
signal \N__7012\ : std_logic;
signal \N__7009\ : std_logic;
signal \N__7006\ : std_logic;
signal \N__7003\ : std_logic;
signal \N__7000\ : std_logic;
signal \N__6997\ : std_logic;
signal \N__6994\ : std_logic;
signal \N__6991\ : std_logic;
signal \N__6988\ : std_logic;
signal \N__6985\ : std_logic;
signal \N__6982\ : std_logic;
signal \N__6979\ : std_logic;
signal \N__6976\ : std_logic;
signal \N__6973\ : std_logic;
signal \N__6970\ : std_logic;
signal \N__6967\ : std_logic;
signal \N__6964\ : std_logic;
signal \N__6961\ : std_logic;
signal \N__6958\ : std_logic;
signal \N__6955\ : std_logic;
signal \N__6952\ : std_logic;
signal \N__6949\ : std_logic;
signal \N__6946\ : std_logic;
signal \N__6943\ : std_logic;
signal \N__6940\ : std_logic;
signal \N__6937\ : std_logic;
signal \N__6934\ : std_logic;
signal \N__6931\ : std_logic;
signal \N__6928\ : std_logic;
signal \N__6925\ : std_logic;
signal \N__6922\ : std_logic;
signal \N__6919\ : std_logic;
signal \N__6916\ : std_logic;
signal \N__6913\ : std_logic;
signal \N__6910\ : std_logic;
signal \N__6907\ : std_logic;
signal \N__6904\ : std_logic;
signal \N__6901\ : std_logic;
signal \N__6898\ : std_logic;
signal \N__6895\ : std_logic;
signal \N__6892\ : std_logic;
signal \N__6889\ : std_logic;
signal \N__6886\ : std_logic;
signal \N__6883\ : std_logic;
signal \N__6880\ : std_logic;
signal \N__6877\ : std_logic;
signal \N__6874\ : std_logic;
signal \N__6871\ : std_logic;
signal \N__6868\ : std_logic;
signal \N__6865\ : std_logic;
signal \N__6862\ : std_logic;
signal \N__6859\ : std_logic;
signal \N__6856\ : std_logic;
signal \N__6853\ : std_logic;
signal \N__6850\ : std_logic;
signal \N__6847\ : std_logic;
signal \N__6844\ : std_logic;
signal \N__6841\ : std_logic;
signal \N__6838\ : std_logic;
signal \N__6835\ : std_logic;
signal \N__6832\ : std_logic;
signal \N__6829\ : std_logic;
signal \N__6826\ : std_logic;
signal \N__6823\ : std_logic;
signal \N__6820\ : std_logic;
signal \N__6817\ : std_logic;
signal \N__6812\ : std_logic;
signal \N__6809\ : std_logic;
signal \N__6806\ : std_logic;
signal \N__6803\ : std_logic;
signal \N__6800\ : std_logic;
signal \N__6799\ : std_logic;
signal \N__6796\ : std_logic;
signal \N__6793\ : std_logic;
signal \N__6790\ : std_logic;
signal \N__6787\ : std_logic;
signal \N__6784\ : std_logic;
signal \N__6781\ : std_logic;
signal \N__6778\ : std_logic;
signal \N__6775\ : std_logic;
signal \N__6772\ : std_logic;
signal \N__6769\ : std_logic;
signal \N__6766\ : std_logic;
signal \N__6763\ : std_logic;
signal \N__6760\ : std_logic;
signal \N__6757\ : std_logic;
signal \N__6754\ : std_logic;
signal \N__6751\ : std_logic;
signal \N__6748\ : std_logic;
signal \N__6745\ : std_logic;
signal \N__6742\ : std_logic;
signal \N__6739\ : std_logic;
signal \N__6736\ : std_logic;
signal \N__6733\ : std_logic;
signal \N__6730\ : std_logic;
signal \N__6727\ : std_logic;
signal \N__6724\ : std_logic;
signal \N__6721\ : std_logic;
signal \N__6718\ : std_logic;
signal \N__6715\ : std_logic;
signal \N__6712\ : std_logic;
signal \N__6709\ : std_logic;
signal \N__6706\ : std_logic;
signal \N__6703\ : std_logic;
signal \N__6700\ : std_logic;
signal \N__6697\ : std_logic;
signal \N__6694\ : std_logic;
signal \N__6691\ : std_logic;
signal \N__6688\ : std_logic;
signal \N__6685\ : std_logic;
signal \N__6682\ : std_logic;
signal \N__6679\ : std_logic;
signal \N__6676\ : std_logic;
signal \N__6673\ : std_logic;
signal \N__6670\ : std_logic;
signal \N__6667\ : std_logic;
signal \N__6664\ : std_logic;
signal \N__6661\ : std_logic;
signal \N__6658\ : std_logic;
signal \N__6655\ : std_logic;
signal \N__6652\ : std_logic;
signal \N__6649\ : std_logic;
signal \N__6646\ : std_logic;
signal \N__6643\ : std_logic;
signal \N__6640\ : std_logic;
signal \N__6637\ : std_logic;
signal \N__6634\ : std_logic;
signal \N__6631\ : std_logic;
signal \N__6628\ : std_logic;
signal \N__6625\ : std_logic;
signal \N__6622\ : std_logic;
signal \N__6619\ : std_logic;
signal \N__6616\ : std_logic;
signal \N__6613\ : std_logic;
signal \N__6610\ : std_logic;
signal \N__6607\ : std_logic;
signal \N__6604\ : std_logic;
signal \N__6601\ : std_logic;
signal \N__6596\ : std_logic;
signal \N__6593\ : std_logic;
signal \N__6590\ : std_logic;
signal \N__6587\ : std_logic;
signal \N__6584\ : std_logic;
signal \N__6583\ : std_logic;
signal \N__6580\ : std_logic;
signal \N__6577\ : std_logic;
signal \N__6574\ : std_logic;
signal \N__6571\ : std_logic;
signal \N__6568\ : std_logic;
signal \N__6565\ : std_logic;
signal \N__6562\ : std_logic;
signal \N__6559\ : std_logic;
signal \N__6556\ : std_logic;
signal \N__6553\ : std_logic;
signal \N__6550\ : std_logic;
signal \N__6547\ : std_logic;
signal \N__6544\ : std_logic;
signal \N__6541\ : std_logic;
signal \N__6538\ : std_logic;
signal \N__6535\ : std_logic;
signal \N__6532\ : std_logic;
signal \N__6529\ : std_logic;
signal \N__6526\ : std_logic;
signal \N__6523\ : std_logic;
signal \N__6520\ : std_logic;
signal \N__6517\ : std_logic;
signal \N__6514\ : std_logic;
signal \N__6511\ : std_logic;
signal \N__6508\ : std_logic;
signal \N__6505\ : std_logic;
signal \N__6502\ : std_logic;
signal \N__6499\ : std_logic;
signal \N__6496\ : std_logic;
signal \N__6493\ : std_logic;
signal \N__6490\ : std_logic;
signal \N__6487\ : std_logic;
signal \N__6484\ : std_logic;
signal \N__6481\ : std_logic;
signal \N__6478\ : std_logic;
signal \N__6475\ : std_logic;
signal \N__6472\ : std_logic;
signal \N__6469\ : std_logic;
signal \N__6466\ : std_logic;
signal \N__6463\ : std_logic;
signal \N__6460\ : std_logic;
signal \N__6457\ : std_logic;
signal \N__6454\ : std_logic;
signal \N__6451\ : std_logic;
signal \N__6448\ : std_logic;
signal \N__6445\ : std_logic;
signal \N__6442\ : std_logic;
signal \N__6439\ : std_logic;
signal \N__6436\ : std_logic;
signal \N__6433\ : std_logic;
signal \N__6430\ : std_logic;
signal \N__6427\ : std_logic;
signal \N__6424\ : std_logic;
signal \N__6421\ : std_logic;
signal \N__6418\ : std_logic;
signal \N__6415\ : std_logic;
signal \N__6412\ : std_logic;
signal \N__6409\ : std_logic;
signal \N__6406\ : std_logic;
signal \N__6403\ : std_logic;
signal \N__6400\ : std_logic;
signal \N__6397\ : std_logic;
signal \N__6394\ : std_logic;
signal \N__6391\ : std_logic;
signal \N__6388\ : std_logic;
signal \N__6385\ : std_logic;
signal \N__6380\ : std_logic;
signal \N__6377\ : std_logic;
signal \N__6374\ : std_logic;
signal \N__6371\ : std_logic;
signal \N__6368\ : std_logic;
signal \N__6367\ : std_logic;
signal \N__6364\ : std_logic;
signal \N__6361\ : std_logic;
signal \N__6358\ : std_logic;
signal \N__6355\ : std_logic;
signal \N__6352\ : std_logic;
signal \N__6349\ : std_logic;
signal \N__6346\ : std_logic;
signal \N__6343\ : std_logic;
signal \N__6340\ : std_logic;
signal \N__6337\ : std_logic;
signal \N__6334\ : std_logic;
signal \N__6331\ : std_logic;
signal \N__6328\ : std_logic;
signal \N__6325\ : std_logic;
signal \N__6322\ : std_logic;
signal \N__6319\ : std_logic;
signal \N__6316\ : std_logic;
signal \N__6313\ : std_logic;
signal \N__6310\ : std_logic;
signal \N__6307\ : std_logic;
signal \N__6304\ : std_logic;
signal \N__6301\ : std_logic;
signal \N__6298\ : std_logic;
signal \N__6295\ : std_logic;
signal \N__6292\ : std_logic;
signal \N__6289\ : std_logic;
signal \N__6286\ : std_logic;
signal \N__6283\ : std_logic;
signal \N__6280\ : std_logic;
signal \N__6277\ : std_logic;
signal \N__6274\ : std_logic;
signal \N__6271\ : std_logic;
signal \N__6268\ : std_logic;
signal \N__6265\ : std_logic;
signal \N__6262\ : std_logic;
signal \N__6259\ : std_logic;
signal \N__6256\ : std_logic;
signal \N__6253\ : std_logic;
signal \N__6250\ : std_logic;
signal \N__6247\ : std_logic;
signal \N__6244\ : std_logic;
signal \N__6241\ : std_logic;
signal \N__6238\ : std_logic;
signal \N__6235\ : std_logic;
signal \N__6232\ : std_logic;
signal \N__6229\ : std_logic;
signal \N__6226\ : std_logic;
signal \N__6223\ : std_logic;
signal \N__6220\ : std_logic;
signal \N__6217\ : std_logic;
signal \N__6214\ : std_logic;
signal \N__6211\ : std_logic;
signal \N__6208\ : std_logic;
signal \N__6205\ : std_logic;
signal \N__6202\ : std_logic;
signal \N__6199\ : std_logic;
signal \N__6196\ : std_logic;
signal \N__6193\ : std_logic;
signal \N__6190\ : std_logic;
signal \N__6187\ : std_logic;
signal \N__6184\ : std_logic;
signal \N__6181\ : std_logic;
signal \N__6178\ : std_logic;
signal \N__6175\ : std_logic;
signal \N__6172\ : std_logic;
signal \N__6169\ : std_logic;
signal \N__6166\ : std_logic;
signal \N__6163\ : std_logic;
signal \N__6158\ : std_logic;
signal \N__6155\ : std_logic;
signal \N__6152\ : std_logic;
signal \N__6149\ : std_logic;
signal \N__6146\ : std_logic;
signal \N__6145\ : std_logic;
signal \N__6142\ : std_logic;
signal \N__6139\ : std_logic;
signal \N__6136\ : std_logic;
signal \N__6133\ : std_logic;
signal \N__6130\ : std_logic;
signal \N__6127\ : std_logic;
signal \N__6124\ : std_logic;
signal \N__6121\ : std_logic;
signal \N__6118\ : std_logic;
signal \N__6115\ : std_logic;
signal \N__6112\ : std_logic;
signal \N__6109\ : std_logic;
signal \N__6106\ : std_logic;
signal \N__6103\ : std_logic;
signal \N__6100\ : std_logic;
signal \N__6097\ : std_logic;
signal \N__6094\ : std_logic;
signal \N__6091\ : std_logic;
signal \N__6088\ : std_logic;
signal \N__6085\ : std_logic;
signal \N__6082\ : std_logic;
signal \N__6079\ : std_logic;
signal \N__6076\ : std_logic;
signal \N__6073\ : std_logic;
signal \N__6070\ : std_logic;
signal \N__6067\ : std_logic;
signal \N__6064\ : std_logic;
signal \N__6061\ : std_logic;
signal \N__6058\ : std_logic;
signal \N__6055\ : std_logic;
signal \N__6052\ : std_logic;
signal \N__6049\ : std_logic;
signal \N__6046\ : std_logic;
signal \N__6043\ : std_logic;
signal \N__6040\ : std_logic;
signal \N__6037\ : std_logic;
signal \N__6034\ : std_logic;
signal \N__6031\ : std_logic;
signal \N__6028\ : std_logic;
signal \N__6025\ : std_logic;
signal \N__6022\ : std_logic;
signal \N__6019\ : std_logic;
signal \N__6016\ : std_logic;
signal \N__6013\ : std_logic;
signal \N__6010\ : std_logic;
signal \N__6007\ : std_logic;
signal \N__6004\ : std_logic;
signal \N__6001\ : std_logic;
signal \N__5998\ : std_logic;
signal \N__5995\ : std_logic;
signal \N__5992\ : std_logic;
signal \N__5989\ : std_logic;
signal \N__5986\ : std_logic;
signal \N__5983\ : std_logic;
signal \N__5980\ : std_logic;
signal \N__5977\ : std_logic;
signal \N__5974\ : std_logic;
signal \N__5971\ : std_logic;
signal \N__5968\ : std_logic;
signal \N__5965\ : std_logic;
signal \N__5962\ : std_logic;
signal \N__5959\ : std_logic;
signal \N__5956\ : std_logic;
signal \N__5953\ : std_logic;
signal \N__5948\ : std_logic;
signal \N__5945\ : std_logic;
signal \N__5942\ : std_logic;
signal \N__5939\ : std_logic;
signal \N__5936\ : std_logic;
signal \N__5933\ : std_logic;
signal \N__5930\ : std_logic;
signal \N__5929\ : std_logic;
signal \N__5926\ : std_logic;
signal \N__5923\ : std_logic;
signal \N__5920\ : std_logic;
signal \N__5917\ : std_logic;
signal \N__5914\ : std_logic;
signal \N__5911\ : std_logic;
signal \N__5908\ : std_logic;
signal \N__5905\ : std_logic;
signal \N__5902\ : std_logic;
signal \N__5899\ : std_logic;
signal \N__5896\ : std_logic;
signal \N__5893\ : std_logic;
signal \N__5890\ : std_logic;
signal \N__5887\ : std_logic;
signal \N__5884\ : std_logic;
signal \N__5881\ : std_logic;
signal \N__5878\ : std_logic;
signal \N__5875\ : std_logic;
signal \N__5872\ : std_logic;
signal \N__5869\ : std_logic;
signal \N__5866\ : std_logic;
signal \N__5863\ : std_logic;
signal \N__5860\ : std_logic;
signal \N__5857\ : std_logic;
signal \N__5854\ : std_logic;
signal \N__5851\ : std_logic;
signal \N__5848\ : std_logic;
signal \N__5845\ : std_logic;
signal \N__5842\ : std_logic;
signal \N__5839\ : std_logic;
signal \N__5836\ : std_logic;
signal \N__5833\ : std_logic;
signal \N__5830\ : std_logic;
signal \N__5827\ : std_logic;
signal \N__5824\ : std_logic;
signal \N__5821\ : std_logic;
signal \N__5818\ : std_logic;
signal \N__5815\ : std_logic;
signal \N__5812\ : std_logic;
signal \N__5809\ : std_logic;
signal \N__5806\ : std_logic;
signal \N__5803\ : std_logic;
signal \N__5800\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5794\ : std_logic;
signal \N__5791\ : std_logic;
signal \N__5788\ : std_logic;
signal \N__5785\ : std_logic;
signal \N__5782\ : std_logic;
signal \N__5779\ : std_logic;
signal \N__5776\ : std_logic;
signal \N__5773\ : std_logic;
signal \N__5770\ : std_logic;
signal \N__5767\ : std_logic;
signal \N__5764\ : std_logic;
signal \N__5761\ : std_logic;
signal \N__5758\ : std_logic;
signal \N__5755\ : std_logic;
signal \N__5752\ : std_logic;
signal \N__5749\ : std_logic;
signal \N__5746\ : std_logic;
signal \N__5743\ : std_logic;
signal \N__5740\ : std_logic;
signal \N__5737\ : std_logic;
signal \N__5734\ : std_logic;
signal \N__5731\ : std_logic;
signal \N__5726\ : std_logic;
signal \N__5723\ : std_logic;
signal \N__5720\ : std_logic;
signal \N__5719\ : std_logic;
signal \N__5716\ : std_logic;
signal \N__5713\ : std_logic;
signal \N__5710\ : std_logic;
signal \N__5707\ : std_logic;
signal \N__5704\ : std_logic;
signal \N__5701\ : std_logic;
signal \N__5698\ : std_logic;
signal \N__5695\ : std_logic;
signal \N__5692\ : std_logic;
signal \N__5689\ : std_logic;
signal \N__5686\ : std_logic;
signal \N__5683\ : std_logic;
signal \N__5680\ : std_logic;
signal \N__5677\ : std_logic;
signal \N__5674\ : std_logic;
signal \N__5671\ : std_logic;
signal \N__5668\ : std_logic;
signal \N__5665\ : std_logic;
signal \N__5662\ : std_logic;
signal \N__5659\ : std_logic;
signal \N__5656\ : std_logic;
signal \N__5653\ : std_logic;
signal \N__5650\ : std_logic;
signal \N__5647\ : std_logic;
signal \N__5644\ : std_logic;
signal \N__5641\ : std_logic;
signal \N__5638\ : std_logic;
signal \N__5635\ : std_logic;
signal \N__5632\ : std_logic;
signal \N__5629\ : std_logic;
signal \N__5626\ : std_logic;
signal \N__5623\ : std_logic;
signal \N__5620\ : std_logic;
signal \N__5617\ : std_logic;
signal \N__5614\ : std_logic;
signal \N__5611\ : std_logic;
signal \N__5608\ : std_logic;
signal \N__5605\ : std_logic;
signal \N__5602\ : std_logic;
signal \N__5599\ : std_logic;
signal \N__5596\ : std_logic;
signal \N__5593\ : std_logic;
signal \N__5590\ : std_logic;
signal \N__5587\ : std_logic;
signal \N__5584\ : std_logic;
signal \N__5581\ : std_logic;
signal \N__5578\ : std_logic;
signal \N__5575\ : std_logic;
signal \N__5572\ : std_logic;
signal \N__5569\ : std_logic;
signal \N__5566\ : std_logic;
signal \N__5563\ : std_logic;
signal \N__5560\ : std_logic;
signal \N__5557\ : std_logic;
signal \N__5554\ : std_logic;
signal \N__5551\ : std_logic;
signal \N__5548\ : std_logic;
signal \N__5545\ : std_logic;
signal \N__5542\ : std_logic;
signal \N__5539\ : std_logic;
signal \N__5536\ : std_logic;
signal \N__5533\ : std_logic;
signal \N__5530\ : std_logic;
signal \N__5527\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5521\ : std_logic;
signal \N__5518\ : std_logic;
signal \N__5515\ : std_logic;
signal \N__5512\ : std_logic;
signal \N__5509\ : std_logic;
signal \N__5506\ : std_logic;
signal \N__5503\ : std_logic;
signal \N__5498\ : std_logic;
signal \N__5495\ : std_logic;
signal \N__5492\ : std_logic;
signal \N__5491\ : std_logic;
signal \N__5488\ : std_logic;
signal \N__5485\ : std_logic;
signal \N__5482\ : std_logic;
signal \N__5479\ : std_logic;
signal \N__5476\ : std_logic;
signal \N__5473\ : std_logic;
signal \N__5470\ : std_logic;
signal \N__5467\ : std_logic;
signal \N__5464\ : std_logic;
signal \N__5461\ : std_logic;
signal \N__5458\ : std_logic;
signal \N__5455\ : std_logic;
signal \N__5452\ : std_logic;
signal \N__5449\ : std_logic;
signal \N__5446\ : std_logic;
signal \N__5443\ : std_logic;
signal \N__5440\ : std_logic;
signal \N__5437\ : std_logic;
signal \N__5434\ : std_logic;
signal \N__5431\ : std_logic;
signal \N__5428\ : std_logic;
signal \N__5425\ : std_logic;
signal \N__5422\ : std_logic;
signal \N__5419\ : std_logic;
signal \N__5416\ : std_logic;
signal \N__5413\ : std_logic;
signal \N__5410\ : std_logic;
signal \N__5407\ : std_logic;
signal \N__5404\ : std_logic;
signal \N__5401\ : std_logic;
signal \N__5398\ : std_logic;
signal \N__5395\ : std_logic;
signal \N__5392\ : std_logic;
signal \N__5389\ : std_logic;
signal \N__5386\ : std_logic;
signal \N__5383\ : std_logic;
signal \N__5380\ : std_logic;
signal \N__5377\ : std_logic;
signal \N__5374\ : std_logic;
signal \N__5371\ : std_logic;
signal \N__5368\ : std_logic;
signal \N__5365\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5359\ : std_logic;
signal \N__5356\ : std_logic;
signal \N__5353\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5347\ : std_logic;
signal \N__5344\ : std_logic;
signal \N__5341\ : std_logic;
signal \N__5338\ : std_logic;
signal \N__5335\ : std_logic;
signal \N__5332\ : std_logic;
signal \N__5329\ : std_logic;
signal \N__5326\ : std_logic;
signal \N__5323\ : std_logic;
signal \N__5320\ : std_logic;
signal \N__5317\ : std_logic;
signal \N__5314\ : std_logic;
signal \N__5311\ : std_logic;
signal \N__5308\ : std_logic;
signal \N__5305\ : std_logic;
signal \N__5302\ : std_logic;
signal \N__5299\ : std_logic;
signal \N__5296\ : std_logic;
signal \N__5293\ : std_logic;
signal \N__5290\ : std_logic;
signal \N__5287\ : std_logic;
signal \N__5284\ : std_logic;
signal \N__5281\ : std_logic;
signal \N__5278\ : std_logic;
signal \N__5275\ : std_logic;
signal \N__5270\ : std_logic;
signal \N__5267\ : std_logic;
signal \N__5264\ : std_logic;
signal \N__5261\ : std_logic;
signal \N__5258\ : std_logic;
signal \N__5257\ : std_logic;
signal \N__5254\ : std_logic;
signal \N__5251\ : std_logic;
signal \N__5248\ : std_logic;
signal \N__5245\ : std_logic;
signal \N__5242\ : std_logic;
signal \N__5239\ : std_logic;
signal \N__5236\ : std_logic;
signal \N__5233\ : std_logic;
signal \N__5230\ : std_logic;
signal \N__5227\ : std_logic;
signal \N__5224\ : std_logic;
signal \N__5221\ : std_logic;
signal \N__5218\ : std_logic;
signal \N__5215\ : std_logic;
signal \N__5212\ : std_logic;
signal \N__5209\ : std_logic;
signal \N__5206\ : std_logic;
signal \N__5203\ : std_logic;
signal \N__5200\ : std_logic;
signal \N__5197\ : std_logic;
signal \N__5194\ : std_logic;
signal \N__5191\ : std_logic;
signal \N__5188\ : std_logic;
signal \N__5185\ : std_logic;
signal \N__5182\ : std_logic;
signal \N__5179\ : std_logic;
signal \N__5176\ : std_logic;
signal \N__5173\ : std_logic;
signal \N__5170\ : std_logic;
signal \N__5167\ : std_logic;
signal \N__5164\ : std_logic;
signal \N__5161\ : std_logic;
signal \N__5158\ : std_logic;
signal \N__5155\ : std_logic;
signal \N__5152\ : std_logic;
signal \N__5149\ : std_logic;
signal \N__5146\ : std_logic;
signal \N__5143\ : std_logic;
signal \N__5140\ : std_logic;
signal \N__5137\ : std_logic;
signal \N__5134\ : std_logic;
signal \N__5131\ : std_logic;
signal \N__5128\ : std_logic;
signal \N__5125\ : std_logic;
signal \N__5122\ : std_logic;
signal \N__5119\ : std_logic;
signal \N__5116\ : std_logic;
signal \N__5113\ : std_logic;
signal \N__5110\ : std_logic;
signal \N__5107\ : std_logic;
signal \N__5104\ : std_logic;
signal \N__5101\ : std_logic;
signal \N__5098\ : std_logic;
signal \N__5095\ : std_logic;
signal \N__5092\ : std_logic;
signal \N__5089\ : std_logic;
signal \N__5086\ : std_logic;
signal \N__5083\ : std_logic;
signal \N__5080\ : std_logic;
signal \N__5077\ : std_logic;
signal \N__5074\ : std_logic;
signal \N__5071\ : std_logic;
signal \N__5068\ : std_logic;
signal \N__5065\ : std_logic;
signal \N__5060\ : std_logic;
signal \N__5057\ : std_logic;
signal \N__5054\ : std_logic;
signal \N__5051\ : std_logic;
signal \N__5050\ : std_logic;
signal \N__5047\ : std_logic;
signal \N__5044\ : std_logic;
signal \N__5041\ : std_logic;
signal \N__5040\ : std_logic;
signal \N__5037\ : std_logic;
signal \N__5036\ : std_logic;
signal \N__5033\ : std_logic;
signal \N__5030\ : std_logic;
signal \N__5027\ : std_logic;
signal \N__5024\ : std_logic;
signal \N__5019\ : std_logic;
signal \N__5018\ : std_logic;
signal \N__5015\ : std_logic;
signal \N__5012\ : std_logic;
signal \N__5011\ : std_logic;
signal \N__5008\ : std_logic;
signal \N__5005\ : std_logic;
signal \N__5000\ : std_logic;
signal \N__4997\ : std_logic;
signal \N__4992\ : std_logic;
signal \N__4991\ : std_logic;
signal \N__4988\ : std_logic;
signal \N__4985\ : std_logic;
signal \N__4984\ : std_logic;
signal \N__4981\ : std_logic;
signal \N__4978\ : std_logic;
signal \N__4973\ : std_logic;
signal \N__4970\ : std_logic;
signal \N__4965\ : std_logic;
signal \N__4962\ : std_logic;
signal \N__4959\ : std_logic;
signal \N__4956\ : std_logic;
signal \N__4951\ : std_logic;
signal \N__4948\ : std_logic;
signal \N__4945\ : std_logic;
signal \N__4942\ : std_logic;
signal \N__4939\ : std_logic;
signal \N__4934\ : std_logic;
signal \N__4933\ : std_logic;
signal \N__4932\ : std_logic;
signal \N__4931\ : std_logic;
signal \N__4930\ : std_logic;
signal \N__4929\ : std_logic;
signal \N__4928\ : std_logic;
signal \N__4927\ : std_logic;
signal \N__4926\ : std_logic;
signal \N__4925\ : std_logic;
signal \N__4924\ : std_logic;
signal \N__4923\ : std_logic;
signal \N__4922\ : std_logic;
signal \N__4921\ : std_logic;
signal \N__4920\ : std_logic;
signal \N__4919\ : std_logic;
signal \N__4918\ : std_logic;
signal \N__4917\ : std_logic;
signal \N__4916\ : std_logic;
signal \N__4915\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4913\ : std_logic;
signal \N__4912\ : std_logic;
signal \N__4911\ : std_logic;
signal \N__4910\ : std_logic;
signal \N__4909\ : std_logic;
signal \N__4908\ : std_logic;
signal \N__4907\ : std_logic;
signal \N__4906\ : std_logic;
signal \N__4905\ : std_logic;
signal \N__4904\ : std_logic;
signal \N__4903\ : std_logic;
signal \N__4902\ : std_logic;
signal \N__4901\ : std_logic;
signal \N__4900\ : std_logic;
signal \N__4829\ : std_logic;
signal \N__4826\ : std_logic;
signal \N__4823\ : std_logic;
signal \N__4820\ : std_logic;
signal \N__4817\ : std_logic;
signal \N__4814\ : std_logic;
signal \N__4811\ : std_logic;
signal \N__4810\ : std_logic;
signal \N__4807\ : std_logic;
signal \N__4804\ : std_logic;
signal \N__4801\ : std_logic;
signal \N__4798\ : std_logic;
signal \N__4795\ : std_logic;
signal \N__4792\ : std_logic;
signal \N__4789\ : std_logic;
signal \N__4786\ : std_logic;
signal \N__4783\ : std_logic;
signal \N__4780\ : std_logic;
signal \N__4777\ : std_logic;
signal \N__4774\ : std_logic;
signal \N__4771\ : std_logic;
signal \N__4768\ : std_logic;
signal \N__4765\ : std_logic;
signal \N__4762\ : std_logic;
signal \N__4759\ : std_logic;
signal \N__4756\ : std_logic;
signal \N__4753\ : std_logic;
signal \N__4750\ : std_logic;
signal \N__4747\ : std_logic;
signal \N__4744\ : std_logic;
signal \N__4741\ : std_logic;
signal \N__4738\ : std_logic;
signal \N__4735\ : std_logic;
signal \N__4732\ : std_logic;
signal \N__4729\ : std_logic;
signal \N__4726\ : std_logic;
signal \N__4723\ : std_logic;
signal \N__4720\ : std_logic;
signal \N__4717\ : std_logic;
signal \N__4714\ : std_logic;
signal \N__4711\ : std_logic;
signal \N__4708\ : std_logic;
signal \N__4705\ : std_logic;
signal \N__4702\ : std_logic;
signal \N__4699\ : std_logic;
signal \N__4696\ : std_logic;
signal \N__4693\ : std_logic;
signal \N__4690\ : std_logic;
signal \N__4687\ : std_logic;
signal \N__4684\ : std_logic;
signal \N__4681\ : std_logic;
signal \N__4678\ : std_logic;
signal \N__4675\ : std_logic;
signal \N__4672\ : std_logic;
signal \N__4669\ : std_logic;
signal \N__4666\ : std_logic;
signal \N__4663\ : std_logic;
signal \N__4660\ : std_logic;
signal \N__4657\ : std_logic;
signal \N__4654\ : std_logic;
signal \N__4651\ : std_logic;
signal \N__4648\ : std_logic;
signal \N__4645\ : std_logic;
signal \N__4642\ : std_logic;
signal \N__4639\ : std_logic;
signal \N__4636\ : std_logic;
signal \N__4633\ : std_logic;
signal \N__4630\ : std_logic;
signal \N__4627\ : std_logic;
signal \N__4624\ : std_logic;
signal \N__4621\ : std_logic;
signal \N__4618\ : std_logic;
signal \N__4615\ : std_logic;
signal \N__4612\ : std_logic;
signal \N__4609\ : std_logic;
signal \N__4606\ : std_logic;
signal \N__4601\ : std_logic;
signal \N__4598\ : std_logic;
signal \N__4595\ : std_logic;
signal \N__4592\ : std_logic;
signal \N__4589\ : std_logic;
signal \N__4586\ : std_logic;
signal \N__4585\ : std_logic;
signal \N__4582\ : std_logic;
signal \N__4579\ : std_logic;
signal \N__4576\ : std_logic;
signal \N__4573\ : std_logic;
signal \N__4570\ : std_logic;
signal \N__4567\ : std_logic;
signal \N__4564\ : std_logic;
signal \N__4561\ : std_logic;
signal \N__4558\ : std_logic;
signal \N__4555\ : std_logic;
signal \N__4552\ : std_logic;
signal \N__4549\ : std_logic;
signal \N__4546\ : std_logic;
signal \N__4543\ : std_logic;
signal \N__4540\ : std_logic;
signal \N__4537\ : std_logic;
signal \N__4534\ : std_logic;
signal \N__4531\ : std_logic;
signal \N__4528\ : std_logic;
signal \N__4525\ : std_logic;
signal \N__4522\ : std_logic;
signal \N__4519\ : std_logic;
signal \N__4516\ : std_logic;
signal \N__4513\ : std_logic;
signal \N__4510\ : std_logic;
signal \N__4507\ : std_logic;
signal \N__4504\ : std_logic;
signal \N__4501\ : std_logic;
signal \N__4498\ : std_logic;
signal \N__4495\ : std_logic;
signal \N__4492\ : std_logic;
signal \N__4489\ : std_logic;
signal \N__4486\ : std_logic;
signal \N__4483\ : std_logic;
signal \N__4480\ : std_logic;
signal \N__4477\ : std_logic;
signal \N__4474\ : std_logic;
signal \N__4471\ : std_logic;
signal \N__4468\ : std_logic;
signal \N__4465\ : std_logic;
signal \N__4462\ : std_logic;
signal \N__4459\ : std_logic;
signal \N__4456\ : std_logic;
signal \N__4453\ : std_logic;
signal \N__4450\ : std_logic;
signal \N__4447\ : std_logic;
signal \N__4444\ : std_logic;
signal \N__4441\ : std_logic;
signal \N__4438\ : std_logic;
signal \N__4435\ : std_logic;
signal \N__4432\ : std_logic;
signal \N__4429\ : std_logic;
signal \N__4426\ : std_logic;
signal \N__4423\ : std_logic;
signal \N__4420\ : std_logic;
signal \N__4417\ : std_logic;
signal \N__4414\ : std_logic;
signal \N__4411\ : std_logic;
signal \N__4408\ : std_logic;
signal \N__4405\ : std_logic;
signal \N__4402\ : std_logic;
signal \N__4399\ : std_logic;
signal \N__4396\ : std_logic;
signal \N__4393\ : std_logic;
signal \N__4390\ : std_logic;
signal \N__4387\ : std_logic;
signal \N__4382\ : std_logic;
signal \N__4379\ : std_logic;
signal \N__4376\ : std_logic;
signal \N__4373\ : std_logic;
signal \N__4372\ : std_logic;
signal \N__4369\ : std_logic;
signal \N__4368\ : std_logic;
signal \N__4365\ : std_logic;
signal \N__4362\ : std_logic;
signal \N__4359\ : std_logic;
signal \N__4356\ : std_logic;
signal \N__4355\ : std_logic;
signal \N__4350\ : std_logic;
signal \N__4349\ : std_logic;
signal \N__4346\ : std_logic;
signal \N__4343\ : std_logic;
signal \N__4340\ : std_logic;
signal \N__4337\ : std_logic;
signal \N__4334\ : std_logic;
signal \N__4331\ : std_logic;
signal \N__4330\ : std_logic;
signal \N__4325\ : std_logic;
signal \N__4324\ : std_logic;
signal \N__4319\ : std_logic;
signal \N__4316\ : std_logic;
signal \N__4313\ : std_logic;
signal \N__4310\ : std_logic;
signal \N__4307\ : std_logic;
signal \N__4304\ : std_logic;
signal \N__4303\ : std_logic;
signal \N__4298\ : std_logic;
signal \N__4293\ : std_logic;
signal \N__4290\ : std_logic;
signal \N__4287\ : std_logic;
signal \N__4284\ : std_logic;
signal \N__4281\ : std_logic;
signal \N__4278\ : std_logic;
signal \N__4273\ : std_logic;
signal \N__4270\ : std_logic;
signal \N__4267\ : std_logic;
signal \N__4262\ : std_logic;
signal \N__4261\ : std_logic;
signal \N__4258\ : std_logic;
signal \N__4255\ : std_logic;
signal \N__4252\ : std_logic;
signal \N__4251\ : std_logic;
signal \N__4248\ : std_logic;
signal \N__4247\ : std_logic;
signal \N__4244\ : std_logic;
signal \N__4241\ : std_logic;
signal \N__4240\ : std_logic;
signal \N__4237\ : std_logic;
signal \N__4234\ : std_logic;
signal \N__4229\ : std_logic;
signal \N__4228\ : std_logic;
signal \N__4225\ : std_logic;
signal \N__4220\ : std_logic;
signal \N__4219\ : std_logic;
signal \N__4216\ : std_logic;
signal \N__4213\ : std_logic;
signal \N__4210\ : std_logic;
signal \N__4207\ : std_logic;
signal \N__4204\ : std_logic;
signal \N__4199\ : std_logic;
signal \N__4196\ : std_logic;
signal \N__4191\ : std_logic;
signal \N__4190\ : std_logic;
signal \N__4185\ : std_logic;
signal \N__4182\ : std_logic;
signal \N__4179\ : std_logic;
signal \N__4176\ : std_logic;
signal \N__4171\ : std_logic;
signal \N__4168\ : std_logic;
signal \N__4165\ : std_logic;
signal \N__4162\ : std_logic;
signal \N__4159\ : std_logic;
signal \N__4154\ : std_logic;
signal \N__4151\ : std_logic;
signal \N__4148\ : std_logic;
signal \N__4147\ : std_logic;
signal \N__4146\ : std_logic;
signal \N__4145\ : std_logic;
signal \N__4144\ : std_logic;
signal \N__4141\ : std_logic;
signal \N__4138\ : std_logic;
signal \N__4135\ : std_logic;
signal \N__4132\ : std_logic;
signal \N__4131\ : std_logic;
signal \N__4128\ : std_logic;
signal \N__4123\ : std_logic;
signal \N__4122\ : std_logic;
signal \N__4119\ : std_logic;
signal \N__4116\ : std_logic;
signal \N__4113\ : std_logic;
signal \N__4110\ : std_logic;
signal \N__4107\ : std_logic;
signal \N__4104\ : std_logic;
signal \N__4103\ : std_logic;
signal \N__4100\ : std_logic;
signal \N__4095\ : std_logic;
signal \N__4092\ : std_logic;
signal \N__4087\ : std_logic;
signal \N__4084\ : std_logic;
signal \N__4081\ : std_logic;
signal \N__4076\ : std_logic;
signal \N__4073\ : std_logic;
signal \N__4070\ : std_logic;
signal \N__4067\ : std_logic;
signal \N__4064\ : std_logic;
signal \N__4059\ : std_logic;
signal \N__4054\ : std_logic;
signal \N__4051\ : std_logic;
signal \N__4046\ : std_logic;
signal \N__4043\ : std_logic;
signal \N__4040\ : std_logic;
signal \N__4039\ : std_logic;
signal \N__4036\ : std_logic;
signal \N__4033\ : std_logic;
signal \N__4028\ : std_logic;
signal \N__4027\ : std_logic;
signal \N__4024\ : std_logic;
signal \N__4021\ : std_logic;
signal \N__4016\ : std_logic;
signal \N__4015\ : std_logic;
signal \N__4014\ : std_logic;
signal \N__4011\ : std_logic;
signal \N__4008\ : std_logic;
signal \N__4007\ : std_logic;
signal \N__4004\ : std_logic;
signal \N__3999\ : std_logic;
signal \N__3998\ : std_logic;
signal \N__3995\ : std_logic;
signal \N__3992\ : std_logic;
signal \N__3989\ : std_logic;
signal \N__3986\ : std_logic;
signal \N__3983\ : std_logic;
signal \N__3982\ : std_logic;
signal \N__3979\ : std_logic;
signal \N__3976\ : std_logic;
signal \N__3973\ : std_logic;
signal \N__3970\ : std_logic;
signal \N__3967\ : std_logic;
signal \N__3964\ : std_logic;
signal \N__3961\ : std_logic;
signal \N__3958\ : std_logic;
signal \N__3953\ : std_logic;
signal \N__3950\ : std_logic;
signal \N__3947\ : std_logic;
signal \N__3944\ : std_logic;
signal \N__3941\ : std_logic;
signal \N__3932\ : std_logic;
signal \N__3929\ : std_logic;
signal \N__3926\ : std_logic;
signal \N__3925\ : std_logic;
signal \N__3922\ : std_logic;
signal \N__3919\ : std_logic;
signal \N__3914\ : std_logic;
signal \N__3913\ : std_logic;
signal \N__3910\ : std_logic;
signal \N__3907\ : std_logic;
signal \N__3906\ : std_logic;
signal \N__3901\ : std_logic;
signal \N__3898\ : std_logic;
signal \N__3895\ : std_logic;
signal \N__3892\ : std_logic;
signal \N__3891\ : std_logic;
signal \N__3890\ : std_logic;
signal \N__3885\ : std_logic;
signal \N__3882\ : std_logic;
signal \N__3881\ : std_logic;
signal \N__3878\ : std_logic;
signal \N__3875\ : std_logic;
signal \N__3872\ : std_logic;
signal \N__3869\ : std_logic;
signal \N__3868\ : std_logic;
signal \N__3865\ : std_logic;
signal \N__3862\ : std_logic;
signal \N__3857\ : std_logic;
signal \N__3854\ : std_logic;
signal \N__3851\ : std_logic;
signal \N__3844\ : std_logic;
signal \GNDG0\ : std_logic;
signal din_c_3 : std_logic;
signal din_c_2 : std_logic;
signal \VCCG0\ : std_logic;
signal din_c_6 : std_logic;
signal din_c_7 : std_logic;
signal din_c_4 : std_logic;
signal din_c_5 : std_logic;
signal raddr_c_5 : std_logic;
signal waddr_c_3 : std_logic;
signal waddr_c_6 : std_logic;
signal wclk_c_g : std_logic;
signal raddr_c_2 : std_logic;
signal raddr_c_7 : std_logic;
signal waddr_c_5 : std_logic;
signal din_c_1 : std_logic;
signal raddr_c_8 : std_logic;
signal waddr_c_4 : std_logic;
signal raddr_c_10 : std_logic;
signal raddr_c_4 : std_logic;
signal waddr_c_9 : std_logic;
signal raddr_c_9 : std_logic;
signal waddr_c_7 : std_logic;
signal raddr_c_0 : std_logic;
signal waddr_c_10 : std_logic;
signal waddr_c_8 : std_logic;
signal raddr_c_1 : std_logic;
signal raddr_c_6 : std_logic;
signal waddr_c_2 : std_logic;
signal din_c_0 : std_logic;
signal rclk_c_g : std_logic;
signal raddr_c_3 : std_logic;
signal waddr_c_1 : std_logic;
signal waddr_c_0 : std_logic;
signal \mem_WE_4\ : std_logic;
signal \mem_WE_0\ : std_logic;
signal \mem_WE_8\ : std_logic;
signal \mem_WE_12\ : std_logic;
signal \mem_WE_16\ : std_logic;
signal \mem_WE_20\ : std_logic;
signal \mem_WE_24\ : std_logic;
signal write_en_c : std_logic;
signal waddr_c_13 : std_logic;
signal waddr_c_11 : std_logic;
signal waddr_c_12 : std_logic;
signal \mem_WE_28\ : std_logic;
signal mem_out_bus0_0 : std_logic;
signal mem_out_bus4_0 : std_logic;
signal mem_out_bus0_1 : std_logic;
signal mem_out_bus4_1 : std_logic;
signal mem_out_bus4_7 : std_logic;
signal mem_out_bus0_7 : std_logic;
signal mem_out_bus0_6 : std_logic;
signal mem_out_bus4_6 : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal mem_out_bus5_1 : std_logic;
signal mem_out_bus1_1 : std_logic;
signal mem_out_bus5_0 : std_logic;
signal mem_out_bus1_0 : std_logic;
signal \dout_obuf_RNO_4Z0Z_1\ : std_logic;
signal \mem_N_162_cascade_\ : std_logic;
signal dout_c_1 : std_logic;
signal \dout_obuf_RNO_4Z0Z_0\ : std_logic;
signal \mem_N_156_cascade_\ : std_logic;
signal dout_c_0 : std_logic;
signal \dout_obuf_RNO_2Z0Z_1\ : std_logic;
signal \mem_N_160\ : std_logic;
signal \dout_obuf_RNO_2Z0Z_0\ : std_logic;
signal \mem_N_154\ : std_logic;
signal mem_out_bus5_2 : std_logic;
signal mem_out_bus1_2 : std_logic;
signal \dout_obuf_RNO_2Z0Z_2\ : std_logic;
signal \mem_N_166_cascade_\ : std_logic;
signal dout_c_2 : std_logic;
signal \dout_obuf_RNO_4Z0Z_7\ : std_logic;
signal mem_out_bus5_7 : std_logic;
signal mem_out_bus1_7 : std_logic;
signal \dout_obuf_RNO_2Z0Z_7_cascade_\ : std_logic;
signal \mem_N_150\ : std_logic;
signal \mem_N_149_cascade_\ : std_logic;
signal dout_c_7 : std_logic;
signal mem_out_bus2_1 : std_logic;
signal mem_out_bus6_1 : std_logic;
signal \dout_obuf_RNO_5Z0Z_1\ : std_logic;
signal mem_out_bus6_0 : std_logic;
signal mem_out_bus2_0 : std_logic;
signal \dout_obuf_RNO_5Z0Z_0\ : std_logic;
signal mem_out_bus6_3 : std_logic;
signal mem_out_bus2_3 : std_logic;
signal mem_out_bus7_0 : std_logic;
signal mem_out_bus3_0 : std_logic;
signal \dout_obuf_RNO_3Z0Z_0\ : std_logic;
signal mem_out_bus7_2 : std_logic;
signal mem_out_bus3_2 : std_logic;
signal \dout_obuf_RNO_3Z0Z_2\ : std_logic;
signal mem_out_bus7_3 : std_logic;
signal mem_out_bus3_3 : std_logic;
signal mem_out_bus4_2 : std_logic;
signal mem_out_bus0_2 : std_logic;
signal mem_out_bus4_3 : std_logic;
signal mem_out_bus0_3 : std_logic;
signal mem_out_bus4_5 : std_logic;
signal mem_out_bus0_5 : std_logic;
signal mem_out_bus0_4 : std_logic;
signal mem_out_bus4_4 : std_logic;
signal \dout_obuf_RNO_4Z0Z_4\ : std_logic;
signal \mem_N_180_cascade_\ : std_logic;
signal dout_c_4 : std_logic;
signal \dout_obuf_RNO_4Z0Z_6\ : std_logic;
signal \mem_N_145_cascade_\ : std_logic;
signal dout_c_6 : std_logic;
signal \dout_obuf_RNO_4Z0Z_3\ : std_logic;
signal \dout_obuf_RNO_5Z0Z_3\ : std_logic;
signal mem_out_bus5_3 : std_logic;
signal mem_out_bus1_3 : std_logic;
signal \dout_obuf_RNO_3Z0Z_3\ : std_logic;
signal \dout_obuf_RNO_2Z0Z_3_cascade_\ : std_logic;
signal \mem_N_174\ : std_logic;
signal \mem_N_172_cascade_\ : std_logic;
signal dout_c_3 : std_logic;
signal \dout_obuf_RNO_4Z0Z_2\ : std_logic;
signal \mem_N_168\ : std_logic;
signal mem_out_bus1_4 : std_logic;
signal mem_out_bus5_4 : std_logic;
signal \dout_obuf_RNO_2Z0Z_4_cascade_\ : std_logic;
signal \mem_N_178\ : std_logic;
signal mem_out_bus1_6 : std_logic;
signal mem_out_bus5_6 : std_logic;
signal \dout_obuf_RNO_2Z0Z_6_cascade_\ : std_logic;
signal \mem_N_144\ : std_logic;
signal mem_out_bus6_4 : std_logic;
signal mem_out_bus2_4 : std_logic;
signal \dout_obuf_RNO_5Z0Z_4\ : std_logic;
signal mem_out_bus2_2 : std_logic;
signal mem_out_bus6_2 : std_logic;
signal \dout_obuf_RNO_5Z0Z_2\ : std_logic;
signal mem_out_bus6_6 : std_logic;
signal mem_out_bus2_6 : std_logic;
signal \dout_obuf_RNO_5Z0Z_6\ : std_logic;
signal mem_out_bus6_7 : std_logic;
signal mem_out_bus2_7 : std_logic;
signal \dout_obuf_RNO_5Z0Z_7\ : std_logic;
signal mem_out_bus7_1 : std_logic;
signal mem_out_bus3_1 : std_logic;
signal \dout_obuf_RNO_3Z0Z_1\ : std_logic;
signal mem_out_bus7_4 : std_logic;
signal mem_out_bus3_4 : std_logic;
signal \dout_obuf_RNO_3Z0Z_4\ : std_logic;
signal mem_out_bus7_7 : std_logic;
signal mem_out_bus3_7 : std_logic;
signal \dout_obuf_RNO_3Z0Z_7\ : std_logic;
signal mem_out_bus7_6 : std_logic;
signal mem_out_bus3_6 : std_logic;
signal \dout_obuf_RNO_3Z0Z_6\ : std_logic;
signal \dout_obuf_RNO_4Z0Z_5\ : std_logic;
signal mem_out_bus1_5 : std_logic;
signal mem_out_bus5_5 : std_logic;
signal \mem_radregZ0Z_12\ : std_logic;
signal \dout_obuf_RNO_2Z0Z_5_cascade_\ : std_logic;
signal \mem_N_140\ : std_logic;
signal \mem_radregZ0Z_11\ : std_logic;
signal \mem_N_139\ : std_logic;
signal dout_c_5 : std_logic;
signal mem_out_bus6_5 : std_logic;
signal mem_out_bus2_5 : std_logic;
signal \dout_obuf_RNO_5Z0Z_5\ : std_logic;
signal \mem_radregZ0Z_13\ : std_logic;
signal mem_out_bus7_5 : std_logic;
signal mem_out_bus3_5 : std_logic;
signal \dout_obuf_RNO_3Z0Z_5\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal wclk_wire : std_logic;
signal rclk_wire : std_logic;
signal waddr_wire : std_logic_vector(13 downto 0);
signal dout_wire : std_logic_vector(7 downto 0);
signal raddr_wire : std_logic_vector(13 downto 0);
signal din_wire : std_logic_vector(7 downto 0);
signal write_en_wire : std_logic;
signal \mem_mem_3_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_3_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_3_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_3_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_3_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_5_2_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_5_2_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_5_2_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_5_2_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_5_2_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_2_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_2_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_2_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_2_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_2_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_1_3_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_1_3_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_1_3_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_1_3_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_1_3_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_4_2_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_4_2_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_4_2_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_4_2_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_4_2_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_7_2_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_7_2_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_7_2_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_7_2_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_7_2_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_3_3_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_3_3_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_3_3_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_3_3_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_3_3_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_6_2_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_6_2_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_6_2_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_6_2_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_6_2_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_5_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_5_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_5_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_5_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_5_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_2_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_2_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_2_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_2_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_2_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_1_2_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_1_2_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_1_2_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_1_2_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_1_2_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_4_3_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_4_3_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_4_3_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_4_3_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_4_3_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_0_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_0_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_0_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_0_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_0_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_3_2_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_3_2_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_3_2_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_3_2_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_3_2_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_6_3_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_6_3_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_6_3_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_6_3_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_6_3_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_5_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_5_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_5_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_5_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_5_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_2_2_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_2_2_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_2_2_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_2_2_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_2_2_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_7_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_7_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_7_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_7_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_7_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_1_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_1_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_1_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_1_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_1_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_4_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_4_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_4_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_4_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_4_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_2_3_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_2_3_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_2_3_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_2_3_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_2_3_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_7_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_7_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_7_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_7_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_7_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_1_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_1_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_1_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_1_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_1_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_4_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_4_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_4_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_4_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_4_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_0_2_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_0_2_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_0_2_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_0_2_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_0_2_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_3_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_3_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_3_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_3_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_3_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_6_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_6_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_6_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_6_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_6_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_5_3_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_5_3_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_5_3_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_5_3_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_5_3_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_7_3_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_7_3_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_7_3_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_7_3_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_7_3_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_0_3_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_0_3_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_0_3_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_0_3_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_0_3_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_6_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_6_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_6_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \mem_mem_6_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \mem_mem_6_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    wclk_wire <= wclk;
    rclk_wire <= rclk;
    waddr_wire <= waddr;
    dout <= dout_wire;
    raddr_wire <= raddr;
    din_wire <= din;
    write_en_wire <= write_en;
    mem_out_bus3_1 <= \mem_mem_3_0_physical_RDATA_wire\(11);
    mem_out_bus3_0 <= \mem_mem_3_0_physical_RDATA_wire\(3);
    \mem_mem_3_0_physical_RADDR_wire\ <= \N__7339\&\N__6676\&\N__7774\&\N__8308\&\N__5356\&\N__9289\&\N__7114\&\N__4693\&\N__8533\&\N__5584\&\N__6244\;
    \mem_mem_3_0_physical_WADDR_wire\ <= \N__6028\&\N__6892\&\N__5806\&\N__6460\&\N__8857\&\N__8101\&\N__7558\&\N__9070\&\N__5140\&\N__4468\&\N__9685\;
    \mem_mem_3_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \mem_mem_3_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8012\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__4991\&'0'&'0'&'0';
    mem_out_bus5_5 <= \mem_mem_5_2_physical_RDATA_wire\(11);
    mem_out_bus5_4 <= \mem_mem_5_2_physical_RDATA_wire\(3);
    \mem_mem_5_2_physical_RADDR_wire\ <= \N__7390\&\N__6727\&\N__7831\&\N__8365\&\N__5419\&\N__9340\&\N__7177\&\N__4738\&\N__8590\&\N__5647\&\N__6295\;
    \mem_mem_5_2_physical_WADDR_wire\ <= \N__6073\&\N__6943\&\N__5857\&\N__6511\&\N__8896\&\N__8140\&\N__7609\&\N__9121\&\N__5185\&\N__4513\&\N__9742\;
    \mem_mem_5_2_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \mem_mem_5_2_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__9524\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__4368\&'0'&'0'&'0';
    mem_out_bus2_1 <= \mem_mem_2_0_physical_RDATA_wire\(11);
    mem_out_bus2_0 <= \mem_mem_2_0_physical_RDATA_wire\(3);
    \mem_mem_2_0_physical_RADDR_wire\ <= \N__7387\&\N__6724\&\N__7822\&\N__8356\&\N__5404\&\N__9337\&\N__7162\&\N__4741\&\N__8581\&\N__5632\&\N__6292\;
    \mem_mem_2_0_physical_WADDR_wire\ <= \N__6076\&\N__6940\&\N__5854\&\N__6508\&\N__8905\&\N__8149\&\N__7606\&\N__9118\&\N__5188\&\N__4516\&\N__9733\;
    \mem_mem_2_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \mem_mem_2_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8004\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__5018\&'0'&'0'&'0';
    mem_out_bus1_7 <= \mem_mem_1_3_physical_RDATA_wire\(11);
    mem_out_bus1_6 <= \mem_mem_1_3_physical_RDATA_wire\(3);
    \mem_mem_1_3_physical_RADDR_wire\ <= \N__7399\&\N__6736\&\N__7834\&\N__8368\&\N__5416\&\N__9349\&\N__7174\&\N__4753\&\N__8593\&\N__5644\&\N__6304\;
    \mem_mem_1_3_physical_WADDR_wire\ <= \N__6088\&\N__6952\&\N__5866\&\N__6520\&\N__8917\&\N__8161\&\N__7618\&\N__9130\&\N__5200\&\N__4528\&\N__9745\;
    \mem_mem_1_3_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \mem_mem_1_3_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__4147\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__4247\&'0'&'0'&'0';
    mem_out_bus4_5 <= \mem_mem_4_2_physical_RDATA_wire\(11);
    mem_out_bus4_4 <= \mem_mem_4_2_physical_RDATA_wire\(3);
    \mem_mem_4_2_physical_RADDR_wire\ <= \N__7438\&\N__6775\&\N__7879\&\N__8413\&\N__5467\&\N__9388\&\N__7225\&\N__4786\&\N__8638\&\N__5695\&\N__6343\;
    \mem_mem_4_2_physical_WADDR_wire\ <= \N__6121\&\N__6991\&\N__5905\&\N__6559\&\N__8944\&\N__8188\&\N__7657\&\N__9169\&\N__5233\&\N__4561\&\N__9790\;
    \mem_mem_4_2_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \mem_mem_4_2_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__9522\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__4376\&'0'&'0'&'0';
    mem_out_bus7_5 <= \mem_mem_7_2_physical_RDATA_wire\(11);
    mem_out_bus7_4 <= \mem_mem_7_2_physical_RDATA_wire\(3);
    \mem_mem_7_2_physical_RADDR_wire\ <= \N__7294\&\N__6631\&\N__7735\&\N__8269\&\N__5323\&\N__9244\&\N__7081\&\N__4642\&\N__8494\&\N__5551\&\N__6199\;
    \mem_mem_7_2_physical_WADDR_wire\ <= \N__5977\&\N__6847\&\N__5761\&\N__6415\&\N__8800\&\N__8044\&\N__7513\&\N__9025\&\N__5089\&\N__4417\&\N__9646\;
    \mem_mem_7_2_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \mem_mem_7_2_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__9523\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__4324\&'0'&'0'&'0';
    mem_out_bus0_1 <= \mem_mem_0_0_physical_RDATA_wire\(11);
    mem_out_bus0_0 <= \mem_mem_0_0_physical_RDATA_wire\(3);
    \mem_mem_0_0_physical_RADDR_wire\ <= \N__7472\&\N__6809\&\N__7910\&\N__8444\&\N__5495\&\N__9422\&\N__7253\&\N__4823\&\N__8669\&\N__5723\&\N__6377\;
    \mem_mem_0_0_physical_WADDR_wire\ <= \N__6158\&\N__7025\&\N__5939\&\N__6593\&\N__8984\&\N__8228\&\N__7691\&\N__9203\&\N__5270\&\N__4598\&\N__9821\;
    \mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \mem_mem_0_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8014\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__5051\&'0'&'0'&'0';
    mem_out_bus3_7 <= \mem_mem_3_3_physical_RDATA_wire\(11);
    mem_out_bus3_6 <= \mem_mem_3_3_physical_RDATA_wire\(3);
    \mem_mem_3_3_physical_RADDR_wire\ <= \N__7303\&\N__6640\&\N__7738\&\N__8272\&\N__5320\&\N__9253\&\N__7078\&\N__4657\&\N__8497\&\N__5548\&\N__6208\;
    \mem_mem_3_3_physical_WADDR_wire\ <= \N__5992\&\N__6856\&\N__5770\&\N__6424\&\N__8821\&\N__8065\&\N__7522\&\N__9034\&\N__5104\&\N__4432\&\N__9649\;
    \mem_mem_3_3_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \mem_mem_3_3_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__4103\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__4190\&'0'&'0'&'0';
    mem_out_bus6_5 <= \mem_mem_6_2_physical_RDATA_wire\(11);
    mem_out_bus6_4 <= \mem_mem_6_2_physical_RDATA_wire\(3);
    \mem_mem_6_2_physical_RADDR_wire\ <= \N__7342\&\N__6679\&\N__7783\&\N__8317\&\N__5371\&\N__9292\&\N__7129\&\N__4690\&\N__8542\&\N__5599\&\N__6247\;
    \mem_mem_6_2_physical_WADDR_wire\ <= \N__6025\&\N__6895\&\N__5809\&\N__6463\&\N__8848\&\N__8092\&\N__7561\&\N__9073\&\N__5137\&\N__4465\&\N__9694\;
    \mem_mem_6_2_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \mem_mem_6_2_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__9516\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__4349\&'0'&'0'&'0';
    mem_out_bus5_3 <= \mem_mem_5_1_physical_RDATA_wire\(11);
    mem_out_bus5_2 <= \mem_mem_5_1_physical_RDATA_wire\(3);
    \mem_mem_5_1_physical_RADDR_wire\ <= \N__7402\&\N__6739\&\N__7843\&\N__8377\&\N__5431\&\N__9352\&\N__7189\&\N__4750\&\N__8602\&\N__5659\&\N__6307\;
    \mem_mem_5_1_physical_WADDR_wire\ <= \N__6085\&\N__6955\&\N__5869\&\N__6523\&\N__8908\&\N__8152\&\N__7621\&\N__9133\&\N__5197\&\N__4525\&\N__9754\;
    \mem_mem_5_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \mem_mem_5_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__4039\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__3925\&'0'&'0'&'0';
    mem_out_bus2_3 <= \mem_mem_2_1_physical_RDATA_wire\(11);
    mem_out_bus2_2 <= \mem_mem_2_1_physical_RDATA_wire\(3);
    \mem_mem_2_1_physical_RADDR_wire\ <= \N__7375\&\N__6712\&\N__7810\&\N__8344\&\N__5392\&\N__9325\&\N__7150\&\N__4729\&\N__8569\&\N__5620\&\N__6280\;
    \mem_mem_2_1_physical_WADDR_wire\ <= \N__6064\&\N__6928\&\N__5842\&\N__6496\&\N__8893\&\N__8137\&\N__7594\&\N__9106\&\N__5176\&\N__4504\&\N__9721\;
    \mem_mem_2_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \mem_mem_2_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__4007\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__3881\&'0'&'0'&'0';
    mem_out_bus1_5 <= \mem_mem_1_2_physical_RDATA_wire\(11);
    mem_out_bus1_4 <= \mem_mem_1_2_physical_RDATA_wire\(3);
    \mem_mem_1_2_physical_RADDR_wire\ <= \N__7411\&\N__6748\&\N__7846\&\N__8380\&\N__5428\&\N__9361\&\N__7186\&\N__4765\&\N__8605\&\N__5656\&\N__6316\;
    \mem_mem_1_2_physical_WADDR_wire\ <= \N__6100\&\N__6964\&\N__5878\&\N__6532\&\N__8929\&\N__8173\&\N__7630\&\N__9142\&\N__5212\&\N__4540\&\N__9757\;
    \mem_mem_1_2_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \mem_mem_1_2_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__9520\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__4355\&'0'&'0'&'0';
    mem_out_bus4_7 <= \mem_mem_4_3_physical_RDATA_wire\(11);
    mem_out_bus4_6 <= \mem_mem_4_3_physical_RDATA_wire\(3);
    \mem_mem_4_3_physical_RADDR_wire\ <= \N__7426\&\N__6763\&\N__7867\&\N__8401\&\N__5455\&\N__9376\&\N__7213\&\N__4774\&\N__8626\&\N__5683\&\N__6331\;
    \mem_mem_4_3_physical_WADDR_wire\ <= \N__6109\&\N__6979\&\N__5893\&\N__6547\&\N__8932\&\N__8176\&\N__7645\&\N__9157\&\N__5221\&\N__4549\&\N__9778\;
    \mem_mem_4_3_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \mem_mem_4_3_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__4146\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__4262\&'0'&'0'&'0';
    mem_out_bus0_3 <= \mem_mem_0_1_physical_RDATA_wire\(11);
    mem_out_bus0_2 <= \mem_mem_0_1_physical_RDATA_wire\(3);
    \mem_mem_0_1_physical_RADDR_wire\ <= \N__7466\&\N__6803\&\N__7904\&\N__8438\&\N__5488\&\N__9416\&\N__7246\&\N__4817\&\N__8663\&\N__5716\&\N__6371\;
    \mem_mem_0_1_physical_WADDR_wire\ <= \N__6152\&\N__7019\&\N__5933\&\N__6587\&\N__8978\&\N__8222\&\N__7685\&\N__9197\&\N__5264\&\N__4592\&\N__9815\;
    \mem_mem_0_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \mem_mem_0_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__4014\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__3891\&'0'&'0'&'0';
    mem_out_bus3_5 <= \mem_mem_3_2_physical_RDATA_wire\(11);
    mem_out_bus3_4 <= \mem_mem_3_2_physical_RDATA_wire\(3);
    \mem_mem_3_2_physical_RADDR_wire\ <= \N__7315\&\N__6652\&\N__7750\&\N__8284\&\N__5332\&\N__9265\&\N__7090\&\N__4669\&\N__8509\&\N__5560\&\N__6220\;
    \mem_mem_3_2_physical_WADDR_wire\ <= \N__6004\&\N__6868\&\N__5782\&\N__6436\&\N__8833\&\N__8077\&\N__7534\&\N__9046\&\N__5116\&\N__4444\&\N__9661\;
    \mem_mem_3_2_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \mem_mem_3_2_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__9487\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__4303\&'0'&'0'&'0';
    mem_out_bus6_7 <= \mem_mem_6_3_physical_RDATA_wire\(11);
    mem_out_bus6_6 <= \mem_mem_6_3_physical_RDATA_wire\(3);
    \mem_mem_6_3_physical_RADDR_wire\ <= \N__7330\&\N__6667\&\N__7771\&\N__8305\&\N__5359\&\N__9280\&\N__7117\&\N__4678\&\N__8530\&\N__5587\&\N__6235\;
    \mem_mem_6_3_physical_WADDR_wire\ <= \N__6013\&\N__6883\&\N__5797\&\N__6451\&\N__8836\&\N__8080\&\N__7549\&\N__9061\&\N__5125\&\N__4453\&\N__9682\;
    \mem_mem_6_3_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \mem_mem_6_3_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__4131\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__4228\&'0'&'0'&'0';
    mem_out_bus5_1 <= \mem_mem_5_0_physical_RDATA_wire\(11);
    mem_out_bus5_0 <= \mem_mem_5_0_physical_RDATA_wire\(3);
    \mem_mem_5_0_physical_RADDR_wire\ <= \N__7414\&\N__6751\&\N__7855\&\N__8389\&\N__5443\&\N__9364\&\N__7201\&\N__4762\&\N__8614\&\N__5671\&\N__6319\;
    \mem_mem_5_0_physical_WADDR_wire\ <= \N__6097\&\N__6967\&\N__5881\&\N__6535\&\N__8920\&\N__8164\&\N__7633\&\N__9145\&\N__5209\&\N__4537\&\N__9766\;
    \mem_mem_5_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \mem_mem_5_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8003\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__5036\&'0'&'0'&'0';
    mem_out_bus2_5 <= \mem_mem_2_2_physical_RDATA_wire\(11);
    mem_out_bus2_4 <= \mem_mem_2_2_physical_RDATA_wire\(3);
    \mem_mem_2_2_physical_RADDR_wire\ <= \N__7363\&\N__6700\&\N__7798\&\N__8332\&\N__5380\&\N__9313\&\N__7138\&\N__4717\&\N__8557\&\N__5608\&\N__6268\;
    \mem_mem_2_2_physical_WADDR_wire\ <= \N__6052\&\N__6916\&\N__5830\&\N__6484\&\N__8881\&\N__8125\&\N__7582\&\N__9094\&\N__5164\&\N__4492\&\N__9709\;
    \mem_mem_2_2_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \mem_mem_2_2_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__9497\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__4330\&'0'&'0'&'0';
    mem_out_bus7_3 <= \mem_mem_7_1_physical_RDATA_wire\(11);
    mem_out_bus7_2 <= \mem_mem_7_1_physical_RDATA_wire\(3);
    \mem_mem_7_1_physical_RADDR_wire\ <= \N__7306\&\N__6643\&\N__7747\&\N__8281\&\N__5335\&\N__9256\&\N__7093\&\N__4654\&\N__8506\&\N__5563\&\N__6211\;
    \mem_mem_7_1_physical_WADDR_wire\ <= \N__5989\&\N__6859\&\N__5773\&\N__6427\&\N__8812\&\N__8056\&\N__7525\&\N__9037\&\N__5101\&\N__4429\&\N__9658\;
    \mem_mem_7_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \mem_mem_7_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__4015\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__3906\&'0'&'0'&'0';
    mem_out_bus1_3 <= \mem_mem_1_1_physical_RDATA_wire\(11);
    mem_out_bus1_2 <= \mem_mem_1_1_physical_RDATA_wire\(3);
    \mem_mem_1_1_physical_RADDR_wire\ <= \N__7423\&\N__6760\&\N__7858\&\N__8392\&\N__5440\&\N__9373\&\N__7198\&\N__4777\&\N__8617\&\N__5668\&\N__6328\;
    \mem_mem_1_1_physical_WADDR_wire\ <= \N__6112\&\N__6976\&\N__5890\&\N__6544\&\N__8941\&\N__8185\&\N__7642\&\N__9154\&\N__5224\&\N__4552\&\N__9769\;
    \mem_mem_1_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \mem_mem_1_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__3998\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__3890\&'0'&'0'&'0';
    mem_out_bus4_1 <= \mem_mem_4_0_physical_RDATA_wire\(11);
    mem_out_bus4_0 <= \mem_mem_4_0_physical_RDATA_wire\(3);
    \mem_mem_4_0_physical_RADDR_wire\ <= \N__7462\&\N__6799\&\N__7903\&\N__8437\&\N__5491\&\N__9412\&\N__7249\&\N__4810\&\N__8662\&\N__5719\&\N__6367\;
    \mem_mem_4_0_physical_WADDR_wire\ <= \N__6145\&\N__7015\&\N__5929\&\N__6583\&\N__8968\&\N__8212\&\N__7681\&\N__9193\&\N__5257\&\N__4585\&\N__9814\;
    \mem_mem_4_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \mem_mem_4_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8015\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__5050\&'0'&'0'&'0';
    mem_out_bus2_7 <= \mem_mem_2_3_physical_RDATA_wire\(11);
    mem_out_bus2_6 <= \mem_mem_2_3_physical_RDATA_wire\(3);
    \mem_mem_2_3_physical_RADDR_wire\ <= \N__7351\&\N__6688\&\N__7786\&\N__8320\&\N__5368\&\N__9301\&\N__7126\&\N__4705\&\N__8545\&\N__5596\&\N__6256\;
    \mem_mem_2_3_physical_WADDR_wire\ <= \N__6040\&\N__6904\&\N__5818\&\N__6472\&\N__8869\&\N__8113\&\N__7570\&\N__9082\&\N__5152\&\N__4480\&\N__9697\;
    \mem_mem_2_3_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \mem_mem_2_3_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__4122\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__4219\&'0'&'0'&'0';
    mem_out_bus7_1 <= \mem_mem_7_0_physical_RDATA_wire\(11);
    mem_out_bus7_0 <= \mem_mem_7_0_physical_RDATA_wire\(3);
    \mem_mem_7_0_physical_RADDR_wire\ <= \N__7318\&\N__6655\&\N__7759\&\N__8293\&\N__5347\&\N__9268\&\N__7105\&\N__4666\&\N__8518\&\N__5575\&\N__6223\;
    \mem_mem_7_0_physical_WADDR_wire\ <= \N__6001\&\N__6871\&\N__5785\&\N__6439\&\N__8824\&\N__8068\&\N__7537\&\N__9049\&\N__5113\&\N__4441\&\N__9670\;
    \mem_mem_7_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \mem_mem_7_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8013\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__4984\&'0'&'0'&'0';
    mem_out_bus1_1 <= \mem_mem_1_0_physical_RDATA_wire\(11);
    mem_out_bus1_0 <= \mem_mem_1_0_physical_RDATA_wire\(3);
    \mem_mem_1_0_physical_RADDR_wire\ <= \N__7435\&\N__6772\&\N__7870\&\N__8404\&\N__5452\&\N__9385\&\N__7210\&\N__4789\&\N__8629\&\N__5680\&\N__6340\;
    \mem_mem_1_0_physical_WADDR_wire\ <= \N__6124\&\N__6988\&\N__5902\&\N__6556\&\N__8953\&\N__8197\&\N__7654\&\N__9166\&\N__5236\&\N__4564\&\N__9781\;
    \mem_mem_1_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \mem_mem_1_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8002\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__5040\&'0'&'0'&'0';
    mem_out_bus4_3 <= \mem_mem_4_1_physical_RDATA_wire\(11);
    mem_out_bus4_2 <= \mem_mem_4_1_physical_RDATA_wire\(3);
    \mem_mem_4_1_physical_RADDR_wire\ <= \N__7450\&\N__6787\&\N__7891\&\N__8425\&\N__5479\&\N__9400\&\N__7237\&\N__4798\&\N__8650\&\N__5707\&\N__6355\;
    \mem_mem_4_1_physical_WADDR_wire\ <= \N__6133\&\N__7003\&\N__5917\&\N__6571\&\N__8956\&\N__8200\&\N__7669\&\N__9181\&\N__5245\&\N__4573\&\N__9802\;
    \mem_mem_4_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \mem_mem_4_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__4046\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__3932\&'0'&'0'&'0';
    mem_out_bus0_5 <= \mem_mem_0_2_physical_RDATA_wire\(11);
    mem_out_bus0_4 <= \mem_mem_0_2_physical_RDATA_wire\(3);
    \mem_mem_0_2_physical_RADDR_wire\ <= \N__7459\&\N__6796\&\N__7894\&\N__8428\&\N__5476\&\N__9409\&\N__7234\&\N__4811\&\N__8653\&\N__5704\&\N__6364\;
    \mem_mem_0_2_physical_WADDR_wire\ <= \N__6146\&\N__7012\&\N__5926\&\N__6580\&\N__8972\&\N__8216\&\N__7678\&\N__9190\&\N__5258\&\N__4586\&\N__9805\;
    \mem_mem_0_2_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \mem_mem_0_2_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__9521\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__4372\&'0'&'0'&'0';
    mem_out_bus3_3 <= \mem_mem_3_1_physical_RDATA_wire\(11);
    mem_out_bus3_2 <= \mem_mem_3_1_physical_RDATA_wire\(3);
    \mem_mem_3_1_physical_RADDR_wire\ <= \N__7327\&\N__6664\&\N__7762\&\N__8296\&\N__5344\&\N__9277\&\N__7102\&\N__4681\&\N__8521\&\N__5572\&\N__6232\;
    \mem_mem_3_1_physical_WADDR_wire\ <= \N__6016\&\N__6880\&\N__5794\&\N__6448\&\N__8845\&\N__8089\&\N__7546\&\N__9058\&\N__5128\&\N__4456\&\N__9673\;
    \mem_mem_3_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \mem_mem_3_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__3982\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__3868\&'0'&'0'&'0';
    mem_out_bus6_1 <= \mem_mem_6_0_physical_RDATA_wire\(11);
    mem_out_bus6_0 <= \mem_mem_6_0_physical_RDATA_wire\(3);
    \mem_mem_6_0_physical_RADDR_wire\ <= \N__7366\&\N__6703\&\N__7807\&\N__8341\&\N__5395\&\N__9316\&\N__7153\&\N__4714\&\N__8566\&\N__5623\&\N__6271\;
    \mem_mem_6_0_physical_WADDR_wire\ <= \N__6049\&\N__6919\&\N__5833\&\N__6487\&\N__8872\&\N__8116\&\N__7585\&\N__9097\&\N__5161\&\N__4489\&\N__9718\;
    \mem_mem_6_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \mem_mem_6_0_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__8005\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__5011\&'0'&'0'&'0';
    mem_out_bus5_7 <= \mem_mem_5_3_physical_RDATA_wire\(11);
    mem_out_bus5_6 <= \mem_mem_5_3_physical_RDATA_wire\(3);
    \mem_mem_5_3_physical_RADDR_wire\ <= \N__7378\&\N__6715\&\N__7819\&\N__8353\&\N__5407\&\N__9328\&\N__7165\&\N__4726\&\N__8578\&\N__5635\&\N__6283\;
    \mem_mem_5_3_physical_WADDR_wire\ <= \N__6061\&\N__6931\&\N__5845\&\N__6499\&\N__8884\&\N__8128\&\N__7597\&\N__9109\&\N__5173\&\N__4501\&\N__9730\;
    \mem_mem_5_3_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \mem_mem_5_3_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__4145\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__4251\&'0'&'0'&'0';
    mem_out_bus7_7 <= \mem_mem_7_3_physical_RDATA_wire\(11);
    mem_out_bus7_6 <= \mem_mem_7_3_physical_RDATA_wire\(3);
    \mem_mem_7_3_physical_RADDR_wire\ <= \N__7282\&\N__6619\&\N__7723\&\N__8257\&\N__5311\&\N__9232\&\N__7069\&\N__4630\&\N__8482\&\N__5539\&\N__6187\;
    \mem_mem_7_3_physical_WADDR_wire\ <= \N__5965\&\N__6835\&\N__5749\&\N__6403\&\N__8788\&\N__8032\&\N__7501\&\N__9013\&\N__5077\&\N__4405\&\N__9634\;
    \mem_mem_7_3_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \mem_mem_7_3_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__4144\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__4240\&'0'&'0'&'0';
    mem_out_bus0_7 <= \mem_mem_0_3_physical_RDATA_wire\(11);
    mem_out_bus0_6 <= \mem_mem_0_3_physical_RDATA_wire\(3);
    \mem_mem_0_3_physical_RADDR_wire\ <= \N__7447\&\N__6784\&\N__7882\&\N__8416\&\N__5464\&\N__9397\&\N__7222\&\N__4801\&\N__8641\&\N__5692\&\N__6352\;
    \mem_mem_0_3_physical_WADDR_wire\ <= \N__6136\&\N__7000\&\N__5914\&\N__6568\&\N__8965\&\N__8209\&\N__7666\&\N__9178\&\N__5248\&\N__4576\&\N__9793\;
    \mem_mem_0_3_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \mem_mem_0_3_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__4154\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__4261\&'0'&'0'&'0';
    mem_out_bus6_3 <= \mem_mem_6_1_physical_RDATA_wire\(11);
    mem_out_bus6_2 <= \mem_mem_6_1_physical_RDATA_wire\(3);
    \mem_mem_6_1_physical_RADDR_wire\ <= \N__7354\&\N__6691\&\N__7795\&\N__8329\&\N__5383\&\N__9304\&\N__7141\&\N__4702\&\N__8554\&\N__5611\&\N__6259\;
    \mem_mem_6_1_physical_WADDR_wire\ <= \N__6037\&\N__6907\&\N__5821\&\N__6475\&\N__8860\&\N__8104\&\N__7573\&\N__9085\&\N__5149\&\N__4477\&\N__9706\;
    \mem_mem_6_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \mem_mem_6_1_physical_WDATA_wire\ <= '0'&'0'&'0'&'0'&\N__4027\&'0'&'0'&'0'&'0'&'0'&'0'&'0'&\N__3913\&'0'&'0'&'0';

    \mem_mem_3_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \mem_mem_3_0_physical_RDATA_wire\,
            RADDR => \mem_mem_3_0_physical_RADDR_wire\,
            WADDR => \mem_mem_3_0_physical_WADDR_wire\,
            MASK => \mem_mem_3_0_physical_MASK_wire\,
            WDATA => \mem_mem_3_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__4923\,
            RE => \N__10964\,
            WCLKE => \N__10238\,
            WCLK => \N__8764\,
            WE => \N__10985\
        );

    \mem_mem_5_2_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \mem_mem_5_2_physical_RDATA_wire\,
            RADDR => \mem_mem_5_2_physical_RADDR_wire\,
            WADDR => \mem_mem_5_2_physical_WADDR_wire\,
            MASK => \mem_mem_5_2_physical_MASK_wire\,
            WDATA => \mem_mem_5_2_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__4903\,
            RE => \N__10636\,
            WCLKE => \N__10317\,
            WCLK => \N__8742\,
            WE => \N__10632\
        );

    \mem_mem_2_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \mem_mem_2_0_physical_RDATA_wire\,
            RADDR => \mem_mem_2_0_physical_RADDR_wire\,
            WADDR => \mem_mem_2_0_physical_WADDR_wire\,
            MASK => \mem_mem_2_0_physical_MASK_wire\,
            WDATA => \mem_mem_2_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__4916\,
            RE => \N__10899\,
            WCLKE => \N__10196\,
            WCLK => \N__8757\,
            WE => \N__10924\
        );

    \mem_mem_1_3_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \mem_mem_1_3_physical_RDATA_wire\,
            RADDR => \mem_mem_1_3_physical_RADDR_wire\,
            WADDR => \mem_mem_1_3_physical_WADDR_wire\,
            MASK => \mem_mem_1_3_physical_MASK_wire\,
            WDATA => \mem_mem_1_3_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__4917\,
            RE => \N__10898\,
            WCLKE => \N__10136\,
            WCLK => \N__8756\,
            WE => \N__10878\
        );

    \mem_mem_4_2_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \mem_mem_4_2_physical_RDATA_wire\,
            RADDR => \mem_mem_4_2_physical_RADDR_wire\,
            WADDR => \mem_mem_4_2_physical_WADDR_wire\,
            MASK => \mem_mem_4_2_physical_MASK_wire\,
            WDATA => \mem_mem_4_2_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__4912\,
            RE => \N__10594\,
            WCLKE => \N__10281\,
            WCLK => \N__8751\,
            WE => \N__10703\
        );

    \mem_mem_7_2_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \mem_mem_7_2_physical_RDATA_wire\,
            RADDR => \mem_mem_7_2_physical_RADDR_wire\,
            WADDR => \mem_mem_7_2_physical_WADDR_wire\,
            MASK => \mem_mem_7_2_physical_MASK_wire\,
            WDATA => \mem_mem_7_2_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__4911\,
            RE => \N__10869\,
            WCLKE => \N__9565\,
            WCLK => \N__8752\,
            WE => \N__10921\
        );

    \mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \mem_mem_0_0_physical_WADDR_wire\,
            MASK => \mem_mem_0_0_physical_MASK_wire\,
            WDATA => \mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__4931\,
            RE => \N__10960\,
            WCLKE => \N__9938\,
            WCLK => \N__8770\,
            WE => \N__10931\
        );

    \mem_mem_3_3_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \mem_mem_3_3_physical_RDATA_wire\,
            RADDR => \mem_mem_3_3_physical_RADDR_wire\,
            WADDR => \mem_mem_3_3_physical_WADDR_wire\,
            MASK => \mem_mem_3_3_physical_MASK_wire\,
            WDATA => \mem_mem_3_3_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__4929\,
            RE => \N__10998\,
            WCLKE => \N__10247\,
            WCLK => \N__8771\,
            WE => \N__11000\
        );

    \mem_mem_6_2_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \mem_mem_6_2_physical_RDATA_wire\,
            RADDR => \mem_mem_6_2_physical_RADDR_wire\,
            WADDR => \mem_mem_6_2_physical_WADDR_wire\,
            MASK => \mem_mem_6_2_physical_MASK_wire\,
            WDATA => \mem_mem_6_2_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__4904\,
            RE => \N__10710\,
            WCLKE => \N__9598\,
            WCLK => \N__8745\,
            WE => \N__10787\
        );

    \mem_mem_5_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \mem_mem_5_1_physical_RDATA_wire\,
            RADDR => \mem_mem_5_1_physical_RADDR_wire\,
            WADDR => \mem_mem_5_1_physical_WADDR_wire\,
            MASK => \mem_mem_5_1_physical_MASK_wire\,
            WDATA => \mem_mem_5_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__4905\,
            RE => \N__10582\,
            WCLKE => \N__10324\,
            WCLK => \N__8744\,
            WE => \N__10589\
        );

    \mem_mem_2_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \mem_mem_2_1_physical_RDATA_wire\,
            RADDR => \mem_mem_2_1_physical_RADDR_wire\,
            WADDR => \mem_mem_2_1_physical_WADDR_wire\,
            MASK => \mem_mem_2_1_physical_MASK_wire\,
            WDATA => \mem_mem_2_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__4918\,
            RE => \N__10932\,
            WCLKE => \N__10197\,
            WCLK => \N__8759\,
            WE => \N__10925\
        );

    \mem_mem_1_2_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \mem_mem_1_2_physical_RDATA_wire\,
            RADDR => \mem_mem_1_2_physical_RADDR_wire\,
            WADDR => \mem_mem_1_2_physical_WADDR_wire\,
            MASK => \mem_mem_1_2_physical_MASK_wire\,
            WDATA => \mem_mem_1_2_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__4919\,
            RE => \N__10842\,
            WCLKE => \N__10137\,
            WCLK => \N__8758\,
            WE => \N__10877\
        );

    \mem_mem_4_3_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \mem_mem_4_3_physical_RDATA_wire\,
            RADDR => \mem_mem_4_3_physical_RADDR_wire\,
            WADDR => \mem_mem_4_3_physical_WADDR_wire\,
            MASK => \mem_mem_4_3_physical_MASK_wire\,
            WDATA => \mem_mem_4_3_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__4910\,
            RE => \N__10637\,
            WCLKE => \N__10272\,
            WCLK => \N__8749\,
            WE => \N__10590\
        );

    \mem_mem_0_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \mem_mem_0_1_physical_RDATA_wire\,
            RADDR => \mem_mem_0_1_physical_RADDR_wire\,
            WADDR => \mem_mem_0_1_physical_WADDR_wire\,
            MASK => \mem_mem_0_1_physical_MASK_wire\,
            WDATA => \mem_mem_0_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__4930\,
            RE => \N__10926\,
            WCLKE => \N__9937\,
            WCLK => \N__8769\,
            WE => \N__10927\
        );

    \mem_mem_3_2_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \mem_mem_3_2_physical_RDATA_wire\,
            RADDR => \mem_mem_3_2_physical_RADDR_wire\,
            WADDR => \mem_mem_3_2_physical_WADDR_wire\,
            MASK => \mem_mem_3_2_physical_MASK_wire\,
            WDATA => \mem_mem_3_2_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__4927\,
            RE => \N__10991\,
            WCLKE => \N__10246\,
            WCLK => \N__8768\,
            WE => \N__10999\
        );

    \mem_mem_6_3_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \mem_mem_6_3_physical_RDATA_wire\,
            RADDR => \mem_mem_6_3_physical_RADDR_wire\,
            WADDR => \mem_mem_6_3_physical_WADDR_wire\,
            MASK => \mem_mem_6_3_physical_MASK_wire\,
            WDATA => \mem_mem_6_3_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__4906\,
            RE => \N__10786\,
            WCLKE => \N__9602\,
            WCLK => \N__8747\,
            WE => \N__10788\
        );

    \mem_mem_5_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \mem_mem_5_0_physical_RDATA_wire\,
            RADDR => \mem_mem_5_0_physical_RADDR_wire\,
            WADDR => \mem_mem_5_0_physical_WADDR_wire\,
            MASK => \mem_mem_5_0_physical_MASK_wire\,
            WDATA => \mem_mem_5_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__4908\,
            RE => \N__10530\,
            WCLKE => \N__10325\,
            WCLK => \N__8746\,
            WE => \N__10631\
        );

    \mem_mem_2_2_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \mem_mem_2_2_physical_RDATA_wire\,
            RADDR => \mem_mem_2_2_physical_RADDR_wire\,
            WADDR => \mem_mem_2_2_physical_WADDR_wire\,
            MASK => \mem_mem_2_2_physical_MASK_wire\,
            WDATA => \mem_mem_2_2_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__4920\,
            RE => \N__10933\,
            WCLKE => \N__10198\,
            WCLK => \N__8761\,
            WE => \N__10961\
        );

    \mem_mem_7_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \mem_mem_7_1_physical_RDATA_wire\,
            RADDR => \mem_mem_7_1_physical_RADDR_wire\,
            WADDR => \mem_mem_7_1_physical_WADDR_wire\,
            MASK => \mem_mem_7_1_physical_MASK_wire\,
            WDATA => \mem_mem_7_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__4909\,
            RE => \N__10868\,
            WCLKE => \N__9558\,
            WCLK => \N__8750\,
            WE => \N__10864\
        );

    \mem_mem_1_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \mem_mem_1_1_physical_RDATA_wire\,
            RADDR => \mem_mem_1_1_physical_RADDR_wire\,
            WADDR => \mem_mem_1_1_physical_WADDR_wire\,
            MASK => \mem_mem_1_1_physical_MASK_wire\,
            WDATA => \mem_mem_1_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__4921\,
            RE => \N__10828\,
            WCLKE => \N__10144\,
            WCLK => \N__8760\,
            WE => \N__10816\
        );

    \mem_mem_4_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \mem_mem_4_0_physical_RDATA_wire\,
            RADDR => \mem_mem_4_0_physical_RADDR_wire\,
            WADDR => \mem_mem_4_0_physical_WADDR_wire\,
            MASK => \mem_mem_4_0_physical_MASK_wire\,
            WDATA => \mem_mem_4_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__4915\,
            RE => \N__10811\,
            WCLKE => \N__10289\,
            WCLK => \N__8754\,
            WE => \N__10740\
        );

    \mem_mem_2_3_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \mem_mem_2_3_physical_RDATA_wire\,
            RADDR => \mem_mem_2_3_physical_RADDR_wire\,
            WADDR => \mem_mem_2_3_physical_WADDR_wire\,
            MASK => \mem_mem_2_3_physical_MASK_wire\,
            WDATA => \mem_mem_2_3_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__4922\,
            RE => \N__10963\,
            WCLKE => \N__10202\,
            WCLK => \N__8763\,
            WE => \N__10962\
        );

    \mem_mem_7_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \mem_mem_7_0_physical_RDATA_wire\,
            RADDR => \mem_mem_7_0_physical_RADDR_wire\,
            WADDR => \mem_mem_7_0_physical_WADDR_wire\,
            MASK => \mem_mem_7_0_physical_MASK_wire\,
            WDATA => \mem_mem_7_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__4907\,
            RE => \N__10798\,
            WCLKE => \N__9541\,
            WCLK => \N__8748\,
            WE => \N__10863\
        );

    \mem_mem_1_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \mem_mem_1_0_physical_RDATA_wire\,
            RADDR => \mem_mem_1_0_physical_RADDR_wire\,
            WADDR => \mem_mem_1_0_physical_WADDR_wire\,
            MASK => \mem_mem_1_0_physical_MASK_wire\,
            WDATA => \mem_mem_1_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__4924\,
            RE => \N__10876\,
            WCLKE => \N__10145\,
            WCLK => \N__8762\,
            WE => \N__10812\
        );

    \mem_mem_4_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \mem_mem_4_1_physical_RDATA_wire\,
            RADDR => \mem_mem_4_1_physical_RADDR_wire\,
            WADDR => \mem_mem_4_1_physical_WADDR_wire\,
            MASK => \mem_mem_4_1_physical_MASK_wire\,
            WDATA => \mem_mem_4_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__4914\,
            RE => \N__10638\,
            WCLKE => \N__10288\,
            WCLK => \N__8753\,
            WE => \N__10736\
        );

    \mem_mem_0_2_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \mem_mem_0_2_physical_RDATA_wire\,
            RADDR => \mem_mem_0_2_physical_RADDR_wire\,
            WADDR => \mem_mem_0_2_physical_WADDR_wire\,
            MASK => \mem_mem_0_2_physical_MASK_wire\,
            WDATA => \mem_mem_0_2_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__4928\,
            RE => \N__10920\,
            WCLKE => \N__9936\,
            WCLK => \N__8767\,
            WE => \N__10862\
        );

    \mem_mem_3_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \mem_mem_3_1_physical_RDATA_wire\,
            RADDR => \mem_mem_3_1_physical_RADDR_wire\,
            WADDR => \mem_mem_3_1_physical_WADDR_wire\,
            MASK => \mem_mem_3_1_physical_MASK_wire\,
            WDATA => \mem_mem_3_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__4925\,
            RE => \N__10990\,
            WCLKE => \N__10239\,
            WCLK => \N__8766\,
            WE => \N__10986\
        );

    \mem_mem_6_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \mem_mem_6_0_physical_RDATA_wire\,
            RADDR => \mem_mem_6_0_physical_RADDR_wire\,
            WADDR => \mem_mem_6_0_physical_WADDR_wire\,
            MASK => \mem_mem_6_0_physical_MASK_wire\,
            WDATA => \mem_mem_6_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__4900\,
            RE => \N__10641\,
            WCLKE => \N__9587\,
            WCLK => \N__8741\,
            WE => \N__10704\
        );

    \mem_mem_5_3_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \mem_mem_5_3_physical_RDATA_wire\,
            RADDR => \mem_mem_5_3_physical_RADDR_wire\,
            WADDR => \mem_mem_5_3_physical_WADDR_wire\,
            MASK => \mem_mem_5_3_physical_MASK_wire\,
            WDATA => \mem_mem_5_3_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__4901\,
            RE => \N__10640\,
            WCLKE => \N__10300\,
            WCLK => \N__8740\,
            WE => \N__10639\
        );

    \mem_mem_7_3_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \mem_mem_7_3_physical_RDATA_wire\,
            RADDR => \mem_mem_7_3_physical_RADDR_wire\,
            WADDR => \mem_mem_7_3_physical_WADDR_wire\,
            MASK => \mem_mem_7_3_physical_MASK_wire\,
            WDATA => \mem_mem_7_3_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__4913\,
            RE => \N__10922\,
            WCLKE => \N__9566\,
            WCLK => \N__8755\,
            WE => \N__10923\
        );

    \mem_mem_0_3_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \mem_mem_0_3_physical_RDATA_wire\,
            RADDR => \mem_mem_0_3_physical_RADDR_wire\,
            WADDR => \mem_mem_0_3_physical_WADDR_wire\,
            MASK => \mem_mem_0_3_physical_MASK_wire\,
            WDATA => \mem_mem_0_3_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__4926\,
            RE => \N__10885\,
            WCLKE => \N__9935\,
            WCLK => \N__8765\,
            WE => \N__10858\
        );

    \mem_mem_6_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 3,
            READ_MODE => 3,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \mem_mem_6_1_physical_RDATA_wire\,
            RADDR => \mem_mem_6_1_physical_RADDR_wire\,
            WADDR => \mem_mem_6_1_physical_WADDR_wire\,
            MASK => \mem_mem_6_1_physical_MASK_wire\,
            WDATA => \mem_mem_6_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__4902\,
            RE => \N__10709\,
            WCLKE => \N__9597\,
            WCLK => \N__8743\,
            WE => \N__10705\
        );

    \wclk_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__13189\,
            GLOBALBUFFEROUTPUT => wclk_c_g
        );

    \wclk_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13191\,
            DIN => \N__13190\,
            DOUT => \N__13189\,
            PACKAGEPIN => wclk_wire
        );

    \wclk_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13191\,
            PADOUT => \N__13190\,
            PADIN => \N__13189\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \rclk_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__13179\,
            GLOBALBUFFEROUTPUT => rclk_c_g
        );

    \rclk_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13181\,
            DIN => \N__13180\,
            DOUT => \N__13179\,
            PACKAGEPIN => rclk_wire
        );

    \rclk_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13181\,
            PADOUT => \N__13180\,
            PADIN => \N__13179\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \waddr_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13170\,
            DIN => \N__13169\,
            DOUT => \N__13168\,
            PACKAGEPIN => waddr_wire(0)
        );

    \waddr_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13170\,
            PADOUT => \N__13169\,
            PADIN => \N__13168\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => waddr_c_0,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \dout_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13161\,
            DIN => \N__13160\,
            DOUT => \N__13159\,
            PACKAGEPIN => dout_wire(3)
        );

    \dout_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13161\,
            PADOUT => \N__13160\,
            PADIN => \N__13159\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11819\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \waddr_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13152\,
            DIN => \N__13151\,
            DOUT => \N__13150\,
            PACKAGEPIN => waddr_wire(12)
        );

    \waddr_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13152\,
            PADOUT => \N__13151\,
            PADIN => \N__13150\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => waddr_c_12,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \waddr_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13143\,
            DIN => \N__13142\,
            DOUT => \N__13141\,
            PACKAGEPIN => waddr_wire(4)
        );

    \waddr_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13143\,
            PADOUT => \N__13142\,
            PADIN => \N__13141\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => waddr_c_4,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \dout_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13134\,
            DIN => \N__13133\,
            DOUT => \N__13132\,
            PACKAGEPIN => dout_wire(6)
        );

    \dout_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13134\,
            PADOUT => \N__13133\,
            PADIN => \N__13132\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11522\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \raddr_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13125\,
            DIN => \N__13124\,
            DOUT => \N__13123\,
            PACKAGEPIN => raddr_wire(3)
        );

    \raddr_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13125\,
            PADOUT => \N__13124\,
            PADIN => \N__13123\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => raddr_c_3,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \din_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13116\,
            DIN => \N__13115\,
            DOUT => \N__13114\,
            PACKAGEPIN => din_wire(0)
        );

    \din_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13116\,
            PADOUT => \N__13115\,
            PADIN => \N__13114\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => din_c_0,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \waddr_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13107\,
            DIN => \N__13106\,
            DOUT => \N__13105\,
            PACKAGEPIN => waddr_wire(3)
        );

    \waddr_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13107\,
            PADOUT => \N__13106\,
            PADIN => \N__13105\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => waddr_c_3,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \raddr_ibuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13098\,
            DIN => \N__13097\,
            DOUT => \N__13096\,
            PACKAGEPIN => raddr_wire(11)
        );

    \raddr_ibuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000000"
        )
    port map (
            PADOEN => \N__13098\,
            PADOUT => \N__13097\,
            PADIN => \N__13096\,
            CLOCKENABLE => \VCCG0\,
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \mem_radregZ0Z_11\,
            DOUT0 => '0',
            INPUTCLK => \N__4932\,
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \raddr_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13089\,
            DIN => \N__13088\,
            DOUT => \N__13087\,
            PACKAGEPIN => raddr_wire(4)
        );

    \raddr_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13089\,
            PADOUT => \N__13088\,
            PADIN => \N__13087\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => raddr_c_4,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \waddr_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13080\,
            DIN => \N__13079\,
            DOUT => \N__13078\,
            PACKAGEPIN => waddr_wire(8)
        );

    \waddr_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13080\,
            PADOUT => \N__13079\,
            PADIN => \N__13078\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => waddr_c_8,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \dout_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13071\,
            DIN => \N__13070\,
            DOUT => \N__13069\,
            PACKAGEPIN => dout_wire(2)
        );

    \dout_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13071\,
            PADOUT => \N__13070\,
            PADIN => \N__13069\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11102\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \waddr_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13062\,
            DIN => \N__13061\,
            DOUT => \N__13060\,
            PACKAGEPIN => waddr_wire(13)
        );

    \waddr_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13062\,
            PADOUT => \N__13061\,
            PADIN => \N__13060\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => waddr_c_13,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \din_ibuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13053\,
            DIN => \N__13052\,
            DOUT => \N__13051\,
            PACKAGEPIN => din_wire(4)
        );

    \din_ibuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13053\,
            PADOUT => \N__13052\,
            PADIN => \N__13051\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => din_c_4,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \waddr_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13044\,
            DIN => \N__13043\,
            DOUT => \N__13042\,
            PACKAGEPIN => waddr_wire(7)
        );

    \waddr_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13044\,
            PADOUT => \N__13043\,
            PADIN => \N__13042\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => waddr_c_7,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \dout_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13035\,
            DIN => \N__13034\,
            DOUT => \N__13033\,
            PACKAGEPIN => dout_wire(5)
        );

    \dout_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__13035\,
            PADOUT => \N__13034\,
            PADIN => \N__13033\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__12482\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \raddr_ibuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13026\,
            DIN => \N__13025\,
            DOUT => \N__13024\,
            PACKAGEPIN => raddr_wire(0)
        );

    \raddr_ibuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13026\,
            PADOUT => \N__13025\,
            PADIN => \N__13024\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => raddr_c_0,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \din_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13017\,
            DIN => \N__13016\,
            DOUT => \N__13015\,
            PACKAGEPIN => din_wire(1)
        );

    \din_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13017\,
            PADOUT => \N__13016\,
            PADIN => \N__13015\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => din_c_1,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \waddr_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__13008\,
            DIN => \N__13007\,
            DOUT => \N__13006\,
            PACKAGEPIN => waddr_wire(2)
        );

    \waddr_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__13008\,
            PADOUT => \N__13007\,
            PADIN => \N__13006\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => waddr_c_2,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \raddr_ibuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12999\,
            DIN => \N__12998\,
            DOUT => \N__12997\,
            PACKAGEPIN => raddr_wire(10)
        );

    \raddr_ibuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12999\,
            PADOUT => \N__12998\,
            PADIN => \N__12997\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => raddr_c_10,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \raddr_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12990\,
            DIN => \N__12989\,
            DOUT => \N__12988\,
            PACKAGEPIN => raddr_wire(5)
        );

    \raddr_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12990\,
            PADOUT => \N__12989\,
            PADIN => \N__12988\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => raddr_c_5,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \dout_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12981\,
            DIN => \N__12980\,
            DOUT => \N__12979\,
            PACKAGEPIN => dout_wire(1)
        );

    \dout_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12981\,
            PADOUT => \N__12980\,
            PADIN => \N__12979\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10370\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \din_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12972\,
            DIN => \N__12971\,
            DOUT => \N__12970\,
            PACKAGEPIN => din_wire(5)
        );

    \din_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12972\,
            PADOUT => \N__12971\,
            PADIN => \N__12970\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => din_c_5,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \waddr_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12963\,
            DIN => \N__12962\,
            DOUT => \N__12961\,
            PACKAGEPIN => waddr_wire(6)
        );

    \waddr_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12963\,
            PADOUT => \N__12962\,
            PADIN => \N__12961\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => waddr_c_6,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \dout_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12954\,
            DIN => \N__12953\,
            DOUT => \N__12952\,
            PACKAGEPIN => dout_wire(4)
        );

    \dout_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12954\,
            PADOUT => \N__12953\,
            PADIN => \N__12952\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11552\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \raddr_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12945\,
            DIN => \N__12944\,
            DOUT => \N__12943\,
            PACKAGEPIN => raddr_wire(1)
        );

    \raddr_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12945\,
            PADOUT => \N__12944\,
            PADIN => \N__12943\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => raddr_c_1,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \raddr_ibuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12936\,
            DIN => \N__12935\,
            DOUT => \N__12934\,
            PACKAGEPIN => raddr_wire(8)
        );

    \raddr_ibuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12936\,
            PADOUT => \N__12935\,
            PADIN => \N__12934\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => raddr_c_8,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \waddr_ibuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12927\,
            DIN => \N__12926\,
            DOUT => \N__12925\,
            PACKAGEPIN => waddr_wire(10)
        );

    \waddr_ibuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12927\,
            PADOUT => \N__12926\,
            PADIN => \N__12925\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => waddr_c_10,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \din_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12918\,
            DIN => \N__12917\,
            DOUT => \N__12916\,
            PACKAGEPIN => din_wire(2)
        );

    \din_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12918\,
            PADOUT => \N__12917\,
            PADIN => \N__12916\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => din_c_2,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \raddr_ibuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12909\,
            DIN => \N__12908\,
            DOUT => \N__12907\,
            PACKAGEPIN => raddr_wire(13)
        );

    \raddr_ibuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000000"
        )
    port map (
            PADOEN => \N__12909\,
            PADOUT => \N__12908\,
            PADIN => \N__12907\,
            CLOCKENABLE => \VCCG0\,
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \mem_radregZ0Z_13\,
            DOUT0 => '0',
            INPUTCLK => \N__4934\,
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \dout_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12900\,
            DIN => \N__12899\,
            DOUT => \N__12898\,
            PACKAGEPIN => dout_wire(0)
        );

    \dout_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12900\,
            PADOUT => \N__12899\,
            PADIN => \N__12898\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__10343\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \din_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12891\,
            DIN => \N__12890\,
            DOUT => \N__12889\,
            PACKAGEPIN => din_wire(6)
        );

    \din_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12891\,
            PADOUT => \N__12890\,
            PADIN => \N__12889\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => din_c_6,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \waddr_ibuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12882\,
            DIN => \N__12881\,
            DOUT => \N__12880\,
            PACKAGEPIN => waddr_wire(1)
        );

    \waddr_ibuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12882\,
            PADOUT => \N__12881\,
            PADIN => \N__12880\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => waddr_c_1,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \raddr_ibuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12873\,
            DIN => \N__12872\,
            DOUT => \N__12871\,
            PACKAGEPIN => raddr_wire(6)
        );

    \raddr_ibuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12873\,
            PADOUT => \N__12872\,
            PADIN => \N__12871\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => raddr_c_6,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \raddr_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12864\,
            DIN => \N__12863\,
            DOUT => \N__12862\,
            PACKAGEPIN => raddr_wire(9)
        );

    \raddr_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12864\,
            PADOUT => \N__12863\,
            PADIN => \N__12862\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => raddr_c_9,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \waddr_ibuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12855\,
            DIN => \N__12854\,
            DOUT => \N__12853\,
            PACKAGEPIN => waddr_wire(11)
        );

    \waddr_ibuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12855\,
            PADOUT => \N__12854\,
            PADIN => \N__12853\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => waddr_c_11,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \din_ibuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12846\,
            DIN => \N__12845\,
            DOUT => \N__12844\,
            PACKAGEPIN => din_wire(3)
        );

    \din_ibuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12846\,
            PADOUT => \N__12845\,
            PADIN => \N__12844\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => din_c_3,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \raddr_ibuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12837\,
            DIN => \N__12836\,
            DOUT => \N__12835\,
            PACKAGEPIN => raddr_wire(12)
        );

    \raddr_ibuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000000"
        )
    port map (
            PADOEN => \N__12837\,
            PADOUT => \N__12836\,
            PADIN => \N__12835\,
            CLOCKENABLE => \VCCG0\,
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => \mem_radregZ0Z_12\,
            DOUT0 => '0',
            INPUTCLK => \N__4933\,
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \waddr_ibuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12828\,
            DIN => \N__12827\,
            DOUT => \N__12826\,
            PACKAGEPIN => waddr_wire(5)
        );

    \waddr_ibuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12828\,
            PADOUT => \N__12827\,
            PADIN => \N__12826\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => waddr_c_5,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \write_en_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12819\,
            DIN => \N__12818\,
            DOUT => \N__12817\,
            PACKAGEPIN => write_en_wire
        );

    \write_en_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12819\,
            PADOUT => \N__12818\,
            PADIN => \N__12817\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => write_en_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \dout_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12810\,
            DIN => \N__12809\,
            DOUT => \N__12808\,
            PACKAGEPIN => dout_wire(7)
        );

    \dout_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__12810\,
            PADOUT => \N__12809\,
            PADIN => \N__12808\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__11048\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \raddr_ibuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12801\,
            DIN => \N__12800\,
            DOUT => \N__12799\,
            PACKAGEPIN => raddr_wire(2)
        );

    \raddr_ibuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12801\,
            PADOUT => \N__12800\,
            PADIN => \N__12799\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => raddr_c_2,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \din_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12792\,
            DIN => \N__12791\,
            DOUT => \N__12790\,
            PACKAGEPIN => din_wire(7)
        );

    \din_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12792\,
            PADOUT => \N__12791\,
            PADIN => \N__12790\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => din_c_7,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \raddr_ibuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12783\,
            DIN => \N__12782\,
            DOUT => \N__12781\,
            PACKAGEPIN => raddr_wire(7)
        );

    \raddr_ibuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12783\,
            PADOUT => \N__12782\,
            PADIN => \N__12781\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => raddr_c_7,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \waddr_ibuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__12774\,
            DIN => \N__12773\,
            DOUT => \N__12772\,
            PACKAGEPIN => waddr_wire(9)
        );

    \waddr_ibuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__12774\,
            PADOUT => \N__12773\,
            PADIN => \N__12772\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => waddr_c_9,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__3118\ : InMux
    port map (
            O => \N__12755\,
            I => \N__12752\
        );

    \I__3117\ : LocalMux
    port map (
            O => \N__12752\,
            I => \N__12744\
        );

    \I__3116\ : InMux
    port map (
            O => \N__12751\,
            I => \N__12739\
        );

    \I__3115\ : InMux
    port map (
            O => \N__12750\,
            I => \N__12739\
        );

    \I__3114\ : InMux
    port map (
            O => \N__12749\,
            I => \N__12736\
        );

    \I__3113\ : InMux
    port map (
            O => \N__12748\,
            I => \N__12731\
        );

    \I__3112\ : InMux
    port map (
            O => \N__12747\,
            I => \N__12731\
        );

    \I__3111\ : Span4Mux_v
    port map (
            O => \N__12744\,
            I => \N__12719\
        );

    \I__3110\ : LocalMux
    port map (
            O => \N__12739\,
            I => \N__12719\
        );

    \I__3109\ : LocalMux
    port map (
            O => \N__12736\,
            I => \N__12719\
        );

    \I__3108\ : LocalMux
    port map (
            O => \N__12731\,
            I => \N__12719\
        );

    \I__3107\ : InMux
    port map (
            O => \N__12730\,
            I => \N__12716\
        );

    \I__3106\ : InMux
    port map (
            O => \N__12729\,
            I => \N__12708\
        );

    \I__3105\ : InMux
    port map (
            O => \N__12728\,
            I => \N__12705\
        );

    \I__3104\ : Span4Mux_h
    port map (
            O => \N__12719\,
            I => \N__12700\
        );

    \I__3103\ : LocalMux
    port map (
            O => \N__12716\,
            I => \N__12700\
        );

    \I__3102\ : InMux
    port map (
            O => \N__12715\,
            I => \N__12697\
        );

    \I__3101\ : InMux
    port map (
            O => \N__12714\,
            I => \N__12694\
        );

    \I__3100\ : InMux
    port map (
            O => \N__12713\,
            I => \N__12691\
        );

    \I__3099\ : InMux
    port map (
            O => \N__12712\,
            I => \N__12688\
        );

    \I__3098\ : InMux
    port map (
            O => \N__12711\,
            I => \N__12685\
        );

    \I__3097\ : LocalMux
    port map (
            O => \N__12708\,
            I => \N__12680\
        );

    \I__3096\ : LocalMux
    port map (
            O => \N__12705\,
            I => \N__12677\
        );

    \I__3095\ : Span4Mux_v
    port map (
            O => \N__12700\,
            I => \N__12674\
        );

    \I__3094\ : LocalMux
    port map (
            O => \N__12697\,
            I => \N__12667\
        );

    \I__3093\ : LocalMux
    port map (
            O => \N__12694\,
            I => \N__12667\
        );

    \I__3092\ : LocalMux
    port map (
            O => \N__12691\,
            I => \N__12667\
        );

    \I__3091\ : LocalMux
    port map (
            O => \N__12688\,
            I => \N__12662\
        );

    \I__3090\ : LocalMux
    port map (
            O => \N__12685\,
            I => \N__12662\
        );

    \I__3089\ : InMux
    port map (
            O => \N__12684\,
            I => \N__12659\
        );

    \I__3088\ : InMux
    port map (
            O => \N__12683\,
            I => \N__12656\
        );

    \I__3087\ : Span4Mux_v
    port map (
            O => \N__12680\,
            I => \N__12651\
        );

    \I__3086\ : Span4Mux_v
    port map (
            O => \N__12677\,
            I => \N__12651\
        );

    \I__3085\ : Span4Mux_h
    port map (
            O => \N__12674\,
            I => \N__12648\
        );

    \I__3084\ : Span4Mux_h
    port map (
            O => \N__12667\,
            I => \N__12645\
        );

    \I__3083\ : Span4Mux_h
    port map (
            O => \N__12662\,
            I => \N__12638\
        );

    \I__3082\ : LocalMux
    port map (
            O => \N__12659\,
            I => \N__12638\
        );

    \I__3081\ : LocalMux
    port map (
            O => \N__12656\,
            I => \N__12638\
        );

    \I__3080\ : Span4Mux_h
    port map (
            O => \N__12651\,
            I => \N__12635\
        );

    \I__3079\ : Span4Mux_h
    port map (
            O => \N__12648\,
            I => \N__12632\
        );

    \I__3078\ : Span4Mux_h
    port map (
            O => \N__12645\,
            I => \N__12629\
        );

    \I__3077\ : Span4Mux_h
    port map (
            O => \N__12638\,
            I => \N__12626\
        );

    \I__3076\ : Sp12to4
    port map (
            O => \N__12635\,
            I => \N__12623\
        );

    \I__3075\ : Sp12to4
    port map (
            O => \N__12632\,
            I => \N__12620\
        );

    \I__3074\ : Sp12to4
    port map (
            O => \N__12629\,
            I => \N__12615\
        );

    \I__3073\ : Sp12to4
    port map (
            O => \N__12626\,
            I => \N__12615\
        );

    \I__3072\ : Span12Mux_h
    port map (
            O => \N__12623\,
            I => \N__12612\
        );

    \I__3071\ : Span12Mux_h
    port map (
            O => \N__12620\,
            I => \N__12609\
        );

    \I__3070\ : Span12Mux_v
    port map (
            O => \N__12615\,
            I => \N__12606\
        );

    \I__3069\ : Span12Mux_v
    port map (
            O => \N__12612\,
            I => \N__12603\
        );

    \I__3068\ : Span12Mux_v
    port map (
            O => \N__12609\,
            I => \N__12598\
        );

    \I__3067\ : Span12Mux_h
    port map (
            O => \N__12606\,
            I => \N__12598\
        );

    \I__3066\ : Odrv12
    port map (
            O => \N__12603\,
            I => \mem_radregZ0Z_12\
        );

    \I__3065\ : Odrv12
    port map (
            O => \N__12598\,
            I => \mem_radregZ0Z_12\
        );

    \I__3064\ : CascadeMux
    port map (
            O => \N__12593\,
            I => \dout_obuf_RNO_2Z0Z_5_cascade_\
        );

    \I__3063\ : InMux
    port map (
            O => \N__12590\,
            I => \N__12587\
        );

    \I__3062\ : LocalMux
    port map (
            O => \N__12587\,
            I => \mem_N_140\
        );

    \I__3061\ : InMux
    port map (
            O => \N__12584\,
            I => \N__12581\
        );

    \I__3060\ : LocalMux
    port map (
            O => \N__12581\,
            I => \N__12575\
        );

    \I__3059\ : InMux
    port map (
            O => \N__12580\,
            I => \N__12572\
        );

    \I__3058\ : InMux
    port map (
            O => \N__12579\,
            I => \N__12567\
        );

    \I__3057\ : InMux
    port map (
            O => \N__12578\,
            I => \N__12567\
        );

    \I__3056\ : Span4Mux_v
    port map (
            O => \N__12575\,
            I => \N__12561\
        );

    \I__3055\ : LocalMux
    port map (
            O => \N__12572\,
            I => \N__12561\
        );

    \I__3054\ : LocalMux
    port map (
            O => \N__12567\,
            I => \N__12555\
        );

    \I__3053\ : InMux
    port map (
            O => \N__12566\,
            I => \N__12552\
        );

    \I__3052\ : Span4Mux_v
    port map (
            O => \N__12561\,
            I => \N__12549\
        );

    \I__3051\ : InMux
    port map (
            O => \N__12560\,
            I => \N__12546\
        );

    \I__3050\ : InMux
    port map (
            O => \N__12559\,
            I => \N__12543\
        );

    \I__3049\ : InMux
    port map (
            O => \N__12558\,
            I => \N__12540\
        );

    \I__3048\ : Span4Mux_v
    port map (
            O => \N__12555\,
            I => \N__12535\
        );

    \I__3047\ : LocalMux
    port map (
            O => \N__12552\,
            I => \N__12535\
        );

    \I__3046\ : Span4Mux_h
    port map (
            O => \N__12549\,
            I => \N__12532\
        );

    \I__3045\ : LocalMux
    port map (
            O => \N__12546\,
            I => \N__12529\
        );

    \I__3044\ : LocalMux
    port map (
            O => \N__12543\,
            I => \N__12524\
        );

    \I__3043\ : LocalMux
    port map (
            O => \N__12540\,
            I => \N__12524\
        );

    \I__3042\ : Span4Mux_h
    port map (
            O => \N__12535\,
            I => \N__12521\
        );

    \I__3041\ : Sp12to4
    port map (
            O => \N__12532\,
            I => \N__12516\
        );

    \I__3040\ : Span12Mux_h
    port map (
            O => \N__12529\,
            I => \N__12516\
        );

    \I__3039\ : Span12Mux_h
    port map (
            O => \N__12524\,
            I => \N__12513\
        );

    \I__3038\ : Sp12to4
    port map (
            O => \N__12521\,
            I => \N__12510\
        );

    \I__3037\ : Span12Mux_h
    port map (
            O => \N__12516\,
            I => \N__12507\
        );

    \I__3036\ : Span12Mux_h
    port map (
            O => \N__12513\,
            I => \N__12504\
        );

    \I__3035\ : Span12Mux_v
    port map (
            O => \N__12510\,
            I => \N__12501\
        );

    \I__3034\ : Span12Mux_v
    port map (
            O => \N__12507\,
            I => \N__12498\
        );

    \I__3033\ : Span12Mux_v
    port map (
            O => \N__12504\,
            I => \N__12493\
        );

    \I__3032\ : Span12Mux_h
    port map (
            O => \N__12501\,
            I => \N__12493\
        );

    \I__3031\ : Odrv12
    port map (
            O => \N__12498\,
            I => \mem_radregZ0Z_11\
        );

    \I__3030\ : Odrv12
    port map (
            O => \N__12493\,
            I => \mem_radregZ0Z_11\
        );

    \I__3029\ : InMux
    port map (
            O => \N__12488\,
            I => \N__12485\
        );

    \I__3028\ : LocalMux
    port map (
            O => \N__12485\,
            I => \mem_N_139\
        );

    \I__3027\ : IoInMux
    port map (
            O => \N__12482\,
            I => \N__12479\
        );

    \I__3026\ : LocalMux
    port map (
            O => \N__12479\,
            I => \N__12476\
        );

    \I__3025\ : IoSpan4Mux
    port map (
            O => \N__12476\,
            I => \N__12473\
        );

    \I__3024\ : Span4Mux_s2_h
    port map (
            O => \N__12473\,
            I => \N__12470\
        );

    \I__3023\ : Span4Mux_h
    port map (
            O => \N__12470\,
            I => \N__12467\
        );

    \I__3022\ : Span4Mux_h
    port map (
            O => \N__12467\,
            I => \N__12464\
        );

    \I__3021\ : Odrv4
    port map (
            O => \N__12464\,
            I => dout_c_5
        );

    \I__3020\ : InMux
    port map (
            O => \N__12461\,
            I => \N__12458\
        );

    \I__3019\ : LocalMux
    port map (
            O => \N__12458\,
            I => \N__12455\
        );

    \I__3018\ : Odrv12
    port map (
            O => \N__12455\,
            I => mem_out_bus6_5
        );

    \I__3017\ : InMux
    port map (
            O => \N__12452\,
            I => \N__12449\
        );

    \I__3016\ : LocalMux
    port map (
            O => \N__12449\,
            I => \N__12446\
        );

    \I__3015\ : Span12Mux_h
    port map (
            O => \N__12446\,
            I => \N__12443\
        );

    \I__3014\ : Odrv12
    port map (
            O => \N__12443\,
            I => mem_out_bus2_5
        );

    \I__3013\ : InMux
    port map (
            O => \N__12440\,
            I => \N__12437\
        );

    \I__3012\ : LocalMux
    port map (
            O => \N__12437\,
            I => \N__12434\
        );

    \I__3011\ : Odrv12
    port map (
            O => \N__12434\,
            I => \dout_obuf_RNO_5Z0Z_5\
        );

    \I__3010\ : InMux
    port map (
            O => \N__12431\,
            I => \N__12425\
        );

    \I__3009\ : InMux
    port map (
            O => \N__12430\,
            I => \N__12425\
        );

    \I__3008\ : LocalMux
    port map (
            O => \N__12425\,
            I => \N__12420\
        );

    \I__3007\ : InMux
    port map (
            O => \N__12424\,
            I => \N__12415\
        );

    \I__3006\ : InMux
    port map (
            O => \N__12423\,
            I => \N__12415\
        );

    \I__3005\ : Span4Mux_s2_v
    port map (
            O => \N__12420\,
            I => \N__12408\
        );

    \I__3004\ : LocalMux
    port map (
            O => \N__12415\,
            I => \N__12408\
        );

    \I__3003\ : InMux
    port map (
            O => \N__12414\,
            I => \N__12403\
        );

    \I__3002\ : InMux
    port map (
            O => \N__12413\,
            I => \N__12403\
        );

    \I__3001\ : Span4Mux_v
    port map (
            O => \N__12408\,
            I => \N__12394\
        );

    \I__3000\ : LocalMux
    port map (
            O => \N__12403\,
            I => \N__12394\
        );

    \I__2999\ : InMux
    port map (
            O => \N__12402\,
            I => \N__12391\
        );

    \I__2998\ : CascadeMux
    port map (
            O => \N__12401\,
            I => \N__12388\
        );

    \I__2997\ : CascadeMux
    port map (
            O => \N__12400\,
            I => \N__12385\
        );

    \I__2996\ : InMux
    port map (
            O => \N__12399\,
            I => \N__12381\
        );

    \I__2995\ : Span4Mux_v
    port map (
            O => \N__12394\,
            I => \N__12376\
        );

    \I__2994\ : LocalMux
    port map (
            O => \N__12391\,
            I => \N__12376\
        );

    \I__2993\ : InMux
    port map (
            O => \N__12388\,
            I => \N__12369\
        );

    \I__2992\ : InMux
    port map (
            O => \N__12385\,
            I => \N__12369\
        );

    \I__2991\ : InMux
    port map (
            O => \N__12384\,
            I => \N__12369\
        );

    \I__2990\ : LocalMux
    port map (
            O => \N__12381\,
            I => \N__12366\
        );

    \I__2989\ : Span4Mux_v
    port map (
            O => \N__12376\,
            I => \N__12359\
        );

    \I__2988\ : LocalMux
    port map (
            O => \N__12369\,
            I => \N__12359\
        );

    \I__2987\ : Span4Mux_v
    port map (
            O => \N__12366\,
            I => \N__12354\
        );

    \I__2986\ : InMux
    port map (
            O => \N__12365\,
            I => \N__12351\
        );

    \I__2985\ : CascadeMux
    port map (
            O => \N__12364\,
            I => \N__12346\
        );

    \I__2984\ : Span4Mux_v
    port map (
            O => \N__12359\,
            I => \N__12342\
        );

    \I__2983\ : InMux
    port map (
            O => \N__12358\,
            I => \N__12339\
        );

    \I__2982\ : InMux
    port map (
            O => \N__12357\,
            I => \N__12336\
        );

    \I__2981\ : Span4Mux_v
    port map (
            O => \N__12354\,
            I => \N__12330\
        );

    \I__2980\ : LocalMux
    port map (
            O => \N__12351\,
            I => \N__12330\
        );

    \I__2979\ : InMux
    port map (
            O => \N__12350\,
            I => \N__12322\
        );

    \I__2978\ : InMux
    port map (
            O => \N__12349\,
            I => \N__12322\
        );

    \I__2977\ : InMux
    port map (
            O => \N__12346\,
            I => \N__12315\
        );

    \I__2976\ : InMux
    port map (
            O => \N__12345\,
            I => \N__12315\
        );

    \I__2975\ : Span4Mux_v
    port map (
            O => \N__12342\,
            I => \N__12306\
        );

    \I__2974\ : LocalMux
    port map (
            O => \N__12339\,
            I => \N__12306\
        );

    \I__2973\ : LocalMux
    port map (
            O => \N__12336\,
            I => \N__12306\
        );

    \I__2972\ : InMux
    port map (
            O => \N__12335\,
            I => \N__12303\
        );

    \I__2971\ : Span4Mux_v
    port map (
            O => \N__12330\,
            I => \N__12300\
        );

    \I__2970\ : InMux
    port map (
            O => \N__12329\,
            I => \N__12297\
        );

    \I__2969\ : InMux
    port map (
            O => \N__12328\,
            I => \N__12294\
        );

    \I__2968\ : InMux
    port map (
            O => \N__12327\,
            I => \N__12291\
        );

    \I__2967\ : LocalMux
    port map (
            O => \N__12322\,
            I => \N__12286\
        );

    \I__2966\ : InMux
    port map (
            O => \N__12321\,
            I => \N__12283\
        );

    \I__2965\ : InMux
    port map (
            O => \N__12320\,
            I => \N__12280\
        );

    \I__2964\ : LocalMux
    port map (
            O => \N__12315\,
            I => \N__12275\
        );

    \I__2963\ : InMux
    port map (
            O => \N__12314\,
            I => \N__12270\
        );

    \I__2962\ : InMux
    port map (
            O => \N__12313\,
            I => \N__12270\
        );

    \I__2961\ : Span4Mux_v
    port map (
            O => \N__12306\,
            I => \N__12265\
        );

    \I__2960\ : LocalMux
    port map (
            O => \N__12303\,
            I => \N__12265\
        );

    \I__2959\ : Span4Mux_v
    port map (
            O => \N__12300\,
            I => \N__12258\
        );

    \I__2958\ : LocalMux
    port map (
            O => \N__12297\,
            I => \N__12258\
        );

    \I__2957\ : LocalMux
    port map (
            O => \N__12294\,
            I => \N__12253\
        );

    \I__2956\ : LocalMux
    port map (
            O => \N__12291\,
            I => \N__12253\
        );

    \I__2955\ : InMux
    port map (
            O => \N__12290\,
            I => \N__12248\
        );

    \I__2954\ : InMux
    port map (
            O => \N__12289\,
            I => \N__12248\
        );

    \I__2953\ : Span12Mux_h
    port map (
            O => \N__12286\,
            I => \N__12245\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__12283\,
            I => \N__12240\
        );

    \I__2951\ : LocalMux
    port map (
            O => \N__12280\,
            I => \N__12240\
        );

    \I__2950\ : InMux
    port map (
            O => \N__12279\,
            I => \N__12235\
        );

    \I__2949\ : InMux
    port map (
            O => \N__12278\,
            I => \N__12235\
        );

    \I__2948\ : Span12Mux_h
    port map (
            O => \N__12275\,
            I => \N__12232\
        );

    \I__2947\ : LocalMux
    port map (
            O => \N__12270\,
            I => \N__12229\
        );

    \I__2946\ : Span4Mux_v
    port map (
            O => \N__12265\,
            I => \N__12226\
        );

    \I__2945\ : InMux
    port map (
            O => \N__12264\,
            I => \N__12221\
        );

    \I__2944\ : InMux
    port map (
            O => \N__12263\,
            I => \N__12221\
        );

    \I__2943\ : Span4Mux_v
    port map (
            O => \N__12258\,
            I => \N__12218\
        );

    \I__2942\ : Span12Mux_h
    port map (
            O => \N__12253\,
            I => \N__12215\
        );

    \I__2941\ : LocalMux
    port map (
            O => \N__12248\,
            I => \N__12212\
        );

    \I__2940\ : Span12Mux_h
    port map (
            O => \N__12245\,
            I => \N__12209\
        );

    \I__2939\ : Span12Mux_h
    port map (
            O => \N__12240\,
            I => \N__12206\
        );

    \I__2938\ : LocalMux
    port map (
            O => \N__12235\,
            I => \N__12203\
        );

    \I__2937\ : Span12Mux_h
    port map (
            O => \N__12232\,
            I => \N__12200\
        );

    \I__2936\ : Span12Mux_h
    port map (
            O => \N__12229\,
            I => \N__12197\
        );

    \I__2935\ : Sp12to4
    port map (
            O => \N__12226\,
            I => \N__12192\
        );

    \I__2934\ : LocalMux
    port map (
            O => \N__12221\,
            I => \N__12192\
        );

    \I__2933\ : Span4Mux_h
    port map (
            O => \N__12218\,
            I => \N__12189\
        );

    \I__2932\ : Span12Mux_h
    port map (
            O => \N__12215\,
            I => \N__12186\
        );

    \I__2931\ : Span12Mux_h
    port map (
            O => \N__12212\,
            I => \N__12183\
        );

    \I__2930\ : Span12Mux_v
    port map (
            O => \N__12209\,
            I => \N__12178\
        );

    \I__2929\ : Span12Mux_h
    port map (
            O => \N__12206\,
            I => \N__12178\
        );

    \I__2928\ : Span12Mux_h
    port map (
            O => \N__12203\,
            I => \N__12175\
        );

    \I__2927\ : Span12Mux_v
    port map (
            O => \N__12200\,
            I => \N__12170\
        );

    \I__2926\ : Span12Mux_h
    port map (
            O => \N__12197\,
            I => \N__12170\
        );

    \I__2925\ : Span12Mux_h
    port map (
            O => \N__12192\,
            I => \N__12165\
        );

    \I__2924\ : Sp12to4
    port map (
            O => \N__12189\,
            I => \N__12165\
        );

    \I__2923\ : Span12Mux_v
    port map (
            O => \N__12186\,
            I => \N__12160\
        );

    \I__2922\ : Span12Mux_h
    port map (
            O => \N__12183\,
            I => \N__12160\
        );

    \I__2921\ : Span12Mux_v
    port map (
            O => \N__12178\,
            I => \N__12155\
        );

    \I__2920\ : Span12Mux_h
    port map (
            O => \N__12175\,
            I => \N__12155\
        );

    \I__2919\ : Span12Mux_v
    port map (
            O => \N__12170\,
            I => \N__12150\
        );

    \I__2918\ : Span12Mux_h
    port map (
            O => \N__12165\,
            I => \N__12150\
        );

    \I__2917\ : Odrv12
    port map (
            O => \N__12160\,
            I => \mem_radregZ0Z_13\
        );

    \I__2916\ : Odrv12
    port map (
            O => \N__12155\,
            I => \mem_radregZ0Z_13\
        );

    \I__2915\ : Odrv12
    port map (
            O => \N__12150\,
            I => \mem_radregZ0Z_13\
        );

    \I__2914\ : InMux
    port map (
            O => \N__12143\,
            I => \N__12140\
        );

    \I__2913\ : LocalMux
    port map (
            O => \N__12140\,
            I => \N__12137\
        );

    \I__2912\ : Odrv12
    port map (
            O => \N__12137\,
            I => mem_out_bus7_5
        );

    \I__2911\ : InMux
    port map (
            O => \N__12134\,
            I => \N__12131\
        );

    \I__2910\ : LocalMux
    port map (
            O => \N__12131\,
            I => \N__12128\
        );

    \I__2909\ : Span12Mux_h
    port map (
            O => \N__12128\,
            I => \N__12125\
        );

    \I__2908\ : Odrv12
    port map (
            O => \N__12125\,
            I => mem_out_bus3_5
        );

    \I__2907\ : InMux
    port map (
            O => \N__12122\,
            I => \N__12119\
        );

    \I__2906\ : LocalMux
    port map (
            O => \N__12119\,
            I => \N__12116\
        );

    \I__2905\ : Span12Mux_v
    port map (
            O => \N__12116\,
            I => \N__12113\
        );

    \I__2904\ : Odrv12
    port map (
            O => \N__12113\,
            I => \dout_obuf_RNO_3Z0Z_5\
        );

    \I__2903\ : InMux
    port map (
            O => \N__12110\,
            I => \N__12107\
        );

    \I__2902\ : LocalMux
    port map (
            O => \N__12107\,
            I => \N__12104\
        );

    \I__2901\ : Span4Mux_v
    port map (
            O => \N__12104\,
            I => \N__12101\
        );

    \I__2900\ : Odrv4
    port map (
            O => \N__12101\,
            I => mem_out_bus6_6
        );

    \I__2899\ : InMux
    port map (
            O => \N__12098\,
            I => \N__12095\
        );

    \I__2898\ : LocalMux
    port map (
            O => \N__12095\,
            I => \N__12092\
        );

    \I__2897\ : Span4Mux_v
    port map (
            O => \N__12092\,
            I => \N__12089\
        );

    \I__2896\ : Sp12to4
    port map (
            O => \N__12089\,
            I => \N__12086\
        );

    \I__2895\ : Span12Mux_h
    port map (
            O => \N__12086\,
            I => \N__12083\
        );

    \I__2894\ : Odrv12
    port map (
            O => \N__12083\,
            I => mem_out_bus2_6
        );

    \I__2893\ : InMux
    port map (
            O => \N__12080\,
            I => \N__12077\
        );

    \I__2892\ : LocalMux
    port map (
            O => \N__12077\,
            I => \N__12074\
        );

    \I__2891\ : Span12Mux_v
    port map (
            O => \N__12074\,
            I => \N__12071\
        );

    \I__2890\ : Odrv12
    port map (
            O => \N__12071\,
            I => \dout_obuf_RNO_5Z0Z_6\
        );

    \I__2889\ : InMux
    port map (
            O => \N__12068\,
            I => \N__12065\
        );

    \I__2888\ : LocalMux
    port map (
            O => \N__12065\,
            I => \N__12062\
        );

    \I__2887\ : Odrv12
    port map (
            O => \N__12062\,
            I => mem_out_bus6_7
        );

    \I__2886\ : InMux
    port map (
            O => \N__12059\,
            I => \N__12056\
        );

    \I__2885\ : LocalMux
    port map (
            O => \N__12056\,
            I => \N__12053\
        );

    \I__2884\ : Span12Mux_h
    port map (
            O => \N__12053\,
            I => \N__12050\
        );

    \I__2883\ : Odrv12
    port map (
            O => \N__12050\,
            I => mem_out_bus2_7
        );

    \I__2882\ : InMux
    port map (
            O => \N__12047\,
            I => \N__12044\
        );

    \I__2881\ : LocalMux
    port map (
            O => \N__12044\,
            I => \N__12041\
        );

    \I__2880\ : Span4Mux_v
    port map (
            O => \N__12041\,
            I => \N__12038\
        );

    \I__2879\ : Span4Mux_v
    port map (
            O => \N__12038\,
            I => \N__12035\
        );

    \I__2878\ : Odrv4
    port map (
            O => \N__12035\,
            I => \dout_obuf_RNO_5Z0Z_7\
        );

    \I__2877\ : InMux
    port map (
            O => \N__12032\,
            I => \N__12029\
        );

    \I__2876\ : LocalMux
    port map (
            O => \N__12029\,
            I => \N__12026\
        );

    \I__2875\ : Odrv4
    port map (
            O => \N__12026\,
            I => mem_out_bus7_1
        );

    \I__2874\ : InMux
    port map (
            O => \N__12023\,
            I => \N__12020\
        );

    \I__2873\ : LocalMux
    port map (
            O => \N__12020\,
            I => \N__12017\
        );

    \I__2872\ : Span12Mux_h
    port map (
            O => \N__12017\,
            I => \N__12014\
        );

    \I__2871\ : Odrv12
    port map (
            O => \N__12014\,
            I => mem_out_bus3_1
        );

    \I__2870\ : InMux
    port map (
            O => \N__12011\,
            I => \N__12008\
        );

    \I__2869\ : LocalMux
    port map (
            O => \N__12008\,
            I => \N__12005\
        );

    \I__2868\ : Sp12to4
    port map (
            O => \N__12005\,
            I => \N__12002\
        );

    \I__2867\ : Span12Mux_v
    port map (
            O => \N__12002\,
            I => \N__11999\
        );

    \I__2866\ : Odrv12
    port map (
            O => \N__11999\,
            I => \dout_obuf_RNO_3Z0Z_1\
        );

    \I__2865\ : InMux
    port map (
            O => \N__11996\,
            I => \N__11993\
        );

    \I__2864\ : LocalMux
    port map (
            O => \N__11993\,
            I => \N__11990\
        );

    \I__2863\ : Span4Mux_v
    port map (
            O => \N__11990\,
            I => \N__11987\
        );

    \I__2862\ : Odrv4
    port map (
            O => \N__11987\,
            I => mem_out_bus7_4
        );

    \I__2861\ : InMux
    port map (
            O => \N__11984\,
            I => \N__11981\
        );

    \I__2860\ : LocalMux
    port map (
            O => \N__11981\,
            I => \N__11978\
        );

    \I__2859\ : Span4Mux_v
    port map (
            O => \N__11978\,
            I => \N__11975\
        );

    \I__2858\ : Sp12to4
    port map (
            O => \N__11975\,
            I => \N__11972\
        );

    \I__2857\ : Span12Mux_h
    port map (
            O => \N__11972\,
            I => \N__11969\
        );

    \I__2856\ : Odrv12
    port map (
            O => \N__11969\,
            I => mem_out_bus3_4
        );

    \I__2855\ : InMux
    port map (
            O => \N__11966\,
            I => \N__11963\
        );

    \I__2854\ : LocalMux
    port map (
            O => \N__11963\,
            I => \N__11960\
        );

    \I__2853\ : Span4Mux_v
    port map (
            O => \N__11960\,
            I => \N__11957\
        );

    \I__2852\ : Span4Mux_v
    port map (
            O => \N__11957\,
            I => \N__11954\
        );

    \I__2851\ : Span4Mux_v
    port map (
            O => \N__11954\,
            I => \N__11951\
        );

    \I__2850\ : Span4Mux_v
    port map (
            O => \N__11951\,
            I => \N__11948\
        );

    \I__2849\ : Odrv4
    port map (
            O => \N__11948\,
            I => \dout_obuf_RNO_3Z0Z_4\
        );

    \I__2848\ : InMux
    port map (
            O => \N__11945\,
            I => \N__11942\
        );

    \I__2847\ : LocalMux
    port map (
            O => \N__11942\,
            I => \N__11939\
        );

    \I__2846\ : Odrv4
    port map (
            O => \N__11939\,
            I => mem_out_bus7_7
        );

    \I__2845\ : InMux
    port map (
            O => \N__11936\,
            I => \N__11933\
        );

    \I__2844\ : LocalMux
    port map (
            O => \N__11933\,
            I => \N__11930\
        );

    \I__2843\ : Span12Mux_h
    port map (
            O => \N__11930\,
            I => \N__11927\
        );

    \I__2842\ : Odrv12
    port map (
            O => \N__11927\,
            I => mem_out_bus3_7
        );

    \I__2841\ : InMux
    port map (
            O => \N__11924\,
            I => \N__11921\
        );

    \I__2840\ : LocalMux
    port map (
            O => \N__11921\,
            I => \N__11918\
        );

    \I__2839\ : Sp12to4
    port map (
            O => \N__11918\,
            I => \N__11915\
        );

    \I__2838\ : Span12Mux_v
    port map (
            O => \N__11915\,
            I => \N__11912\
        );

    \I__2837\ : Odrv12
    port map (
            O => \N__11912\,
            I => \dout_obuf_RNO_3Z0Z_7\
        );

    \I__2836\ : InMux
    port map (
            O => \N__11909\,
            I => \N__11906\
        );

    \I__2835\ : LocalMux
    port map (
            O => \N__11906\,
            I => \N__11903\
        );

    \I__2834\ : Span4Mux_h
    port map (
            O => \N__11903\,
            I => \N__11900\
        );

    \I__2833\ : Odrv4
    port map (
            O => \N__11900\,
            I => mem_out_bus7_6
        );

    \I__2832\ : InMux
    port map (
            O => \N__11897\,
            I => \N__11894\
        );

    \I__2831\ : LocalMux
    port map (
            O => \N__11894\,
            I => \N__11891\
        );

    \I__2830\ : Span4Mux_v
    port map (
            O => \N__11891\,
            I => \N__11888\
        );

    \I__2829\ : Sp12to4
    port map (
            O => \N__11888\,
            I => \N__11885\
        );

    \I__2828\ : Span12Mux_h
    port map (
            O => \N__11885\,
            I => \N__11882\
        );

    \I__2827\ : Odrv12
    port map (
            O => \N__11882\,
            I => mem_out_bus3_6
        );

    \I__2826\ : InMux
    port map (
            O => \N__11879\,
            I => \N__11876\
        );

    \I__2825\ : LocalMux
    port map (
            O => \N__11876\,
            I => \N__11873\
        );

    \I__2824\ : Sp12to4
    port map (
            O => \N__11873\,
            I => \N__11870\
        );

    \I__2823\ : Span12Mux_v
    port map (
            O => \N__11870\,
            I => \N__11867\
        );

    \I__2822\ : Span12Mux_v
    port map (
            O => \N__11867\,
            I => \N__11864\
        );

    \I__2821\ : Odrv12
    port map (
            O => \N__11864\,
            I => \dout_obuf_RNO_3Z0Z_6\
        );

    \I__2820\ : InMux
    port map (
            O => \N__11861\,
            I => \N__11858\
        );

    \I__2819\ : LocalMux
    port map (
            O => \N__11858\,
            I => \N__11855\
        );

    \I__2818\ : Span12Mux_h
    port map (
            O => \N__11855\,
            I => \N__11852\
        );

    \I__2817\ : Odrv12
    port map (
            O => \N__11852\,
            I => \dout_obuf_RNO_4Z0Z_5\
        );

    \I__2816\ : InMux
    port map (
            O => \N__11849\,
            I => \N__11846\
        );

    \I__2815\ : LocalMux
    port map (
            O => \N__11846\,
            I => \N__11843\
        );

    \I__2814\ : Span12Mux_h
    port map (
            O => \N__11843\,
            I => \N__11840\
        );

    \I__2813\ : Odrv12
    port map (
            O => \N__11840\,
            I => mem_out_bus1_5
        );

    \I__2812\ : InMux
    port map (
            O => \N__11837\,
            I => \N__11834\
        );

    \I__2811\ : LocalMux
    port map (
            O => \N__11834\,
            I => \N__11831\
        );

    \I__2810\ : Odrv12
    port map (
            O => \N__11831\,
            I => mem_out_bus5_5
        );

    \I__2809\ : InMux
    port map (
            O => \N__11828\,
            I => \N__11825\
        );

    \I__2808\ : LocalMux
    port map (
            O => \N__11825\,
            I => \mem_N_174\
        );

    \I__2807\ : CascadeMux
    port map (
            O => \N__11822\,
            I => \mem_N_172_cascade_\
        );

    \I__2806\ : IoInMux
    port map (
            O => \N__11819\,
            I => \N__11816\
        );

    \I__2805\ : LocalMux
    port map (
            O => \N__11816\,
            I => \N__11813\
        );

    \I__2804\ : Span12Mux_s8_h
    port map (
            O => \N__11813\,
            I => \N__11810\
        );

    \I__2803\ : Odrv12
    port map (
            O => \N__11810\,
            I => dout_c_3
        );

    \I__2802\ : InMux
    port map (
            O => \N__11807\,
            I => \N__11804\
        );

    \I__2801\ : LocalMux
    port map (
            O => \N__11804\,
            I => \N__11801\
        );

    \I__2800\ : Span12Mux_v
    port map (
            O => \N__11801\,
            I => \N__11798\
        );

    \I__2799\ : Odrv12
    port map (
            O => \N__11798\,
            I => \dout_obuf_RNO_4Z0Z_2\
        );

    \I__2798\ : InMux
    port map (
            O => \N__11795\,
            I => \N__11792\
        );

    \I__2797\ : LocalMux
    port map (
            O => \N__11792\,
            I => \mem_N_168\
        );

    \I__2796\ : InMux
    port map (
            O => \N__11789\,
            I => \N__11786\
        );

    \I__2795\ : LocalMux
    port map (
            O => \N__11786\,
            I => \N__11783\
        );

    \I__2794\ : Span4Mux_v
    port map (
            O => \N__11783\,
            I => \N__11780\
        );

    \I__2793\ : Sp12to4
    port map (
            O => \N__11780\,
            I => \N__11777\
        );

    \I__2792\ : Span12Mux_h
    port map (
            O => \N__11777\,
            I => \N__11774\
        );

    \I__2791\ : Odrv12
    port map (
            O => \N__11774\,
            I => mem_out_bus1_4
        );

    \I__2790\ : InMux
    port map (
            O => \N__11771\,
            I => \N__11768\
        );

    \I__2789\ : LocalMux
    port map (
            O => \N__11768\,
            I => \N__11765\
        );

    \I__2788\ : Span4Mux_v
    port map (
            O => \N__11765\,
            I => \N__11762\
        );

    \I__2787\ : Odrv4
    port map (
            O => \N__11762\,
            I => mem_out_bus5_4
        );

    \I__2786\ : CascadeMux
    port map (
            O => \N__11759\,
            I => \dout_obuf_RNO_2Z0Z_4_cascade_\
        );

    \I__2785\ : InMux
    port map (
            O => \N__11756\,
            I => \N__11753\
        );

    \I__2784\ : LocalMux
    port map (
            O => \N__11753\,
            I => \N__11750\
        );

    \I__2783\ : Span4Mux_v
    port map (
            O => \N__11750\,
            I => \N__11747\
        );

    \I__2782\ : Odrv4
    port map (
            O => \N__11747\,
            I => \mem_N_178\
        );

    \I__2781\ : InMux
    port map (
            O => \N__11744\,
            I => \N__11741\
        );

    \I__2780\ : LocalMux
    port map (
            O => \N__11741\,
            I => \N__11738\
        );

    \I__2779\ : Span4Mux_v
    port map (
            O => \N__11738\,
            I => \N__11735\
        );

    \I__2778\ : Sp12to4
    port map (
            O => \N__11735\,
            I => \N__11732\
        );

    \I__2777\ : Span12Mux_h
    port map (
            O => \N__11732\,
            I => \N__11729\
        );

    \I__2776\ : Odrv12
    port map (
            O => \N__11729\,
            I => mem_out_bus1_6
        );

    \I__2775\ : InMux
    port map (
            O => \N__11726\,
            I => \N__11723\
        );

    \I__2774\ : LocalMux
    port map (
            O => \N__11723\,
            I => \N__11720\
        );

    \I__2773\ : Span4Mux_v
    port map (
            O => \N__11720\,
            I => \N__11717\
        );

    \I__2772\ : Odrv4
    port map (
            O => \N__11717\,
            I => mem_out_bus5_6
        );

    \I__2771\ : CascadeMux
    port map (
            O => \N__11714\,
            I => \dout_obuf_RNO_2Z0Z_6_cascade_\
        );

    \I__2770\ : InMux
    port map (
            O => \N__11711\,
            I => \N__11708\
        );

    \I__2769\ : LocalMux
    port map (
            O => \N__11708\,
            I => \N__11705\
        );

    \I__2768\ : Span4Mux_v
    port map (
            O => \N__11705\,
            I => \N__11702\
        );

    \I__2767\ : Odrv4
    port map (
            O => \N__11702\,
            I => \mem_N_144\
        );

    \I__2766\ : InMux
    port map (
            O => \N__11699\,
            I => \N__11696\
        );

    \I__2765\ : LocalMux
    port map (
            O => \N__11696\,
            I => \N__11693\
        );

    \I__2764\ : Span4Mux_v
    port map (
            O => \N__11693\,
            I => \N__11690\
        );

    \I__2763\ : Odrv4
    port map (
            O => \N__11690\,
            I => mem_out_bus6_4
        );

    \I__2762\ : InMux
    port map (
            O => \N__11687\,
            I => \N__11684\
        );

    \I__2761\ : LocalMux
    port map (
            O => \N__11684\,
            I => \N__11681\
        );

    \I__2760\ : Span4Mux_v
    port map (
            O => \N__11681\,
            I => \N__11678\
        );

    \I__2759\ : Sp12to4
    port map (
            O => \N__11678\,
            I => \N__11675\
        );

    \I__2758\ : Span12Mux_h
    port map (
            O => \N__11675\,
            I => \N__11672\
        );

    \I__2757\ : Odrv12
    port map (
            O => \N__11672\,
            I => mem_out_bus2_4
        );

    \I__2756\ : InMux
    port map (
            O => \N__11669\,
            I => \N__11666\
        );

    \I__2755\ : LocalMux
    port map (
            O => \N__11666\,
            I => \N__11663\
        );

    \I__2754\ : Span12Mux_v
    port map (
            O => \N__11663\,
            I => \N__11660\
        );

    \I__2753\ : Odrv12
    port map (
            O => \N__11660\,
            I => \dout_obuf_RNO_5Z0Z_4\
        );

    \I__2752\ : InMux
    port map (
            O => \N__11657\,
            I => \N__11654\
        );

    \I__2751\ : LocalMux
    port map (
            O => \N__11654\,
            I => \N__11651\
        );

    \I__2750\ : Span4Mux_v
    port map (
            O => \N__11651\,
            I => \N__11648\
        );

    \I__2749\ : Sp12to4
    port map (
            O => \N__11648\,
            I => \N__11645\
        );

    \I__2748\ : Span12Mux_h
    port map (
            O => \N__11645\,
            I => \N__11642\
        );

    \I__2747\ : Odrv12
    port map (
            O => \N__11642\,
            I => mem_out_bus2_2
        );

    \I__2746\ : InMux
    port map (
            O => \N__11639\,
            I => \N__11636\
        );

    \I__2745\ : LocalMux
    port map (
            O => \N__11636\,
            I => \N__11633\
        );

    \I__2744\ : Span4Mux_v
    port map (
            O => \N__11633\,
            I => \N__11630\
        );

    \I__2743\ : Odrv4
    port map (
            O => \N__11630\,
            I => mem_out_bus6_2
        );

    \I__2742\ : InMux
    port map (
            O => \N__11627\,
            I => \N__11624\
        );

    \I__2741\ : LocalMux
    port map (
            O => \N__11624\,
            I => \N__11621\
        );

    \I__2740\ : Odrv12
    port map (
            O => \N__11621\,
            I => \dout_obuf_RNO_5Z0Z_2\
        );

    \I__2739\ : InMux
    port map (
            O => \N__11618\,
            I => \N__11615\
        );

    \I__2738\ : LocalMux
    port map (
            O => \N__11615\,
            I => \N__11612\
        );

    \I__2737\ : Odrv4
    port map (
            O => \N__11612\,
            I => mem_out_bus4_5
        );

    \I__2736\ : InMux
    port map (
            O => \N__11609\,
            I => \N__11606\
        );

    \I__2735\ : LocalMux
    port map (
            O => \N__11606\,
            I => \N__11603\
        );

    \I__2734\ : Span12Mux_h
    port map (
            O => \N__11603\,
            I => \N__11600\
        );

    \I__2733\ : Odrv12
    port map (
            O => \N__11600\,
            I => mem_out_bus0_5
        );

    \I__2732\ : InMux
    port map (
            O => \N__11597\,
            I => \N__11594\
        );

    \I__2731\ : LocalMux
    port map (
            O => \N__11594\,
            I => \N__11591\
        );

    \I__2730\ : Span4Mux_v
    port map (
            O => \N__11591\,
            I => \N__11588\
        );

    \I__2729\ : Sp12to4
    port map (
            O => \N__11588\,
            I => \N__11585\
        );

    \I__2728\ : Span12Mux_h
    port map (
            O => \N__11585\,
            I => \N__11582\
        );

    \I__2727\ : Odrv12
    port map (
            O => \N__11582\,
            I => mem_out_bus0_4
        );

    \I__2726\ : InMux
    port map (
            O => \N__11579\,
            I => \N__11576\
        );

    \I__2725\ : LocalMux
    port map (
            O => \N__11576\,
            I => \N__11573\
        );

    \I__2724\ : Span4Mux_v
    port map (
            O => \N__11573\,
            I => \N__11570\
        );

    \I__2723\ : Odrv4
    port map (
            O => \N__11570\,
            I => mem_out_bus4_4
        );

    \I__2722\ : InMux
    port map (
            O => \N__11567\,
            I => \N__11564\
        );

    \I__2721\ : LocalMux
    port map (
            O => \N__11564\,
            I => \N__11561\
        );

    \I__2720\ : Span4Mux_v
    port map (
            O => \N__11561\,
            I => \N__11558\
        );

    \I__2719\ : Odrv4
    port map (
            O => \N__11558\,
            I => \dout_obuf_RNO_4Z0Z_4\
        );

    \I__2718\ : CascadeMux
    port map (
            O => \N__11555\,
            I => \mem_N_180_cascade_\
        );

    \I__2717\ : IoInMux
    port map (
            O => \N__11552\,
            I => \N__11549\
        );

    \I__2716\ : LocalMux
    port map (
            O => \N__11549\,
            I => \N__11546\
        );

    \I__2715\ : Span4Mux_s2_h
    port map (
            O => \N__11546\,
            I => \N__11543\
        );

    \I__2714\ : Span4Mux_h
    port map (
            O => \N__11543\,
            I => \N__11540\
        );

    \I__2713\ : Span4Mux_h
    port map (
            O => \N__11540\,
            I => \N__11537\
        );

    \I__2712\ : Odrv4
    port map (
            O => \N__11537\,
            I => dout_c_4
        );

    \I__2711\ : InMux
    port map (
            O => \N__11534\,
            I => \N__11531\
        );

    \I__2710\ : LocalMux
    port map (
            O => \N__11531\,
            I => \N__11528\
        );

    \I__2709\ : Odrv4
    port map (
            O => \N__11528\,
            I => \dout_obuf_RNO_4Z0Z_6\
        );

    \I__2708\ : CascadeMux
    port map (
            O => \N__11525\,
            I => \mem_N_145_cascade_\
        );

    \I__2707\ : IoInMux
    port map (
            O => \N__11522\,
            I => \N__11519\
        );

    \I__2706\ : LocalMux
    port map (
            O => \N__11519\,
            I => \N__11516\
        );

    \I__2705\ : Span4Mux_s2_h
    port map (
            O => \N__11516\,
            I => \N__11513\
        );

    \I__2704\ : Span4Mux_h
    port map (
            O => \N__11513\,
            I => \N__11510\
        );

    \I__2703\ : Span4Mux_h
    port map (
            O => \N__11510\,
            I => \N__11507\
        );

    \I__2702\ : Odrv4
    port map (
            O => \N__11507\,
            I => dout_c_6
        );

    \I__2701\ : InMux
    port map (
            O => \N__11504\,
            I => \N__11501\
        );

    \I__2700\ : LocalMux
    port map (
            O => \N__11501\,
            I => \N__11498\
        );

    \I__2699\ : Sp12to4
    port map (
            O => \N__11498\,
            I => \N__11495\
        );

    \I__2698\ : Odrv12
    port map (
            O => \N__11495\,
            I => \dout_obuf_RNO_4Z0Z_3\
        );

    \I__2697\ : InMux
    port map (
            O => \N__11492\,
            I => \N__11489\
        );

    \I__2696\ : LocalMux
    port map (
            O => \N__11489\,
            I => \N__11486\
        );

    \I__2695\ : Span4Mux_v
    port map (
            O => \N__11486\,
            I => \N__11483\
        );

    \I__2694\ : Odrv4
    port map (
            O => \N__11483\,
            I => \dout_obuf_RNO_5Z0Z_3\
        );

    \I__2693\ : InMux
    port map (
            O => \N__11480\,
            I => \N__11477\
        );

    \I__2692\ : LocalMux
    port map (
            O => \N__11477\,
            I => \N__11474\
        );

    \I__2691\ : Odrv4
    port map (
            O => \N__11474\,
            I => mem_out_bus5_3
        );

    \I__2690\ : InMux
    port map (
            O => \N__11471\,
            I => \N__11468\
        );

    \I__2689\ : LocalMux
    port map (
            O => \N__11468\,
            I => \N__11465\
        );

    \I__2688\ : Span12Mux_h
    port map (
            O => \N__11465\,
            I => \N__11462\
        );

    \I__2687\ : Span12Mux_h
    port map (
            O => \N__11462\,
            I => \N__11459\
        );

    \I__2686\ : Odrv12
    port map (
            O => \N__11459\,
            I => mem_out_bus1_3
        );

    \I__2685\ : InMux
    port map (
            O => \N__11456\,
            I => \N__11453\
        );

    \I__2684\ : LocalMux
    port map (
            O => \N__11453\,
            I => \N__11450\
        );

    \I__2683\ : Span12Mux_v
    port map (
            O => \N__11450\,
            I => \N__11447\
        );

    \I__2682\ : Span12Mux_v
    port map (
            O => \N__11447\,
            I => \N__11444\
        );

    \I__2681\ : Odrv12
    port map (
            O => \N__11444\,
            I => \dout_obuf_RNO_3Z0Z_3\
        );

    \I__2680\ : CascadeMux
    port map (
            O => \N__11441\,
            I => \dout_obuf_RNO_2Z0Z_3_cascade_\
        );

    \I__2679\ : InMux
    port map (
            O => \N__11438\,
            I => \N__11435\
        );

    \I__2678\ : LocalMux
    port map (
            O => \N__11435\,
            I => \N__11432\
        );

    \I__2677\ : Span12Mux_h
    port map (
            O => \N__11432\,
            I => \N__11429\
        );

    \I__2676\ : Span12Mux_h
    port map (
            O => \N__11429\,
            I => \N__11426\
        );

    \I__2675\ : Odrv12
    port map (
            O => \N__11426\,
            I => mem_out_bus2_1
        );

    \I__2674\ : InMux
    port map (
            O => \N__11423\,
            I => \N__11420\
        );

    \I__2673\ : LocalMux
    port map (
            O => \N__11420\,
            I => \N__11417\
        );

    \I__2672\ : Odrv12
    port map (
            O => \N__11417\,
            I => mem_out_bus6_1
        );

    \I__2671\ : InMux
    port map (
            O => \N__11414\,
            I => \N__11411\
        );

    \I__2670\ : LocalMux
    port map (
            O => \N__11411\,
            I => \N__11408\
        );

    \I__2669\ : Span4Mux_v
    port map (
            O => \N__11408\,
            I => \N__11405\
        );

    \I__2668\ : Odrv4
    port map (
            O => \N__11405\,
            I => \dout_obuf_RNO_5Z0Z_1\
        );

    \I__2667\ : InMux
    port map (
            O => \N__11402\,
            I => \N__11399\
        );

    \I__2666\ : LocalMux
    port map (
            O => \N__11399\,
            I => \N__11396\
        );

    \I__2665\ : Span4Mux_h
    port map (
            O => \N__11396\,
            I => \N__11393\
        );

    \I__2664\ : Odrv4
    port map (
            O => \N__11393\,
            I => mem_out_bus6_0
        );

    \I__2663\ : InMux
    port map (
            O => \N__11390\,
            I => \N__11387\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__11387\,
            I => \N__11384\
        );

    \I__2661\ : Span4Mux_v
    port map (
            O => \N__11384\,
            I => \N__11381\
        );

    \I__2660\ : Sp12to4
    port map (
            O => \N__11381\,
            I => \N__11378\
        );

    \I__2659\ : Span12Mux_h
    port map (
            O => \N__11378\,
            I => \N__11375\
        );

    \I__2658\ : Odrv12
    port map (
            O => \N__11375\,
            I => mem_out_bus2_0
        );

    \I__2657\ : InMux
    port map (
            O => \N__11372\,
            I => \N__11369\
        );

    \I__2656\ : LocalMux
    port map (
            O => \N__11369\,
            I => \N__11366\
        );

    \I__2655\ : Odrv12
    port map (
            O => \N__11366\,
            I => \dout_obuf_RNO_5Z0Z_0\
        );

    \I__2654\ : InMux
    port map (
            O => \N__11363\,
            I => \N__11360\
        );

    \I__2653\ : LocalMux
    port map (
            O => \N__11360\,
            I => \N__11357\
        );

    \I__2652\ : Span4Mux_v
    port map (
            O => \N__11357\,
            I => \N__11354\
        );

    \I__2651\ : Odrv4
    port map (
            O => \N__11354\,
            I => mem_out_bus6_3
        );

    \I__2650\ : InMux
    port map (
            O => \N__11351\,
            I => \N__11348\
        );

    \I__2649\ : LocalMux
    port map (
            O => \N__11348\,
            I => \N__11345\
        );

    \I__2648\ : Span4Mux_v
    port map (
            O => \N__11345\,
            I => \N__11342\
        );

    \I__2647\ : Sp12to4
    port map (
            O => \N__11342\,
            I => \N__11339\
        );

    \I__2646\ : Span12Mux_h
    port map (
            O => \N__11339\,
            I => \N__11336\
        );

    \I__2645\ : Odrv12
    port map (
            O => \N__11336\,
            I => mem_out_bus2_3
        );

    \I__2644\ : InMux
    port map (
            O => \N__11333\,
            I => \N__11330\
        );

    \I__2643\ : LocalMux
    port map (
            O => \N__11330\,
            I => \N__11327\
        );

    \I__2642\ : Span4Mux_h
    port map (
            O => \N__11327\,
            I => \N__11324\
        );

    \I__2641\ : Odrv4
    port map (
            O => \N__11324\,
            I => mem_out_bus7_0
        );

    \I__2640\ : InMux
    port map (
            O => \N__11321\,
            I => \N__11318\
        );

    \I__2639\ : LocalMux
    port map (
            O => \N__11318\,
            I => \N__11315\
        );

    \I__2638\ : Span4Mux_v
    port map (
            O => \N__11315\,
            I => \N__11312\
        );

    \I__2637\ : Sp12to4
    port map (
            O => \N__11312\,
            I => \N__11309\
        );

    \I__2636\ : Span12Mux_h
    port map (
            O => \N__11309\,
            I => \N__11306\
        );

    \I__2635\ : Odrv12
    port map (
            O => \N__11306\,
            I => mem_out_bus3_0
        );

    \I__2634\ : InMux
    port map (
            O => \N__11303\,
            I => \N__11300\
        );

    \I__2633\ : LocalMux
    port map (
            O => \N__11300\,
            I => \N__11297\
        );

    \I__2632\ : Span12Mux_v
    port map (
            O => \N__11297\,
            I => \N__11294\
        );

    \I__2631\ : Odrv12
    port map (
            O => \N__11294\,
            I => \dout_obuf_RNO_3Z0Z_0\
        );

    \I__2630\ : InMux
    port map (
            O => \N__11291\,
            I => \N__11288\
        );

    \I__2629\ : LocalMux
    port map (
            O => \N__11288\,
            I => \N__11285\
        );

    \I__2628\ : Span4Mux_h
    port map (
            O => \N__11285\,
            I => \N__11282\
        );

    \I__2627\ : Odrv4
    port map (
            O => \N__11282\,
            I => mem_out_bus7_2
        );

    \I__2626\ : InMux
    port map (
            O => \N__11279\,
            I => \N__11276\
        );

    \I__2625\ : LocalMux
    port map (
            O => \N__11276\,
            I => \N__11273\
        );

    \I__2624\ : Span4Mux_v
    port map (
            O => \N__11273\,
            I => \N__11270\
        );

    \I__2623\ : Sp12to4
    port map (
            O => \N__11270\,
            I => \N__11267\
        );

    \I__2622\ : Span12Mux_h
    port map (
            O => \N__11267\,
            I => \N__11264\
        );

    \I__2621\ : Odrv12
    port map (
            O => \N__11264\,
            I => mem_out_bus3_2
        );

    \I__2620\ : InMux
    port map (
            O => \N__11261\,
            I => \N__11258\
        );

    \I__2619\ : LocalMux
    port map (
            O => \N__11258\,
            I => \N__11255\
        );

    \I__2618\ : Span12Mux_v
    port map (
            O => \N__11255\,
            I => \N__11252\
        );

    \I__2617\ : Span12Mux_v
    port map (
            O => \N__11252\,
            I => \N__11249\
        );

    \I__2616\ : Odrv12
    port map (
            O => \N__11249\,
            I => \dout_obuf_RNO_3Z0Z_2\
        );

    \I__2615\ : InMux
    port map (
            O => \N__11246\,
            I => \N__11243\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__11243\,
            I => \N__11240\
        );

    \I__2613\ : Odrv4
    port map (
            O => \N__11240\,
            I => mem_out_bus7_3
        );

    \I__2612\ : InMux
    port map (
            O => \N__11237\,
            I => \N__11234\
        );

    \I__2611\ : LocalMux
    port map (
            O => \N__11234\,
            I => \N__11231\
        );

    \I__2610\ : Span12Mux_h
    port map (
            O => \N__11231\,
            I => \N__11228\
        );

    \I__2609\ : Span12Mux_h
    port map (
            O => \N__11228\,
            I => \N__11225\
        );

    \I__2608\ : Odrv12
    port map (
            O => \N__11225\,
            I => mem_out_bus3_3
        );

    \I__2607\ : InMux
    port map (
            O => \N__11222\,
            I => \N__11219\
        );

    \I__2606\ : LocalMux
    port map (
            O => \N__11219\,
            I => \N__11216\
        );

    \I__2605\ : Span4Mux_s3_v
    port map (
            O => \N__11216\,
            I => \N__11213\
        );

    \I__2604\ : Odrv4
    port map (
            O => \N__11213\,
            I => mem_out_bus4_2
        );

    \I__2603\ : InMux
    port map (
            O => \N__11210\,
            I => \N__11207\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__11207\,
            I => \N__11204\
        );

    \I__2601\ : Span4Mux_s3_v
    port map (
            O => \N__11204\,
            I => \N__11201\
        );

    \I__2600\ : Sp12to4
    port map (
            O => \N__11201\,
            I => \N__11198\
        );

    \I__2599\ : Span12Mux_h
    port map (
            O => \N__11198\,
            I => \N__11195\
        );

    \I__2598\ : Odrv12
    port map (
            O => \N__11195\,
            I => mem_out_bus0_2
        );

    \I__2597\ : InMux
    port map (
            O => \N__11192\,
            I => \N__11189\
        );

    \I__2596\ : LocalMux
    port map (
            O => \N__11189\,
            I => \N__11186\
        );

    \I__2595\ : Odrv4
    port map (
            O => \N__11186\,
            I => mem_out_bus4_3
        );

    \I__2594\ : InMux
    port map (
            O => \N__11183\,
            I => \N__11180\
        );

    \I__2593\ : LocalMux
    port map (
            O => \N__11180\,
            I => \N__11177\
        );

    \I__2592\ : Span12Mux_h
    port map (
            O => \N__11177\,
            I => \N__11174\
        );

    \I__2591\ : Odrv12
    port map (
            O => \N__11174\,
            I => mem_out_bus0_3
        );

    \I__2590\ : InMux
    port map (
            O => \N__11171\,
            I => \N__11168\
        );

    \I__2589\ : LocalMux
    port map (
            O => \N__11168\,
            I => \N__11165\
        );

    \I__2588\ : Odrv12
    port map (
            O => \N__11165\,
            I => \dout_obuf_RNO_2Z0Z_1\
        );

    \I__2587\ : InMux
    port map (
            O => \N__11162\,
            I => \N__11159\
        );

    \I__2586\ : LocalMux
    port map (
            O => \N__11159\,
            I => \mem_N_160\
        );

    \I__2585\ : InMux
    port map (
            O => \N__11156\,
            I => \N__11153\
        );

    \I__2584\ : LocalMux
    port map (
            O => \N__11153\,
            I => \N__11150\
        );

    \I__2583\ : Odrv4
    port map (
            O => \N__11150\,
            I => \dout_obuf_RNO_2Z0Z_0\
        );

    \I__2582\ : InMux
    port map (
            O => \N__11147\,
            I => \N__11144\
        );

    \I__2581\ : LocalMux
    port map (
            O => \N__11144\,
            I => \mem_N_154\
        );

    \I__2580\ : InMux
    port map (
            O => \N__11141\,
            I => \N__11138\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__11138\,
            I => \N__11135\
        );

    \I__2578\ : Span4Mux_h
    port map (
            O => \N__11135\,
            I => \N__11132\
        );

    \I__2577\ : Odrv4
    port map (
            O => \N__11132\,
            I => mem_out_bus5_2
        );

    \I__2576\ : InMux
    port map (
            O => \N__11129\,
            I => \N__11126\
        );

    \I__2575\ : LocalMux
    port map (
            O => \N__11126\,
            I => \N__11123\
        );

    \I__2574\ : Span4Mux_v
    port map (
            O => \N__11123\,
            I => \N__11120\
        );

    \I__2573\ : Sp12to4
    port map (
            O => \N__11120\,
            I => \N__11117\
        );

    \I__2572\ : Span12Mux_h
    port map (
            O => \N__11117\,
            I => \N__11114\
        );

    \I__2571\ : Odrv12
    port map (
            O => \N__11114\,
            I => mem_out_bus1_2
        );

    \I__2570\ : InMux
    port map (
            O => \N__11111\,
            I => \N__11108\
        );

    \I__2569\ : LocalMux
    port map (
            O => \N__11108\,
            I => \dout_obuf_RNO_2Z0Z_2\
        );

    \I__2568\ : CascadeMux
    port map (
            O => \N__11105\,
            I => \mem_N_166_cascade_\
        );

    \I__2567\ : IoInMux
    port map (
            O => \N__11102\,
            I => \N__11099\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__11099\,
            I => \N__11096\
        );

    \I__2565\ : Odrv12
    port map (
            O => \N__11096\,
            I => dout_c_2
        );

    \I__2564\ : InMux
    port map (
            O => \N__11093\,
            I => \N__11090\
        );

    \I__2563\ : LocalMux
    port map (
            O => \N__11090\,
            I => \N__11087\
        );

    \I__2562\ : Odrv12
    port map (
            O => \N__11087\,
            I => \dout_obuf_RNO_4Z0Z_7\
        );

    \I__2561\ : InMux
    port map (
            O => \N__11084\,
            I => \N__11081\
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__11081\,
            I => \N__11078\
        );

    \I__2559\ : Odrv4
    port map (
            O => \N__11078\,
            I => mem_out_bus5_7
        );

    \I__2558\ : InMux
    port map (
            O => \N__11075\,
            I => \N__11072\
        );

    \I__2557\ : LocalMux
    port map (
            O => \N__11072\,
            I => \N__11069\
        );

    \I__2556\ : Span12Mux_h
    port map (
            O => \N__11069\,
            I => \N__11066\
        );

    \I__2555\ : Span12Mux_h
    port map (
            O => \N__11066\,
            I => \N__11063\
        );

    \I__2554\ : Odrv12
    port map (
            O => \N__11063\,
            I => mem_out_bus1_7
        );

    \I__2553\ : CascadeMux
    port map (
            O => \N__11060\,
            I => \dout_obuf_RNO_2Z0Z_7_cascade_\
        );

    \I__2552\ : InMux
    port map (
            O => \N__11057\,
            I => \N__11054\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__11054\,
            I => \mem_N_150\
        );

    \I__2550\ : CascadeMux
    port map (
            O => \N__11051\,
            I => \mem_N_149_cascade_\
        );

    \I__2549\ : IoInMux
    port map (
            O => \N__11048\,
            I => \N__11045\
        );

    \I__2548\ : LocalMux
    port map (
            O => \N__11045\,
            I => \N__11042\
        );

    \I__2547\ : IoSpan4Mux
    port map (
            O => \N__11042\,
            I => \N__11039\
        );

    \I__2546\ : Span4Mux_s3_h
    port map (
            O => \N__11039\,
            I => \N__11036\
        );

    \I__2545\ : Span4Mux_h
    port map (
            O => \N__11036\,
            I => \N__11033\
        );

    \I__2544\ : Odrv4
    port map (
            O => \N__11033\,
            I => dout_c_7
        );

    \I__2543\ : InMux
    port map (
            O => \N__11030\,
            I => \N__11027\
        );

    \I__2542\ : LocalMux
    port map (
            O => \N__11027\,
            I => \N__11024\
        );

    \I__2541\ : Span4Mux_v
    port map (
            O => \N__11024\,
            I => \N__11021\
        );

    \I__2540\ : Sp12to4
    port map (
            O => \N__11021\,
            I => \N__11018\
        );

    \I__2539\ : Span12Mux_h
    port map (
            O => \N__11018\,
            I => \N__11015\
        );

    \I__2538\ : Odrv12
    port map (
            O => \N__11015\,
            I => mem_out_bus0_6
        );

    \I__2537\ : InMux
    port map (
            O => \N__11012\,
            I => \N__11009\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__11009\,
            I => \N__11006\
        );

    \I__2535\ : Span4Mux_h
    port map (
            O => \N__11006\,
            I => \N__11003\
        );

    \I__2534\ : Odrv4
    port map (
            O => \N__11003\,
            I => mem_out_bus4_6
        );

    \I__2533\ : SRMux
    port map (
            O => \N__11000\,
            I => \N__10995\
        );

    \I__2532\ : SRMux
    port map (
            O => \N__10999\,
            I => \N__10992\
        );

    \I__2531\ : SRMux
    port map (
            O => \N__10998\,
            I => \N__10987\
        );

    \I__2530\ : LocalMux
    port map (
            O => \N__10995\,
            I => \N__10980\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__10992\,
            I => \N__10980\
        );

    \I__2528\ : SRMux
    port map (
            O => \N__10991\,
            I => \N__10977\
        );

    \I__2527\ : SRMux
    port map (
            O => \N__10990\,
            I => \N__10974\
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__10987\,
            I => \N__10971\
        );

    \I__2525\ : SRMux
    port map (
            O => \N__10986\,
            I => \N__10968\
        );

    \I__2524\ : SRMux
    port map (
            O => \N__10985\,
            I => \N__10965\
        );

    \I__2523\ : Span4Mux_s3_v
    port map (
            O => \N__10980\,
            I => \N__10953\
        );

    \I__2522\ : LocalMux
    port map (
            O => \N__10977\,
            I => \N__10953\
        );

    \I__2521\ : LocalMux
    port map (
            O => \N__10974\,
            I => \N__10953\
        );

    \I__2520\ : Span4Mux_s3_v
    port map (
            O => \N__10971\,
            I => \N__10946\
        );

    \I__2519\ : LocalMux
    port map (
            O => \N__10968\,
            I => \N__10946\
        );

    \I__2518\ : LocalMux
    port map (
            O => \N__10965\,
            I => \N__10946\
        );

    \I__2517\ : SRMux
    port map (
            O => \N__10964\,
            I => \N__10943\
        );

    \I__2516\ : SRMux
    port map (
            O => \N__10963\,
            I => \N__10940\
        );

    \I__2515\ : SRMux
    port map (
            O => \N__10962\,
            I => \N__10937\
        );

    \I__2514\ : SRMux
    port map (
            O => \N__10961\,
            I => \N__10934\
        );

    \I__2513\ : SRMux
    port map (
            O => \N__10960\,
            I => \N__10928\
        );

    \I__2512\ : Span4Mux_v
    port map (
            O => \N__10953\,
            I => \N__10911\
        );

    \I__2511\ : Span4Mux_v
    port map (
            O => \N__10946\,
            I => \N__10911\
        );

    \I__2510\ : LocalMux
    port map (
            O => \N__10943\,
            I => \N__10911\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__10940\,
            I => \N__10911\
        );

    \I__2508\ : LocalMux
    port map (
            O => \N__10937\,
            I => \N__10906\
        );

    \I__2507\ : LocalMux
    port map (
            O => \N__10934\,
            I => \N__10906\
        );

    \I__2506\ : SRMux
    port map (
            O => \N__10933\,
            I => \N__10903\
        );

    \I__2505\ : SRMux
    port map (
            O => \N__10932\,
            I => \N__10900\
        );

    \I__2504\ : SRMux
    port map (
            O => \N__10931\,
            I => \N__10895\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__10928\,
            I => \N__10892\
        );

    \I__2502\ : SRMux
    port map (
            O => \N__10927\,
            I => \N__10889\
        );

    \I__2501\ : SRMux
    port map (
            O => \N__10926\,
            I => \N__10886\
        );

    \I__2500\ : SRMux
    port map (
            O => \N__10925\,
            I => \N__10882\
        );

    \I__2499\ : SRMux
    port map (
            O => \N__10924\,
            I => \N__10879\
        );

    \I__2498\ : SRMux
    port map (
            O => \N__10923\,
            I => \N__10873\
        );

    \I__2497\ : SRMux
    port map (
            O => \N__10922\,
            I => \N__10870\
        );

    \I__2496\ : SRMux
    port map (
            O => \N__10921\,
            I => \N__10865\
        );

    \I__2495\ : SRMux
    port map (
            O => \N__10920\,
            I => \N__10859\
        );

    \I__2494\ : Span4Mux_v
    port map (
            O => \N__10911\,
            I => \N__10849\
        );

    \I__2493\ : Span4Mux_v
    port map (
            O => \N__10906\,
            I => \N__10849\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__10903\,
            I => \N__10849\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__10900\,
            I => \N__10849\
        );

    \I__2490\ : SRMux
    port map (
            O => \N__10899\,
            I => \N__10846\
        );

    \I__2489\ : SRMux
    port map (
            O => \N__10898\,
            I => \N__10843\
        );

    \I__2488\ : LocalMux
    port map (
            O => \N__10895\,
            I => \N__10835\
        );

    \I__2487\ : Span4Mux_s0_v
    port map (
            O => \N__10892\,
            I => \N__10835\
        );

    \I__2486\ : LocalMux
    port map (
            O => \N__10889\,
            I => \N__10835\
        );

    \I__2485\ : LocalMux
    port map (
            O => \N__10886\,
            I => \N__10832\
        );

    \I__2484\ : SRMux
    port map (
            O => \N__10885\,
            I => \N__10829\
        );

    \I__2483\ : LocalMux
    port map (
            O => \N__10882\,
            I => \N__10823\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__10879\,
            I => \N__10823\
        );

    \I__2481\ : SRMux
    port map (
            O => \N__10878\,
            I => \N__10820\
        );

    \I__2480\ : SRMux
    port map (
            O => \N__10877\,
            I => \N__10817\
        );

    \I__2479\ : SRMux
    port map (
            O => \N__10876\,
            I => \N__10813\
        );

    \I__2478\ : LocalMux
    port map (
            O => \N__10873\,
            I => \N__10808\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__10870\,
            I => \N__10805\
        );

    \I__2476\ : SRMux
    port map (
            O => \N__10869\,
            I => \N__10802\
        );

    \I__2475\ : SRMux
    port map (
            O => \N__10868\,
            I => \N__10799\
        );

    \I__2474\ : LocalMux
    port map (
            O => \N__10865\,
            I => \N__10795\
        );

    \I__2473\ : SRMux
    port map (
            O => \N__10864\,
            I => \N__10792\
        );

    \I__2472\ : SRMux
    port map (
            O => \N__10863\,
            I => \N__10789\
        );

    \I__2471\ : SRMux
    port map (
            O => \N__10862\,
            I => \N__10783\
        );

    \I__2470\ : LocalMux
    port map (
            O => \N__10859\,
            I => \N__10780\
        );

    \I__2469\ : SRMux
    port map (
            O => \N__10858\,
            I => \N__10777\
        );

    \I__2468\ : Span4Mux_v
    port map (
            O => \N__10849\,
            I => \N__10770\
        );

    \I__2467\ : LocalMux
    port map (
            O => \N__10846\,
            I => \N__10770\
        );

    \I__2466\ : LocalMux
    port map (
            O => \N__10843\,
            I => \N__10770\
        );

    \I__2465\ : SRMux
    port map (
            O => \N__10842\,
            I => \N__10767\
        );

    \I__2464\ : Span4Mux_v
    port map (
            O => \N__10835\,
            I => \N__10760\
        );

    \I__2463\ : Span4Mux_v
    port map (
            O => \N__10832\,
            I => \N__10760\
        );

    \I__2462\ : LocalMux
    port map (
            O => \N__10829\,
            I => \N__10760\
        );

    \I__2461\ : SRMux
    port map (
            O => \N__10828\,
            I => \N__10757\
        );

    \I__2460\ : Span4Mux_v
    port map (
            O => \N__10823\,
            I => \N__10750\
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__10820\,
            I => \N__10750\
        );

    \I__2458\ : LocalMux
    port map (
            O => \N__10817\,
            I => \N__10750\
        );

    \I__2457\ : SRMux
    port map (
            O => \N__10816\,
            I => \N__10747\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__10813\,
            I => \N__10744\
        );

    \I__2455\ : SRMux
    port map (
            O => \N__10812\,
            I => \N__10741\
        );

    \I__2454\ : SRMux
    port map (
            O => \N__10811\,
            I => \N__10737\
        );

    \I__2453\ : Span4Mux_s3_v
    port map (
            O => \N__10808\,
            I => \N__10727\
        );

    \I__2452\ : Span4Mux_s3_v
    port map (
            O => \N__10805\,
            I => \N__10727\
        );

    \I__2451\ : LocalMux
    port map (
            O => \N__10802\,
            I => \N__10727\
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__10799\,
            I => \N__10727\
        );

    \I__2449\ : SRMux
    port map (
            O => \N__10798\,
            I => \N__10724\
        );

    \I__2448\ : Span4Mux_s3_v
    port map (
            O => \N__10795\,
            I => \N__10717\
        );

    \I__2447\ : LocalMux
    port map (
            O => \N__10792\,
            I => \N__10717\
        );

    \I__2446\ : LocalMux
    port map (
            O => \N__10789\,
            I => \N__10717\
        );

    \I__2445\ : SRMux
    port map (
            O => \N__10788\,
            I => \N__10714\
        );

    \I__2444\ : SRMux
    port map (
            O => \N__10787\,
            I => \N__10711\
        );

    \I__2443\ : SRMux
    port map (
            O => \N__10786\,
            I => \N__10706\
        );

    \I__2442\ : LocalMux
    port map (
            O => \N__10783\,
            I => \N__10696\
        );

    \I__2441\ : Span4Mux_h
    port map (
            O => \N__10780\,
            I => \N__10696\
        );

    \I__2440\ : LocalMux
    port map (
            O => \N__10777\,
            I => \N__10696\
        );

    \I__2439\ : Span4Mux_v
    port map (
            O => \N__10770\,
            I => \N__10687\
        );

    \I__2438\ : LocalMux
    port map (
            O => \N__10767\,
            I => \N__10687\
        );

    \I__2437\ : Span4Mux_v
    port map (
            O => \N__10760\,
            I => \N__10687\
        );

    \I__2436\ : LocalMux
    port map (
            O => \N__10757\,
            I => \N__10687\
        );

    \I__2435\ : Span4Mux_v
    port map (
            O => \N__10750\,
            I => \N__10678\
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__10747\,
            I => \N__10678\
        );

    \I__2433\ : Span4Mux_h
    port map (
            O => \N__10744\,
            I => \N__10678\
        );

    \I__2432\ : LocalMux
    port map (
            O => \N__10741\,
            I => \N__10678\
        );

    \I__2431\ : SRMux
    port map (
            O => \N__10740\,
            I => \N__10675\
        );

    \I__2430\ : LocalMux
    port map (
            O => \N__10737\,
            I => \N__10672\
        );

    \I__2429\ : SRMux
    port map (
            O => \N__10736\,
            I => \N__10669\
        );

    \I__2428\ : Span4Mux_v
    port map (
            O => \N__10727\,
            I => \N__10664\
        );

    \I__2427\ : LocalMux
    port map (
            O => \N__10724\,
            I => \N__10664\
        );

    \I__2426\ : Span4Mux_v
    port map (
            O => \N__10717\,
            I => \N__10657\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__10714\,
            I => \N__10657\
        );

    \I__2424\ : LocalMux
    port map (
            O => \N__10711\,
            I => \N__10657\
        );

    \I__2423\ : SRMux
    port map (
            O => \N__10710\,
            I => \N__10654\
        );

    \I__2422\ : SRMux
    port map (
            O => \N__10709\,
            I => \N__10651\
        );

    \I__2421\ : LocalMux
    port map (
            O => \N__10706\,
            I => \N__10648\
        );

    \I__2420\ : SRMux
    port map (
            O => \N__10705\,
            I => \N__10645\
        );

    \I__2419\ : SRMux
    port map (
            O => \N__10704\,
            I => \N__10642\
        );

    \I__2418\ : SRMux
    port map (
            O => \N__10703\,
            I => \N__10633\
        );

    \I__2417\ : Span4Mux_v
    port map (
            O => \N__10696\,
            I => \N__10624\
        );

    \I__2416\ : Span4Mux_v
    port map (
            O => \N__10687\,
            I => \N__10624\
        );

    \I__2415\ : Span4Mux_v
    port map (
            O => \N__10678\,
            I => \N__10624\
        );

    \I__2414\ : LocalMux
    port map (
            O => \N__10675\,
            I => \N__10617\
        );

    \I__2413\ : Span4Mux_h
    port map (
            O => \N__10672\,
            I => \N__10617\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__10669\,
            I => \N__10617\
        );

    \I__2411\ : Span4Mux_v
    port map (
            O => \N__10664\,
            I => \N__10608\
        );

    \I__2410\ : Span4Mux_v
    port map (
            O => \N__10657\,
            I => \N__10608\
        );

    \I__2409\ : LocalMux
    port map (
            O => \N__10654\,
            I => \N__10608\
        );

    \I__2408\ : LocalMux
    port map (
            O => \N__10651\,
            I => \N__10608\
        );

    \I__2407\ : Span4Mux_v
    port map (
            O => \N__10648\,
            I => \N__10601\
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__10645\,
            I => \N__10601\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__10642\,
            I => \N__10601\
        );

    \I__2404\ : SRMux
    port map (
            O => \N__10641\,
            I => \N__10598\
        );

    \I__2403\ : SRMux
    port map (
            O => \N__10640\,
            I => \N__10595\
        );

    \I__2402\ : SRMux
    port map (
            O => \N__10639\,
            I => \N__10591\
        );

    \I__2401\ : SRMux
    port map (
            O => \N__10638\,
            I => \N__10586\
        );

    \I__2400\ : SRMux
    port map (
            O => \N__10637\,
            I => \N__10583\
        );

    \I__2399\ : SRMux
    port map (
            O => \N__10636\,
            I => \N__10579\
        );

    \I__2398\ : LocalMux
    port map (
            O => \N__10633\,
            I => \N__10576\
        );

    \I__2397\ : SRMux
    port map (
            O => \N__10632\,
            I => \N__10573\
        );

    \I__2396\ : SRMux
    port map (
            O => \N__10631\,
            I => \N__10570\
        );

    \I__2395\ : Span4Mux_h
    port map (
            O => \N__10624\,
            I => \N__10567\
        );

    \I__2394\ : Span4Mux_v
    port map (
            O => \N__10617\,
            I => \N__10564\
        );

    \I__2393\ : Span4Mux_v
    port map (
            O => \N__10608\,
            I => \N__10555\
        );

    \I__2392\ : Span4Mux_v
    port map (
            O => \N__10601\,
            I => \N__10555\
        );

    \I__2391\ : LocalMux
    port map (
            O => \N__10598\,
            I => \N__10555\
        );

    \I__2390\ : LocalMux
    port map (
            O => \N__10595\,
            I => \N__10555\
        );

    \I__2389\ : SRMux
    port map (
            O => \N__10594\,
            I => \N__10552\
        );

    \I__2388\ : LocalMux
    port map (
            O => \N__10591\,
            I => \N__10549\
        );

    \I__2387\ : SRMux
    port map (
            O => \N__10590\,
            I => \N__10546\
        );

    \I__2386\ : SRMux
    port map (
            O => \N__10589\,
            I => \N__10543\
        );

    \I__2385\ : LocalMux
    port map (
            O => \N__10586\,
            I => \N__10540\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__10583\,
            I => \N__10537\
        );

    \I__2383\ : SRMux
    port map (
            O => \N__10582\,
            I => \N__10534\
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__10579\,
            I => \N__10531\
        );

    \I__2381\ : Span4Mux_h
    port map (
            O => \N__10576\,
            I => \N__10527\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__10573\,
            I => \N__10524\
        );

    \I__2379\ : LocalMux
    port map (
            O => \N__10570\,
            I => \N__10521\
        );

    \I__2378\ : Span4Mux_h
    port map (
            O => \N__10567\,
            I => \N__10518\
        );

    \I__2377\ : Span4Mux_v
    port map (
            O => \N__10564\,
            I => \N__10513\
        );

    \I__2376\ : Span4Mux_v
    port map (
            O => \N__10555\,
            I => \N__10513\
        );

    \I__2375\ : LocalMux
    port map (
            O => \N__10552\,
            I => \N__10510\
        );

    \I__2374\ : Span4Mux_h
    port map (
            O => \N__10549\,
            I => \N__10507\
        );

    \I__2373\ : LocalMux
    port map (
            O => \N__10546\,
            I => \N__10504\
        );

    \I__2372\ : LocalMux
    port map (
            O => \N__10543\,
            I => \N__10501\
        );

    \I__2371\ : Span4Mux_h
    port map (
            O => \N__10540\,
            I => \N__10496\
        );

    \I__2370\ : Span4Mux_h
    port map (
            O => \N__10537\,
            I => \N__10496\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__10534\,
            I => \N__10493\
        );

    \I__2368\ : Span4Mux_h
    port map (
            O => \N__10531\,
            I => \N__10490\
        );

    \I__2367\ : SRMux
    port map (
            O => \N__10530\,
            I => \N__10487\
        );

    \I__2366\ : Span4Mux_v
    port map (
            O => \N__10527\,
            I => \N__10480\
        );

    \I__2365\ : Span4Mux_h
    port map (
            O => \N__10524\,
            I => \N__10480\
        );

    \I__2364\ : Span4Mux_h
    port map (
            O => \N__10521\,
            I => \N__10480\
        );

    \I__2363\ : Span4Mux_h
    port map (
            O => \N__10518\,
            I => \N__10475\
        );

    \I__2362\ : Span4Mux_v
    port map (
            O => \N__10513\,
            I => \N__10475\
        );

    \I__2361\ : Span4Mux_h
    port map (
            O => \N__10510\,
            I => \N__10472\
        );

    \I__2360\ : Span4Mux_v
    port map (
            O => \N__10507\,
            I => \N__10465\
        );

    \I__2359\ : Span4Mux_h
    port map (
            O => \N__10504\,
            I => \N__10465\
        );

    \I__2358\ : Span4Mux_h
    port map (
            O => \N__10501\,
            I => \N__10465\
        );

    \I__2357\ : Sp12to4
    port map (
            O => \N__10496\,
            I => \N__10460\
        );

    \I__2356\ : Span12Mux_s9_h
    port map (
            O => \N__10493\,
            I => \N__10460\
        );

    \I__2355\ : Span4Mux_v
    port map (
            O => \N__10490\,
            I => \N__10455\
        );

    \I__2354\ : LocalMux
    port map (
            O => \N__10487\,
            I => \N__10455\
        );

    \I__2353\ : Span4Mux_v
    port map (
            O => \N__10480\,
            I => \N__10452\
        );

    \I__2352\ : Odrv4
    port map (
            O => \N__10475\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2351\ : Odrv4
    port map (
            O => \N__10472\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2350\ : Odrv4
    port map (
            O => \N__10465\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2349\ : Odrv12
    port map (
            O => \N__10460\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2348\ : Odrv4
    port map (
            O => \N__10455\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2347\ : Odrv4
    port map (
            O => \N__10452\,
            I => \CONSTANT_ONE_NET\
        );

    \I__2346\ : InMux
    port map (
            O => \N__10439\,
            I => \N__10436\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__10436\,
            I => \N__10433\
        );

    \I__2344\ : Odrv4
    port map (
            O => \N__10433\,
            I => mem_out_bus5_1
        );

    \I__2343\ : InMux
    port map (
            O => \N__10430\,
            I => \N__10427\
        );

    \I__2342\ : LocalMux
    port map (
            O => \N__10427\,
            I => \N__10424\
        );

    \I__2341\ : Span12Mux_h
    port map (
            O => \N__10424\,
            I => \N__10421\
        );

    \I__2340\ : Span12Mux_h
    port map (
            O => \N__10421\,
            I => \N__10418\
        );

    \I__2339\ : Odrv12
    port map (
            O => \N__10418\,
            I => mem_out_bus1_1
        );

    \I__2338\ : InMux
    port map (
            O => \N__10415\,
            I => \N__10412\
        );

    \I__2337\ : LocalMux
    port map (
            O => \N__10412\,
            I => \N__10409\
        );

    \I__2336\ : Span4Mux_h
    port map (
            O => \N__10409\,
            I => \N__10406\
        );

    \I__2335\ : Odrv4
    port map (
            O => \N__10406\,
            I => mem_out_bus5_0
        );

    \I__2334\ : InMux
    port map (
            O => \N__10403\,
            I => \N__10400\
        );

    \I__2333\ : LocalMux
    port map (
            O => \N__10400\,
            I => \N__10397\
        );

    \I__2332\ : Span4Mux_v
    port map (
            O => \N__10397\,
            I => \N__10394\
        );

    \I__2331\ : Sp12to4
    port map (
            O => \N__10394\,
            I => \N__10391\
        );

    \I__2330\ : Span12Mux_h
    port map (
            O => \N__10391\,
            I => \N__10388\
        );

    \I__2329\ : Odrv12
    port map (
            O => \N__10388\,
            I => mem_out_bus1_0
        );

    \I__2328\ : InMux
    port map (
            O => \N__10385\,
            I => \N__10382\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__10382\,
            I => \N__10379\
        );

    \I__2326\ : Span12Mux_v
    port map (
            O => \N__10379\,
            I => \N__10376\
        );

    \I__2325\ : Odrv12
    port map (
            O => \N__10376\,
            I => \dout_obuf_RNO_4Z0Z_1\
        );

    \I__2324\ : CascadeMux
    port map (
            O => \N__10373\,
            I => \mem_N_162_cascade_\
        );

    \I__2323\ : IoInMux
    port map (
            O => \N__10370\,
            I => \N__10367\
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__10367\,
            I => \N__10364\
        );

    \I__2321\ : Span12Mux_s9_h
    port map (
            O => \N__10364\,
            I => \N__10361\
        );

    \I__2320\ : Odrv12
    port map (
            O => \N__10361\,
            I => dout_c_1
        );

    \I__2319\ : InMux
    port map (
            O => \N__10358\,
            I => \N__10355\
        );

    \I__2318\ : LocalMux
    port map (
            O => \N__10355\,
            I => \N__10352\
        );

    \I__2317\ : Span12Mux_v
    port map (
            O => \N__10352\,
            I => \N__10349\
        );

    \I__2316\ : Odrv12
    port map (
            O => \N__10349\,
            I => \dout_obuf_RNO_4Z0Z_0\
        );

    \I__2315\ : CascadeMux
    port map (
            O => \N__10346\,
            I => \mem_N_156_cascade_\
        );

    \I__2314\ : IoInMux
    port map (
            O => \N__10343\,
            I => \N__10340\
        );

    \I__2313\ : LocalMux
    port map (
            O => \N__10340\,
            I => \N__10337\
        );

    \I__2312\ : Span4Mux_s2_h
    port map (
            O => \N__10337\,
            I => \N__10334\
        );

    \I__2311\ : Sp12to4
    port map (
            O => \N__10334\,
            I => \N__10331\
        );

    \I__2310\ : Span12Mux_s10_v
    port map (
            O => \N__10331\,
            I => \N__10328\
        );

    \I__2309\ : Odrv12
    port map (
            O => \N__10328\,
            I => dout_c_0
        );

    \I__2308\ : CEMux
    port map (
            O => \N__10325\,
            I => \N__10321\
        );

    \I__2307\ : CEMux
    port map (
            O => \N__10324\,
            I => \N__10318\
        );

    \I__2306\ : LocalMux
    port map (
            O => \N__10321\,
            I => \N__10314\
        );

    \I__2305\ : LocalMux
    port map (
            O => \N__10318\,
            I => \N__10311\
        );

    \I__2304\ : CEMux
    port map (
            O => \N__10317\,
            I => \N__10308\
        );

    \I__2303\ : Span4Mux_v
    port map (
            O => \N__10314\,
            I => \N__10301\
        );

    \I__2302\ : Span4Mux_h
    port map (
            O => \N__10311\,
            I => \N__10301\
        );

    \I__2301\ : LocalMux
    port map (
            O => \N__10308\,
            I => \N__10301\
        );

    \I__2300\ : Span4Mux_v
    port map (
            O => \N__10301\,
            I => \N__10297\
        );

    \I__2299\ : CEMux
    port map (
            O => \N__10300\,
            I => \N__10294\
        );

    \I__2298\ : Odrv4
    port map (
            O => \N__10297\,
            I => \mem_WE_8\
        );

    \I__2297\ : LocalMux
    port map (
            O => \N__10294\,
            I => \mem_WE_8\
        );

    \I__2296\ : CEMux
    port map (
            O => \N__10289\,
            I => \N__10285\
        );

    \I__2295\ : CEMux
    port map (
            O => \N__10288\,
            I => \N__10282\
        );

    \I__2294\ : LocalMux
    port map (
            O => \N__10285\,
            I => \N__10276\
        );

    \I__2293\ : LocalMux
    port map (
            O => \N__10282\,
            I => \N__10276\
        );

    \I__2292\ : CEMux
    port map (
            O => \N__10281\,
            I => \N__10273\
        );

    \I__2291\ : Span4Mux_v
    port map (
            O => \N__10276\,
            I => \N__10267\
        );

    \I__2290\ : LocalMux
    port map (
            O => \N__10273\,
            I => \N__10267\
        );

    \I__2289\ : CEMux
    port map (
            O => \N__10272\,
            I => \N__10264\
        );

    \I__2288\ : Span4Mux_v
    port map (
            O => \N__10267\,
            I => \N__10261\
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__10264\,
            I => \N__10258\
        );

    \I__2286\ : Span4Mux_v
    port map (
            O => \N__10261\,
            I => \N__10255\
        );

    \I__2285\ : Span12Mux_h
    port map (
            O => \N__10258\,
            I => \N__10252\
        );

    \I__2284\ : Odrv4
    port map (
            O => \N__10255\,
            I => \mem_WE_12\
        );

    \I__2283\ : Odrv12
    port map (
            O => \N__10252\,
            I => \mem_WE_12\
        );

    \I__2282\ : CEMux
    port map (
            O => \N__10247\,
            I => \N__10243\
        );

    \I__2281\ : CEMux
    port map (
            O => \N__10246\,
            I => \N__10240\
        );

    \I__2280\ : LocalMux
    port map (
            O => \N__10243\,
            I => \N__10233\
        );

    \I__2279\ : LocalMux
    port map (
            O => \N__10240\,
            I => \N__10233\
        );

    \I__2278\ : CEMux
    port map (
            O => \N__10239\,
            I => \N__10230\
        );

    \I__2277\ : CEMux
    port map (
            O => \N__10238\,
            I => \N__10227\
        );

    \I__2276\ : Span4Mux_s3_v
    port map (
            O => \N__10233\,
            I => \N__10220\
        );

    \I__2275\ : LocalMux
    port map (
            O => \N__10230\,
            I => \N__10220\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__10227\,
            I => \N__10220\
        );

    \I__2273\ : Span4Mux_v
    port map (
            O => \N__10220\,
            I => \N__10217\
        );

    \I__2272\ : Span4Mux_v
    port map (
            O => \N__10217\,
            I => \N__10214\
        );

    \I__2271\ : Span4Mux_v
    port map (
            O => \N__10214\,
            I => \N__10211\
        );

    \I__2270\ : Sp12to4
    port map (
            O => \N__10211\,
            I => \N__10208\
        );

    \I__2269\ : Span12Mux_h
    port map (
            O => \N__10208\,
            I => \N__10205\
        );

    \I__2268\ : Odrv12
    port map (
            O => \N__10205\,
            I => \mem_WE_16\
        );

    \I__2267\ : CEMux
    port map (
            O => \N__10202\,
            I => \N__10199\
        );

    \I__2266\ : LocalMux
    port map (
            O => \N__10199\,
            I => \N__10193\
        );

    \I__2265\ : CEMux
    port map (
            O => \N__10198\,
            I => \N__10190\
        );

    \I__2264\ : CEMux
    port map (
            O => \N__10197\,
            I => \N__10187\
        );

    \I__2263\ : CEMux
    port map (
            O => \N__10196\,
            I => \N__10184\
        );

    \I__2262\ : Span4Mux_v
    port map (
            O => \N__10193\,
            I => \N__10181\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__10190\,
            I => \N__10178\
        );

    \I__2260\ : LocalMux
    port map (
            O => \N__10187\,
            I => \N__10173\
        );

    \I__2259\ : LocalMux
    port map (
            O => \N__10184\,
            I => \N__10173\
        );

    \I__2258\ : Span4Mux_h
    port map (
            O => \N__10181\,
            I => \N__10168\
        );

    \I__2257\ : Span4Mux_h
    port map (
            O => \N__10178\,
            I => \N__10168\
        );

    \I__2256\ : Span4Mux_v
    port map (
            O => \N__10173\,
            I => \N__10165\
        );

    \I__2255\ : Span4Mux_h
    port map (
            O => \N__10168\,
            I => \N__10162\
        );

    \I__2254\ : Span4Mux_h
    port map (
            O => \N__10165\,
            I => \N__10159\
        );

    \I__2253\ : Sp12to4
    port map (
            O => \N__10162\,
            I => \N__10156\
        );

    \I__2252\ : Sp12to4
    port map (
            O => \N__10159\,
            I => \N__10153\
        );

    \I__2251\ : Span12Mux_v
    port map (
            O => \N__10156\,
            I => \N__10148\
        );

    \I__2250\ : Span12Mux_h
    port map (
            O => \N__10153\,
            I => \N__10148\
        );

    \I__2249\ : Odrv12
    port map (
            O => \N__10148\,
            I => \mem_WE_20\
        );

    \I__2248\ : CEMux
    port map (
            O => \N__10145\,
            I => \N__10141\
        );

    \I__2247\ : CEMux
    port map (
            O => \N__10144\,
            I => \N__10138\
        );

    \I__2246\ : LocalMux
    port map (
            O => \N__10141\,
            I => \N__10131\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__10138\,
            I => \N__10131\
        );

    \I__2244\ : CEMux
    port map (
            O => \N__10137\,
            I => \N__10128\
        );

    \I__2243\ : CEMux
    port map (
            O => \N__10136\,
            I => \N__10125\
        );

    \I__2242\ : Span4Mux_v
    port map (
            O => \N__10131\,
            I => \N__10118\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__10128\,
            I => \N__10118\
        );

    \I__2240\ : LocalMux
    port map (
            O => \N__10125\,
            I => \N__10118\
        );

    \I__2239\ : Span4Mux_v
    port map (
            O => \N__10118\,
            I => \N__10115\
        );

    \I__2238\ : Span4Mux_h
    port map (
            O => \N__10115\,
            I => \N__10112\
        );

    \I__2237\ : Span4Mux_h
    port map (
            O => \N__10112\,
            I => \N__10109\
        );

    \I__2236\ : Span4Mux_h
    port map (
            O => \N__10109\,
            I => \N__10106\
        );

    \I__2235\ : Span4Mux_h
    port map (
            O => \N__10106\,
            I => \N__10103\
        );

    \I__2234\ : Odrv4
    port map (
            O => \N__10103\,
            I => \mem_WE_24\
        );

    \I__2233\ : InMux
    port map (
            O => \N__10100\,
            I => \N__10076\
        );

    \I__2232\ : InMux
    port map (
            O => \N__10099\,
            I => \N__10076\
        );

    \I__2231\ : InMux
    port map (
            O => \N__10098\,
            I => \N__10076\
        );

    \I__2230\ : InMux
    port map (
            O => \N__10097\,
            I => \N__10076\
        );

    \I__2229\ : InMux
    port map (
            O => \N__10096\,
            I => \N__10076\
        );

    \I__2228\ : InMux
    port map (
            O => \N__10095\,
            I => \N__10076\
        );

    \I__2227\ : InMux
    port map (
            O => \N__10094\,
            I => \N__10076\
        );

    \I__2226\ : InMux
    port map (
            O => \N__10093\,
            I => \N__10076\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__10076\,
            I => \N__10073\
        );

    \I__2224\ : Span4Mux_v
    port map (
            O => \N__10073\,
            I => \N__10070\
        );

    \I__2223\ : Span4Mux_h
    port map (
            O => \N__10070\,
            I => \N__10067\
        );

    \I__2222\ : Odrv4
    port map (
            O => \N__10067\,
            I => write_en_c
        );

    \I__2221\ : InMux
    port map (
            O => \N__10064\,
            I => \N__10040\
        );

    \I__2220\ : InMux
    port map (
            O => \N__10063\,
            I => \N__10040\
        );

    \I__2219\ : InMux
    port map (
            O => \N__10062\,
            I => \N__10040\
        );

    \I__2218\ : InMux
    port map (
            O => \N__10061\,
            I => \N__10040\
        );

    \I__2217\ : InMux
    port map (
            O => \N__10060\,
            I => \N__10040\
        );

    \I__2216\ : InMux
    port map (
            O => \N__10059\,
            I => \N__10040\
        );

    \I__2215\ : InMux
    port map (
            O => \N__10058\,
            I => \N__10040\
        );

    \I__2214\ : InMux
    port map (
            O => \N__10057\,
            I => \N__10040\
        );

    \I__2213\ : LocalMux
    port map (
            O => \N__10040\,
            I => \N__10037\
        );

    \I__2212\ : Span4Mux_v
    port map (
            O => \N__10037\,
            I => \N__10034\
        );

    \I__2211\ : Sp12to4
    port map (
            O => \N__10034\,
            I => \N__10031\
        );

    \I__2210\ : Odrv12
    port map (
            O => \N__10031\,
            I => waddr_c_13
        );

    \I__2209\ : CascadeMux
    port map (
            O => \N__10028\,
            I => \N__10022\
        );

    \I__2208\ : CascadeMux
    port map (
            O => \N__10027\,
            I => \N__10018\
        );

    \I__2207\ : CascadeMux
    port map (
            O => \N__10026\,
            I => \N__10014\
        );

    \I__2206\ : CascadeMux
    port map (
            O => \N__10025\,
            I => \N__10010\
        );

    \I__2205\ : InMux
    port map (
            O => \N__10022\,
            I => \N__9992\
        );

    \I__2204\ : InMux
    port map (
            O => \N__10021\,
            I => \N__9992\
        );

    \I__2203\ : InMux
    port map (
            O => \N__10018\,
            I => \N__9992\
        );

    \I__2202\ : InMux
    port map (
            O => \N__10017\,
            I => \N__9992\
        );

    \I__2201\ : InMux
    port map (
            O => \N__10014\,
            I => \N__9992\
        );

    \I__2200\ : InMux
    port map (
            O => \N__10013\,
            I => \N__9992\
        );

    \I__2199\ : InMux
    port map (
            O => \N__10010\,
            I => \N__9992\
        );

    \I__2198\ : InMux
    port map (
            O => \N__10009\,
            I => \N__9992\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__9992\,
            I => \N__9989\
        );

    \I__2196\ : Span4Mux_v
    port map (
            O => \N__9989\,
            I => \N__9986\
        );

    \I__2195\ : Span4Mux_h
    port map (
            O => \N__9986\,
            I => \N__9983\
        );

    \I__2194\ : Odrv4
    port map (
            O => \N__9983\,
            I => waddr_c_11
        );

    \I__2193\ : CascadeMux
    port map (
            O => \N__9980\,
            I => \N__9973\
        );

    \I__2192\ : CascadeMux
    port map (
            O => \N__9979\,
            I => \N__9969\
        );

    \I__2191\ : CascadeMux
    port map (
            O => \N__9978\,
            I => \N__9965\
        );

    \I__2190\ : CascadeMux
    port map (
            O => \N__9977\,
            I => \N__9961\
        );

    \I__2189\ : InMux
    port map (
            O => \N__9976\,
            I => \N__9944\
        );

    \I__2188\ : InMux
    port map (
            O => \N__9973\,
            I => \N__9944\
        );

    \I__2187\ : InMux
    port map (
            O => \N__9972\,
            I => \N__9944\
        );

    \I__2186\ : InMux
    port map (
            O => \N__9969\,
            I => \N__9944\
        );

    \I__2185\ : InMux
    port map (
            O => \N__9968\,
            I => \N__9944\
        );

    \I__2184\ : InMux
    port map (
            O => \N__9965\,
            I => \N__9944\
        );

    \I__2183\ : InMux
    port map (
            O => \N__9964\,
            I => \N__9944\
        );

    \I__2182\ : InMux
    port map (
            O => \N__9961\,
            I => \N__9944\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__9944\,
            I => \N__9941\
        );

    \I__2180\ : Odrv12
    port map (
            O => \N__9941\,
            I => waddr_c_12
        );

    \I__2179\ : CEMux
    port map (
            O => \N__9938\,
            I => \N__9932\
        );

    \I__2178\ : CEMux
    port map (
            O => \N__9937\,
            I => \N__9929\
        );

    \I__2177\ : CEMux
    port map (
            O => \N__9936\,
            I => \N__9926\
        );

    \I__2176\ : CEMux
    port map (
            O => \N__9935\,
            I => \N__9923\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__9932\,
            I => \N__9918\
        );

    \I__2174\ : LocalMux
    port map (
            O => \N__9929\,
            I => \N__9918\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__9926\,
            I => \N__9913\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__9923\,
            I => \N__9913\
        );

    \I__2171\ : Span4Mux_v
    port map (
            O => \N__9918\,
            I => \N__9908\
        );

    \I__2170\ : Span4Mux_v
    port map (
            O => \N__9913\,
            I => \N__9908\
        );

    \I__2169\ : Sp12to4
    port map (
            O => \N__9908\,
            I => \N__9905\
        );

    \I__2168\ : Span12Mux_h
    port map (
            O => \N__9905\,
            I => \N__9902\
        );

    \I__2167\ : Span12Mux_v
    port map (
            O => \N__9902\,
            I => \N__9899\
        );

    \I__2166\ : Odrv12
    port map (
            O => \N__9899\,
            I => \mem_WE_28\
        );

    \I__2165\ : InMux
    port map (
            O => \N__9896\,
            I => \N__9893\
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__9893\,
            I => \N__9890\
        );

    \I__2163\ : Span4Mux_s1_v
    port map (
            O => \N__9890\,
            I => \N__9887\
        );

    \I__2162\ : Sp12to4
    port map (
            O => \N__9887\,
            I => \N__9884\
        );

    \I__2161\ : Span12Mux_h
    port map (
            O => \N__9884\,
            I => \N__9881\
        );

    \I__2160\ : Odrv12
    port map (
            O => \N__9881\,
            I => mem_out_bus0_0
        );

    \I__2159\ : InMux
    port map (
            O => \N__9878\,
            I => \N__9875\
        );

    \I__2158\ : LocalMux
    port map (
            O => \N__9875\,
            I => \N__9872\
        );

    \I__2157\ : Span4Mux_s1_v
    port map (
            O => \N__9872\,
            I => \N__9869\
        );

    \I__2156\ : Odrv4
    port map (
            O => \N__9869\,
            I => mem_out_bus4_0
        );

    \I__2155\ : InMux
    port map (
            O => \N__9866\,
            I => \N__9863\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__9863\,
            I => \N__9860\
        );

    \I__2153\ : Span12Mux_h
    port map (
            O => \N__9860\,
            I => \N__9857\
        );

    \I__2152\ : Span12Mux_h
    port map (
            O => \N__9857\,
            I => \N__9854\
        );

    \I__2151\ : Odrv12
    port map (
            O => \N__9854\,
            I => mem_out_bus0_1
        );

    \I__2150\ : InMux
    port map (
            O => \N__9851\,
            I => \N__9848\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__9848\,
            I => \N__9845\
        );

    \I__2148\ : Odrv4
    port map (
            O => \N__9845\,
            I => mem_out_bus4_1
        );

    \I__2147\ : InMux
    port map (
            O => \N__9842\,
            I => \N__9839\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__9839\,
            I => \N__9836\
        );

    \I__2145\ : Odrv12
    port map (
            O => \N__9836\,
            I => mem_out_bus4_7
        );

    \I__2144\ : InMux
    port map (
            O => \N__9833\,
            I => \N__9830\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__9830\,
            I => \N__9827\
        );

    \I__2142\ : Span12Mux_h
    port map (
            O => \N__9827\,
            I => \N__9824\
        );

    \I__2141\ : Odrv12
    port map (
            O => \N__9824\,
            I => mem_out_bus0_7
        );

    \I__2140\ : CascadeMux
    port map (
            O => \N__9821\,
            I => \N__9818\
        );

    \I__2139\ : CascadeBuf
    port map (
            O => \N__9818\,
            I => \N__9815\
        );

    \I__2138\ : CascadeMux
    port map (
            O => \N__9815\,
            I => \N__9811\
        );

    \I__2137\ : CascadeMux
    port map (
            O => \N__9814\,
            I => \N__9808\
        );

    \I__2136\ : CascadeBuf
    port map (
            O => \N__9811\,
            I => \N__9805\
        );

    \I__2135\ : CascadeBuf
    port map (
            O => \N__9808\,
            I => \N__9802\
        );

    \I__2134\ : CascadeMux
    port map (
            O => \N__9805\,
            I => \N__9799\
        );

    \I__2133\ : CascadeMux
    port map (
            O => \N__9802\,
            I => \N__9796\
        );

    \I__2132\ : CascadeBuf
    port map (
            O => \N__9799\,
            I => \N__9793\
        );

    \I__2131\ : CascadeBuf
    port map (
            O => \N__9796\,
            I => \N__9790\
        );

    \I__2130\ : CascadeMux
    port map (
            O => \N__9793\,
            I => \N__9787\
        );

    \I__2129\ : CascadeMux
    port map (
            O => \N__9790\,
            I => \N__9784\
        );

    \I__2128\ : CascadeBuf
    port map (
            O => \N__9787\,
            I => \N__9781\
        );

    \I__2127\ : CascadeBuf
    port map (
            O => \N__9784\,
            I => \N__9778\
        );

    \I__2126\ : CascadeMux
    port map (
            O => \N__9781\,
            I => \N__9775\
        );

    \I__2125\ : CascadeMux
    port map (
            O => \N__9778\,
            I => \N__9772\
        );

    \I__2124\ : CascadeBuf
    port map (
            O => \N__9775\,
            I => \N__9769\
        );

    \I__2123\ : CascadeBuf
    port map (
            O => \N__9772\,
            I => \N__9766\
        );

    \I__2122\ : CascadeMux
    port map (
            O => \N__9769\,
            I => \N__9763\
        );

    \I__2121\ : CascadeMux
    port map (
            O => \N__9766\,
            I => \N__9760\
        );

    \I__2120\ : CascadeBuf
    port map (
            O => \N__9763\,
            I => \N__9757\
        );

    \I__2119\ : CascadeBuf
    port map (
            O => \N__9760\,
            I => \N__9754\
        );

    \I__2118\ : CascadeMux
    port map (
            O => \N__9757\,
            I => \N__9751\
        );

    \I__2117\ : CascadeMux
    port map (
            O => \N__9754\,
            I => \N__9748\
        );

    \I__2116\ : CascadeBuf
    port map (
            O => \N__9751\,
            I => \N__9745\
        );

    \I__2115\ : CascadeBuf
    port map (
            O => \N__9748\,
            I => \N__9742\
        );

    \I__2114\ : CascadeMux
    port map (
            O => \N__9745\,
            I => \N__9739\
        );

    \I__2113\ : CascadeMux
    port map (
            O => \N__9742\,
            I => \N__9736\
        );

    \I__2112\ : CascadeBuf
    port map (
            O => \N__9739\,
            I => \N__9733\
        );

    \I__2111\ : CascadeBuf
    port map (
            O => \N__9736\,
            I => \N__9730\
        );

    \I__2110\ : CascadeMux
    port map (
            O => \N__9733\,
            I => \N__9727\
        );

    \I__2109\ : CascadeMux
    port map (
            O => \N__9730\,
            I => \N__9724\
        );

    \I__2108\ : CascadeBuf
    port map (
            O => \N__9727\,
            I => \N__9721\
        );

    \I__2107\ : CascadeBuf
    port map (
            O => \N__9724\,
            I => \N__9718\
        );

    \I__2106\ : CascadeMux
    port map (
            O => \N__9721\,
            I => \N__9715\
        );

    \I__2105\ : CascadeMux
    port map (
            O => \N__9718\,
            I => \N__9712\
        );

    \I__2104\ : CascadeBuf
    port map (
            O => \N__9715\,
            I => \N__9709\
        );

    \I__2103\ : CascadeBuf
    port map (
            O => \N__9712\,
            I => \N__9706\
        );

    \I__2102\ : CascadeMux
    port map (
            O => \N__9709\,
            I => \N__9703\
        );

    \I__2101\ : CascadeMux
    port map (
            O => \N__9706\,
            I => \N__9700\
        );

    \I__2100\ : CascadeBuf
    port map (
            O => \N__9703\,
            I => \N__9697\
        );

    \I__2099\ : CascadeBuf
    port map (
            O => \N__9700\,
            I => \N__9694\
        );

    \I__2098\ : CascadeMux
    port map (
            O => \N__9697\,
            I => \N__9691\
        );

    \I__2097\ : CascadeMux
    port map (
            O => \N__9694\,
            I => \N__9688\
        );

    \I__2096\ : CascadeBuf
    port map (
            O => \N__9691\,
            I => \N__9685\
        );

    \I__2095\ : CascadeBuf
    port map (
            O => \N__9688\,
            I => \N__9682\
        );

    \I__2094\ : CascadeMux
    port map (
            O => \N__9685\,
            I => \N__9679\
        );

    \I__2093\ : CascadeMux
    port map (
            O => \N__9682\,
            I => \N__9676\
        );

    \I__2092\ : CascadeBuf
    port map (
            O => \N__9679\,
            I => \N__9673\
        );

    \I__2091\ : CascadeBuf
    port map (
            O => \N__9676\,
            I => \N__9670\
        );

    \I__2090\ : CascadeMux
    port map (
            O => \N__9673\,
            I => \N__9667\
        );

    \I__2089\ : CascadeMux
    port map (
            O => \N__9670\,
            I => \N__9664\
        );

    \I__2088\ : CascadeBuf
    port map (
            O => \N__9667\,
            I => \N__9661\
        );

    \I__2087\ : CascadeBuf
    port map (
            O => \N__9664\,
            I => \N__9658\
        );

    \I__2086\ : CascadeMux
    port map (
            O => \N__9661\,
            I => \N__9655\
        );

    \I__2085\ : CascadeMux
    port map (
            O => \N__9658\,
            I => \N__9652\
        );

    \I__2084\ : CascadeBuf
    port map (
            O => \N__9655\,
            I => \N__9649\
        );

    \I__2083\ : CascadeBuf
    port map (
            O => \N__9652\,
            I => \N__9646\
        );

    \I__2082\ : CascadeMux
    port map (
            O => \N__9649\,
            I => \N__9643\
        );

    \I__2081\ : CascadeMux
    port map (
            O => \N__9646\,
            I => \N__9640\
        );

    \I__2080\ : InMux
    port map (
            O => \N__9643\,
            I => \N__9637\
        );

    \I__2079\ : CascadeBuf
    port map (
            O => \N__9640\,
            I => \N__9634\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__9637\,
            I => \N__9631\
        );

    \I__2077\ : CascadeMux
    port map (
            O => \N__9634\,
            I => \N__9628\
        );

    \I__2076\ : Span4Mux_s2_v
    port map (
            O => \N__9631\,
            I => \N__9625\
        );

    \I__2075\ : InMux
    port map (
            O => \N__9628\,
            I => \N__9622\
        );

    \I__2074\ : Span4Mux_h
    port map (
            O => \N__9625\,
            I => \N__9619\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__9622\,
            I => \N__9616\
        );

    \I__2072\ : Sp12to4
    port map (
            O => \N__9619\,
            I => \N__9613\
        );

    \I__2071\ : Span4Mux_s2_v
    port map (
            O => \N__9616\,
            I => \N__9610\
        );

    \I__2070\ : Span12Mux_h
    port map (
            O => \N__9613\,
            I => \N__9605\
        );

    \I__2069\ : Sp12to4
    port map (
            O => \N__9610\,
            I => \N__9605\
        );

    \I__2068\ : Odrv12
    port map (
            O => \N__9605\,
            I => waddr_c_0
        );

    \I__2067\ : CEMux
    port map (
            O => \N__9602\,
            I => \N__9599\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__9599\,
            I => \N__9594\
        );

    \I__2065\ : CEMux
    port map (
            O => \N__9598\,
            I => \N__9591\
        );

    \I__2064\ : CEMux
    port map (
            O => \N__9597\,
            I => \N__9588\
        );

    \I__2063\ : Span4Mux_v
    port map (
            O => \N__9594\,
            I => \N__9580\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__9591\,
            I => \N__9580\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__9588\,
            I => \N__9580\
        );

    \I__2060\ : CEMux
    port map (
            O => \N__9587\,
            I => \N__9577\
        );

    \I__2059\ : Span4Mux_v
    port map (
            O => \N__9580\,
            I => \N__9572\
        );

    \I__2058\ : LocalMux
    port map (
            O => \N__9577\,
            I => \N__9572\
        );

    \I__2057\ : Span4Mux_h
    port map (
            O => \N__9572\,
            I => \N__9569\
        );

    \I__2056\ : Odrv4
    port map (
            O => \N__9569\,
            I => \mem_WE_4\
        );

    \I__2055\ : CEMux
    port map (
            O => \N__9566\,
            I => \N__9562\
        );

    \I__2054\ : CEMux
    port map (
            O => \N__9565\,
            I => \N__9559\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__9562\,
            I => \N__9555\
        );

    \I__2052\ : LocalMux
    port map (
            O => \N__9559\,
            I => \N__9552\
        );

    \I__2051\ : CEMux
    port map (
            O => \N__9558\,
            I => \N__9549\
        );

    \I__2050\ : Span4Mux_s2_v
    port map (
            O => \N__9555\,
            I => \N__9542\
        );

    \I__2049\ : Span4Mux_h
    port map (
            O => \N__9552\,
            I => \N__9542\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__9549\,
            I => \N__9542\
        );

    \I__2047\ : Span4Mux_v
    port map (
            O => \N__9542\,
            I => \N__9538\
        );

    \I__2046\ : CEMux
    port map (
            O => \N__9541\,
            I => \N__9535\
        );

    \I__2045\ : Sp12to4
    port map (
            O => \N__9538\,
            I => \N__9530\
        );

    \I__2044\ : LocalMux
    port map (
            O => \N__9535\,
            I => \N__9530\
        );

    \I__2043\ : Span12Mux_h
    port map (
            O => \N__9530\,
            I => \N__9527\
        );

    \I__2042\ : Odrv12
    port map (
            O => \N__9527\,
            I => \mem_WE_0\
        );

    \I__2041\ : InMux
    port map (
            O => \N__9524\,
            I => \N__9517\
        );

    \I__2040\ : InMux
    port map (
            O => \N__9523\,
            I => \N__9513\
        );

    \I__2039\ : InMux
    port map (
            O => \N__9522\,
            I => \N__9510\
        );

    \I__2038\ : InMux
    port map (
            O => \N__9521\,
            I => \N__9507\
        );

    \I__2037\ : InMux
    port map (
            O => \N__9520\,
            I => \N__9504\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__9517\,
            I => \N__9501\
        );

    \I__2035\ : InMux
    port map (
            O => \N__9516\,
            I => \N__9498\
        );

    \I__2034\ : LocalMux
    port map (
            O => \N__9513\,
            I => \N__9494\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__9510\,
            I => \N__9491\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__9507\,
            I => \N__9488\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__9504\,
            I => \N__9484\
        );

    \I__2030\ : Sp12to4
    port map (
            O => \N__9501\,
            I => \N__9479\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__9498\,
            I => \N__9479\
        );

    \I__2028\ : InMux
    port map (
            O => \N__9497\,
            I => \N__9476\
        );

    \I__2027\ : Span4Mux_h
    port map (
            O => \N__9494\,
            I => \N__9473\
        );

    \I__2026\ : Span12Mux_h
    port map (
            O => \N__9491\,
            I => \N__9468\
        );

    \I__2025\ : Span12Mux_h
    port map (
            O => \N__9488\,
            I => \N__9468\
        );

    \I__2024\ : InMux
    port map (
            O => \N__9487\,
            I => \N__9465\
        );

    \I__2023\ : Span12Mux_h
    port map (
            O => \N__9484\,
            I => \N__9462\
        );

    \I__2022\ : Span12Mux_v
    port map (
            O => \N__9479\,
            I => \N__9459\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__9476\,
            I => \N__9456\
        );

    \I__2020\ : Span4Mux_h
    port map (
            O => \N__9473\,
            I => \N__9453\
        );

    \I__2019\ : Span12Mux_v
    port map (
            O => \N__9468\,
            I => \N__9450\
        );

    \I__2018\ : LocalMux
    port map (
            O => \N__9465\,
            I => \N__9447\
        );

    \I__2017\ : Span12Mux_v
    port map (
            O => \N__9462\,
            I => \N__9442\
        );

    \I__2016\ : Span12Mux_h
    port map (
            O => \N__9459\,
            I => \N__9442\
        );

    \I__2015\ : Span12Mux_h
    port map (
            O => \N__9456\,
            I => \N__9439\
        );

    \I__2014\ : Span4Mux_h
    port map (
            O => \N__9453\,
            I => \N__9436\
        );

    \I__2013\ : Span12Mux_v
    port map (
            O => \N__9450\,
            I => \N__9431\
        );

    \I__2012\ : Span12Mux_h
    port map (
            O => \N__9447\,
            I => \N__9431\
        );

    \I__2011\ : Odrv12
    port map (
            O => \N__9442\,
            I => din_c_5
        );

    \I__2010\ : Odrv12
    port map (
            O => \N__9439\,
            I => din_c_5
        );

    \I__2009\ : Odrv4
    port map (
            O => \N__9436\,
            I => din_c_5
        );

    \I__2008\ : Odrv12
    port map (
            O => \N__9431\,
            I => din_c_5
        );

    \I__2007\ : CascadeMux
    port map (
            O => \N__9422\,
            I => \N__9419\
        );

    \I__2006\ : CascadeBuf
    port map (
            O => \N__9419\,
            I => \N__9416\
        );

    \I__2005\ : CascadeMux
    port map (
            O => \N__9416\,
            I => \N__9413\
        );

    \I__2004\ : CascadeBuf
    port map (
            O => \N__9413\,
            I => \N__9409\
        );

    \I__2003\ : CascadeMux
    port map (
            O => \N__9412\,
            I => \N__9406\
        );

    \I__2002\ : CascadeMux
    port map (
            O => \N__9409\,
            I => \N__9403\
        );

    \I__2001\ : CascadeBuf
    port map (
            O => \N__9406\,
            I => \N__9400\
        );

    \I__2000\ : CascadeBuf
    port map (
            O => \N__9403\,
            I => \N__9397\
        );

    \I__1999\ : CascadeMux
    port map (
            O => \N__9400\,
            I => \N__9394\
        );

    \I__1998\ : CascadeMux
    port map (
            O => \N__9397\,
            I => \N__9391\
        );

    \I__1997\ : CascadeBuf
    port map (
            O => \N__9394\,
            I => \N__9388\
        );

    \I__1996\ : CascadeBuf
    port map (
            O => \N__9391\,
            I => \N__9385\
        );

    \I__1995\ : CascadeMux
    port map (
            O => \N__9388\,
            I => \N__9382\
        );

    \I__1994\ : CascadeMux
    port map (
            O => \N__9385\,
            I => \N__9379\
        );

    \I__1993\ : CascadeBuf
    port map (
            O => \N__9382\,
            I => \N__9376\
        );

    \I__1992\ : CascadeBuf
    port map (
            O => \N__9379\,
            I => \N__9373\
        );

    \I__1991\ : CascadeMux
    port map (
            O => \N__9376\,
            I => \N__9370\
        );

    \I__1990\ : CascadeMux
    port map (
            O => \N__9373\,
            I => \N__9367\
        );

    \I__1989\ : CascadeBuf
    port map (
            O => \N__9370\,
            I => \N__9364\
        );

    \I__1988\ : CascadeBuf
    port map (
            O => \N__9367\,
            I => \N__9361\
        );

    \I__1987\ : CascadeMux
    port map (
            O => \N__9364\,
            I => \N__9358\
        );

    \I__1986\ : CascadeMux
    port map (
            O => \N__9361\,
            I => \N__9355\
        );

    \I__1985\ : CascadeBuf
    port map (
            O => \N__9358\,
            I => \N__9352\
        );

    \I__1984\ : CascadeBuf
    port map (
            O => \N__9355\,
            I => \N__9349\
        );

    \I__1983\ : CascadeMux
    port map (
            O => \N__9352\,
            I => \N__9346\
        );

    \I__1982\ : CascadeMux
    port map (
            O => \N__9349\,
            I => \N__9343\
        );

    \I__1981\ : CascadeBuf
    port map (
            O => \N__9346\,
            I => \N__9340\
        );

    \I__1980\ : CascadeBuf
    port map (
            O => \N__9343\,
            I => \N__9337\
        );

    \I__1979\ : CascadeMux
    port map (
            O => \N__9340\,
            I => \N__9334\
        );

    \I__1978\ : CascadeMux
    port map (
            O => \N__9337\,
            I => \N__9331\
        );

    \I__1977\ : CascadeBuf
    port map (
            O => \N__9334\,
            I => \N__9328\
        );

    \I__1976\ : CascadeBuf
    port map (
            O => \N__9331\,
            I => \N__9325\
        );

    \I__1975\ : CascadeMux
    port map (
            O => \N__9328\,
            I => \N__9322\
        );

    \I__1974\ : CascadeMux
    port map (
            O => \N__9325\,
            I => \N__9319\
        );

    \I__1973\ : CascadeBuf
    port map (
            O => \N__9322\,
            I => \N__9316\
        );

    \I__1972\ : CascadeBuf
    port map (
            O => \N__9319\,
            I => \N__9313\
        );

    \I__1971\ : CascadeMux
    port map (
            O => \N__9316\,
            I => \N__9310\
        );

    \I__1970\ : CascadeMux
    port map (
            O => \N__9313\,
            I => \N__9307\
        );

    \I__1969\ : CascadeBuf
    port map (
            O => \N__9310\,
            I => \N__9304\
        );

    \I__1968\ : CascadeBuf
    port map (
            O => \N__9307\,
            I => \N__9301\
        );

    \I__1967\ : CascadeMux
    port map (
            O => \N__9304\,
            I => \N__9298\
        );

    \I__1966\ : CascadeMux
    port map (
            O => \N__9301\,
            I => \N__9295\
        );

    \I__1965\ : CascadeBuf
    port map (
            O => \N__9298\,
            I => \N__9292\
        );

    \I__1964\ : CascadeBuf
    port map (
            O => \N__9295\,
            I => \N__9289\
        );

    \I__1963\ : CascadeMux
    port map (
            O => \N__9292\,
            I => \N__9286\
        );

    \I__1962\ : CascadeMux
    port map (
            O => \N__9289\,
            I => \N__9283\
        );

    \I__1961\ : CascadeBuf
    port map (
            O => \N__9286\,
            I => \N__9280\
        );

    \I__1960\ : CascadeBuf
    port map (
            O => \N__9283\,
            I => \N__9277\
        );

    \I__1959\ : CascadeMux
    port map (
            O => \N__9280\,
            I => \N__9274\
        );

    \I__1958\ : CascadeMux
    port map (
            O => \N__9277\,
            I => \N__9271\
        );

    \I__1957\ : CascadeBuf
    port map (
            O => \N__9274\,
            I => \N__9268\
        );

    \I__1956\ : CascadeBuf
    port map (
            O => \N__9271\,
            I => \N__9265\
        );

    \I__1955\ : CascadeMux
    port map (
            O => \N__9268\,
            I => \N__9262\
        );

    \I__1954\ : CascadeMux
    port map (
            O => \N__9265\,
            I => \N__9259\
        );

    \I__1953\ : CascadeBuf
    port map (
            O => \N__9262\,
            I => \N__9256\
        );

    \I__1952\ : CascadeBuf
    port map (
            O => \N__9259\,
            I => \N__9253\
        );

    \I__1951\ : CascadeMux
    port map (
            O => \N__9256\,
            I => \N__9250\
        );

    \I__1950\ : CascadeMux
    port map (
            O => \N__9253\,
            I => \N__9247\
        );

    \I__1949\ : CascadeBuf
    port map (
            O => \N__9250\,
            I => \N__9244\
        );

    \I__1948\ : InMux
    port map (
            O => \N__9247\,
            I => \N__9241\
        );

    \I__1947\ : CascadeMux
    port map (
            O => \N__9244\,
            I => \N__9238\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__9241\,
            I => \N__9235\
        );

    \I__1945\ : CascadeBuf
    port map (
            O => \N__9238\,
            I => \N__9232\
        );

    \I__1944\ : Span4Mux_s3_v
    port map (
            O => \N__9235\,
            I => \N__9229\
        );

    \I__1943\ : CascadeMux
    port map (
            O => \N__9232\,
            I => \N__9226\
        );

    \I__1942\ : Span4Mux_v
    port map (
            O => \N__9229\,
            I => \N__9223\
        );

    \I__1941\ : InMux
    port map (
            O => \N__9226\,
            I => \N__9220\
        );

    \I__1940\ : Sp12to4
    port map (
            O => \N__9223\,
            I => \N__9217\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__9220\,
            I => \N__9214\
        );

    \I__1938\ : Span12Mux_h
    port map (
            O => \N__9217\,
            I => \N__9211\
        );

    \I__1937\ : Span12Mux_s7_v
    port map (
            O => \N__9214\,
            I => \N__9208\
        );

    \I__1936\ : Odrv12
    port map (
            O => \N__9211\,
            I => raddr_c_5
        );

    \I__1935\ : Odrv12
    port map (
            O => \N__9208\,
            I => raddr_c_5
        );

    \I__1934\ : CascadeMux
    port map (
            O => \N__9203\,
            I => \N__9200\
        );

    \I__1933\ : CascadeBuf
    port map (
            O => \N__9200\,
            I => \N__9197\
        );

    \I__1932\ : CascadeMux
    port map (
            O => \N__9197\,
            I => \N__9194\
        );

    \I__1931\ : CascadeBuf
    port map (
            O => \N__9194\,
            I => \N__9190\
        );

    \I__1930\ : CascadeMux
    port map (
            O => \N__9193\,
            I => \N__9187\
        );

    \I__1929\ : CascadeMux
    port map (
            O => \N__9190\,
            I => \N__9184\
        );

    \I__1928\ : CascadeBuf
    port map (
            O => \N__9187\,
            I => \N__9181\
        );

    \I__1927\ : CascadeBuf
    port map (
            O => \N__9184\,
            I => \N__9178\
        );

    \I__1926\ : CascadeMux
    port map (
            O => \N__9181\,
            I => \N__9175\
        );

    \I__1925\ : CascadeMux
    port map (
            O => \N__9178\,
            I => \N__9172\
        );

    \I__1924\ : CascadeBuf
    port map (
            O => \N__9175\,
            I => \N__9169\
        );

    \I__1923\ : CascadeBuf
    port map (
            O => \N__9172\,
            I => \N__9166\
        );

    \I__1922\ : CascadeMux
    port map (
            O => \N__9169\,
            I => \N__9163\
        );

    \I__1921\ : CascadeMux
    port map (
            O => \N__9166\,
            I => \N__9160\
        );

    \I__1920\ : CascadeBuf
    port map (
            O => \N__9163\,
            I => \N__9157\
        );

    \I__1919\ : CascadeBuf
    port map (
            O => \N__9160\,
            I => \N__9154\
        );

    \I__1918\ : CascadeMux
    port map (
            O => \N__9157\,
            I => \N__9151\
        );

    \I__1917\ : CascadeMux
    port map (
            O => \N__9154\,
            I => \N__9148\
        );

    \I__1916\ : CascadeBuf
    port map (
            O => \N__9151\,
            I => \N__9145\
        );

    \I__1915\ : CascadeBuf
    port map (
            O => \N__9148\,
            I => \N__9142\
        );

    \I__1914\ : CascadeMux
    port map (
            O => \N__9145\,
            I => \N__9139\
        );

    \I__1913\ : CascadeMux
    port map (
            O => \N__9142\,
            I => \N__9136\
        );

    \I__1912\ : CascadeBuf
    port map (
            O => \N__9139\,
            I => \N__9133\
        );

    \I__1911\ : CascadeBuf
    port map (
            O => \N__9136\,
            I => \N__9130\
        );

    \I__1910\ : CascadeMux
    port map (
            O => \N__9133\,
            I => \N__9127\
        );

    \I__1909\ : CascadeMux
    port map (
            O => \N__9130\,
            I => \N__9124\
        );

    \I__1908\ : CascadeBuf
    port map (
            O => \N__9127\,
            I => \N__9121\
        );

    \I__1907\ : CascadeBuf
    port map (
            O => \N__9124\,
            I => \N__9118\
        );

    \I__1906\ : CascadeMux
    port map (
            O => \N__9121\,
            I => \N__9115\
        );

    \I__1905\ : CascadeMux
    port map (
            O => \N__9118\,
            I => \N__9112\
        );

    \I__1904\ : CascadeBuf
    port map (
            O => \N__9115\,
            I => \N__9109\
        );

    \I__1903\ : CascadeBuf
    port map (
            O => \N__9112\,
            I => \N__9106\
        );

    \I__1902\ : CascadeMux
    port map (
            O => \N__9109\,
            I => \N__9103\
        );

    \I__1901\ : CascadeMux
    port map (
            O => \N__9106\,
            I => \N__9100\
        );

    \I__1900\ : CascadeBuf
    port map (
            O => \N__9103\,
            I => \N__9097\
        );

    \I__1899\ : CascadeBuf
    port map (
            O => \N__9100\,
            I => \N__9094\
        );

    \I__1898\ : CascadeMux
    port map (
            O => \N__9097\,
            I => \N__9091\
        );

    \I__1897\ : CascadeMux
    port map (
            O => \N__9094\,
            I => \N__9088\
        );

    \I__1896\ : CascadeBuf
    port map (
            O => \N__9091\,
            I => \N__9085\
        );

    \I__1895\ : CascadeBuf
    port map (
            O => \N__9088\,
            I => \N__9082\
        );

    \I__1894\ : CascadeMux
    port map (
            O => \N__9085\,
            I => \N__9079\
        );

    \I__1893\ : CascadeMux
    port map (
            O => \N__9082\,
            I => \N__9076\
        );

    \I__1892\ : CascadeBuf
    port map (
            O => \N__9079\,
            I => \N__9073\
        );

    \I__1891\ : CascadeBuf
    port map (
            O => \N__9076\,
            I => \N__9070\
        );

    \I__1890\ : CascadeMux
    port map (
            O => \N__9073\,
            I => \N__9067\
        );

    \I__1889\ : CascadeMux
    port map (
            O => \N__9070\,
            I => \N__9064\
        );

    \I__1888\ : CascadeBuf
    port map (
            O => \N__9067\,
            I => \N__9061\
        );

    \I__1887\ : CascadeBuf
    port map (
            O => \N__9064\,
            I => \N__9058\
        );

    \I__1886\ : CascadeMux
    port map (
            O => \N__9061\,
            I => \N__9055\
        );

    \I__1885\ : CascadeMux
    port map (
            O => \N__9058\,
            I => \N__9052\
        );

    \I__1884\ : CascadeBuf
    port map (
            O => \N__9055\,
            I => \N__9049\
        );

    \I__1883\ : CascadeBuf
    port map (
            O => \N__9052\,
            I => \N__9046\
        );

    \I__1882\ : CascadeMux
    port map (
            O => \N__9049\,
            I => \N__9043\
        );

    \I__1881\ : CascadeMux
    port map (
            O => \N__9046\,
            I => \N__9040\
        );

    \I__1880\ : CascadeBuf
    port map (
            O => \N__9043\,
            I => \N__9037\
        );

    \I__1879\ : CascadeBuf
    port map (
            O => \N__9040\,
            I => \N__9034\
        );

    \I__1878\ : CascadeMux
    port map (
            O => \N__9037\,
            I => \N__9031\
        );

    \I__1877\ : CascadeMux
    port map (
            O => \N__9034\,
            I => \N__9028\
        );

    \I__1876\ : CascadeBuf
    port map (
            O => \N__9031\,
            I => \N__9025\
        );

    \I__1875\ : InMux
    port map (
            O => \N__9028\,
            I => \N__9022\
        );

    \I__1874\ : CascadeMux
    port map (
            O => \N__9025\,
            I => \N__9019\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__9022\,
            I => \N__9016\
        );

    \I__1872\ : CascadeBuf
    port map (
            O => \N__9019\,
            I => \N__9013\
        );

    \I__1871\ : Span4Mux_s3_v
    port map (
            O => \N__9016\,
            I => \N__9010\
        );

    \I__1870\ : CascadeMux
    port map (
            O => \N__9013\,
            I => \N__9007\
        );

    \I__1869\ : Sp12to4
    port map (
            O => \N__9010\,
            I => \N__9004\
        );

    \I__1868\ : InMux
    port map (
            O => \N__9007\,
            I => \N__9001\
        );

    \I__1867\ : Span12Mux_h
    port map (
            O => \N__9004\,
            I => \N__8998\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__9001\,
            I => \N__8995\
        );

    \I__1865\ : Span12Mux_h
    port map (
            O => \N__8998\,
            I => \N__8992\
        );

    \I__1864\ : IoSpan4Mux
    port map (
            O => \N__8995\,
            I => \N__8989\
        );

    \I__1863\ : Odrv12
    port map (
            O => \N__8992\,
            I => waddr_c_3
        );

    \I__1862\ : Odrv4
    port map (
            O => \N__8989\,
            I => waddr_c_3
        );

    \I__1861\ : CascadeMux
    port map (
            O => \N__8984\,
            I => \N__8981\
        );

    \I__1860\ : CascadeBuf
    port map (
            O => \N__8981\,
            I => \N__8978\
        );

    \I__1859\ : CascadeMux
    port map (
            O => \N__8978\,
            I => \N__8975\
        );

    \I__1858\ : CascadeBuf
    port map (
            O => \N__8975\,
            I => \N__8972\
        );

    \I__1857\ : CascadeMux
    port map (
            O => \N__8972\,
            I => \N__8969\
        );

    \I__1856\ : CascadeBuf
    port map (
            O => \N__8969\,
            I => \N__8965\
        );

    \I__1855\ : CascadeMux
    port map (
            O => \N__8968\,
            I => \N__8962\
        );

    \I__1854\ : CascadeMux
    port map (
            O => \N__8965\,
            I => \N__8959\
        );

    \I__1853\ : CascadeBuf
    port map (
            O => \N__8962\,
            I => \N__8956\
        );

    \I__1852\ : CascadeBuf
    port map (
            O => \N__8959\,
            I => \N__8953\
        );

    \I__1851\ : CascadeMux
    port map (
            O => \N__8956\,
            I => \N__8950\
        );

    \I__1850\ : CascadeMux
    port map (
            O => \N__8953\,
            I => \N__8947\
        );

    \I__1849\ : CascadeBuf
    port map (
            O => \N__8950\,
            I => \N__8944\
        );

    \I__1848\ : CascadeBuf
    port map (
            O => \N__8947\,
            I => \N__8941\
        );

    \I__1847\ : CascadeMux
    port map (
            O => \N__8944\,
            I => \N__8938\
        );

    \I__1846\ : CascadeMux
    port map (
            O => \N__8941\,
            I => \N__8935\
        );

    \I__1845\ : CascadeBuf
    port map (
            O => \N__8938\,
            I => \N__8932\
        );

    \I__1844\ : CascadeBuf
    port map (
            O => \N__8935\,
            I => \N__8929\
        );

    \I__1843\ : CascadeMux
    port map (
            O => \N__8932\,
            I => \N__8926\
        );

    \I__1842\ : CascadeMux
    port map (
            O => \N__8929\,
            I => \N__8923\
        );

    \I__1841\ : CascadeBuf
    port map (
            O => \N__8926\,
            I => \N__8920\
        );

    \I__1840\ : CascadeBuf
    port map (
            O => \N__8923\,
            I => \N__8917\
        );

    \I__1839\ : CascadeMux
    port map (
            O => \N__8920\,
            I => \N__8914\
        );

    \I__1838\ : CascadeMux
    port map (
            O => \N__8917\,
            I => \N__8911\
        );

    \I__1837\ : CascadeBuf
    port map (
            O => \N__8914\,
            I => \N__8908\
        );

    \I__1836\ : CascadeBuf
    port map (
            O => \N__8911\,
            I => \N__8905\
        );

    \I__1835\ : CascadeMux
    port map (
            O => \N__8908\,
            I => \N__8902\
        );

    \I__1834\ : CascadeMux
    port map (
            O => \N__8905\,
            I => \N__8899\
        );

    \I__1833\ : CascadeBuf
    port map (
            O => \N__8902\,
            I => \N__8896\
        );

    \I__1832\ : CascadeBuf
    port map (
            O => \N__8899\,
            I => \N__8893\
        );

    \I__1831\ : CascadeMux
    port map (
            O => \N__8896\,
            I => \N__8890\
        );

    \I__1830\ : CascadeMux
    port map (
            O => \N__8893\,
            I => \N__8887\
        );

    \I__1829\ : CascadeBuf
    port map (
            O => \N__8890\,
            I => \N__8884\
        );

    \I__1828\ : CascadeBuf
    port map (
            O => \N__8887\,
            I => \N__8881\
        );

    \I__1827\ : CascadeMux
    port map (
            O => \N__8884\,
            I => \N__8878\
        );

    \I__1826\ : CascadeMux
    port map (
            O => \N__8881\,
            I => \N__8875\
        );

    \I__1825\ : CascadeBuf
    port map (
            O => \N__8878\,
            I => \N__8872\
        );

    \I__1824\ : CascadeBuf
    port map (
            O => \N__8875\,
            I => \N__8869\
        );

    \I__1823\ : CascadeMux
    port map (
            O => \N__8872\,
            I => \N__8866\
        );

    \I__1822\ : CascadeMux
    port map (
            O => \N__8869\,
            I => \N__8863\
        );

    \I__1821\ : CascadeBuf
    port map (
            O => \N__8866\,
            I => \N__8860\
        );

    \I__1820\ : CascadeBuf
    port map (
            O => \N__8863\,
            I => \N__8857\
        );

    \I__1819\ : CascadeMux
    port map (
            O => \N__8860\,
            I => \N__8854\
        );

    \I__1818\ : CascadeMux
    port map (
            O => \N__8857\,
            I => \N__8851\
        );

    \I__1817\ : CascadeBuf
    port map (
            O => \N__8854\,
            I => \N__8848\
        );

    \I__1816\ : CascadeBuf
    port map (
            O => \N__8851\,
            I => \N__8845\
        );

    \I__1815\ : CascadeMux
    port map (
            O => \N__8848\,
            I => \N__8842\
        );

    \I__1814\ : CascadeMux
    port map (
            O => \N__8845\,
            I => \N__8839\
        );

    \I__1813\ : CascadeBuf
    port map (
            O => \N__8842\,
            I => \N__8836\
        );

    \I__1812\ : CascadeBuf
    port map (
            O => \N__8839\,
            I => \N__8833\
        );

    \I__1811\ : CascadeMux
    port map (
            O => \N__8836\,
            I => \N__8830\
        );

    \I__1810\ : CascadeMux
    port map (
            O => \N__8833\,
            I => \N__8827\
        );

    \I__1809\ : CascadeBuf
    port map (
            O => \N__8830\,
            I => \N__8824\
        );

    \I__1808\ : CascadeBuf
    port map (
            O => \N__8827\,
            I => \N__8821\
        );

    \I__1807\ : CascadeMux
    port map (
            O => \N__8824\,
            I => \N__8818\
        );

    \I__1806\ : CascadeMux
    port map (
            O => \N__8821\,
            I => \N__8815\
        );

    \I__1805\ : CascadeBuf
    port map (
            O => \N__8818\,
            I => \N__8812\
        );

    \I__1804\ : InMux
    port map (
            O => \N__8815\,
            I => \N__8809\
        );

    \I__1803\ : CascadeMux
    port map (
            O => \N__8812\,
            I => \N__8806\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__8809\,
            I => \N__8803\
        );

    \I__1801\ : CascadeBuf
    port map (
            O => \N__8806\,
            I => \N__8800\
        );

    \I__1800\ : Span4Mux_s3_v
    port map (
            O => \N__8803\,
            I => \N__8797\
        );

    \I__1799\ : CascadeMux
    port map (
            O => \N__8800\,
            I => \N__8794\
        );

    \I__1798\ : Span4Mux_h
    port map (
            O => \N__8797\,
            I => \N__8791\
        );

    \I__1797\ : CascadeBuf
    port map (
            O => \N__8794\,
            I => \N__8788\
        );

    \I__1796\ : Sp12to4
    port map (
            O => \N__8791\,
            I => \N__8785\
        );

    \I__1795\ : CascadeMux
    port map (
            O => \N__8788\,
            I => \N__8782\
        );

    \I__1794\ : Span12Mux_h
    port map (
            O => \N__8785\,
            I => \N__8779\
        );

    \I__1793\ : InMux
    port map (
            O => \N__8782\,
            I => \N__8776\
        );

    \I__1792\ : Odrv12
    port map (
            O => \N__8779\,
            I => waddr_c_6
        );

    \I__1791\ : LocalMux
    port map (
            O => \N__8776\,
            I => waddr_c_6
        );

    \I__1790\ : ClkMux
    port map (
            O => \N__8771\,
            I => \N__8675\
        );

    \I__1789\ : ClkMux
    port map (
            O => \N__8770\,
            I => \N__8675\
        );

    \I__1788\ : ClkMux
    port map (
            O => \N__8769\,
            I => \N__8675\
        );

    \I__1787\ : ClkMux
    port map (
            O => \N__8768\,
            I => \N__8675\
        );

    \I__1786\ : ClkMux
    port map (
            O => \N__8767\,
            I => \N__8675\
        );

    \I__1785\ : ClkMux
    port map (
            O => \N__8766\,
            I => \N__8675\
        );

    \I__1784\ : ClkMux
    port map (
            O => \N__8765\,
            I => \N__8675\
        );

    \I__1783\ : ClkMux
    port map (
            O => \N__8764\,
            I => \N__8675\
        );

    \I__1782\ : ClkMux
    port map (
            O => \N__8763\,
            I => \N__8675\
        );

    \I__1781\ : ClkMux
    port map (
            O => \N__8762\,
            I => \N__8675\
        );

    \I__1780\ : ClkMux
    port map (
            O => \N__8761\,
            I => \N__8675\
        );

    \I__1779\ : ClkMux
    port map (
            O => \N__8760\,
            I => \N__8675\
        );

    \I__1778\ : ClkMux
    port map (
            O => \N__8759\,
            I => \N__8675\
        );

    \I__1777\ : ClkMux
    port map (
            O => \N__8758\,
            I => \N__8675\
        );

    \I__1776\ : ClkMux
    port map (
            O => \N__8757\,
            I => \N__8675\
        );

    \I__1775\ : ClkMux
    port map (
            O => \N__8756\,
            I => \N__8675\
        );

    \I__1774\ : ClkMux
    port map (
            O => \N__8755\,
            I => \N__8675\
        );

    \I__1773\ : ClkMux
    port map (
            O => \N__8754\,
            I => \N__8675\
        );

    \I__1772\ : ClkMux
    port map (
            O => \N__8753\,
            I => \N__8675\
        );

    \I__1771\ : ClkMux
    port map (
            O => \N__8752\,
            I => \N__8675\
        );

    \I__1770\ : ClkMux
    port map (
            O => \N__8751\,
            I => \N__8675\
        );

    \I__1769\ : ClkMux
    port map (
            O => \N__8750\,
            I => \N__8675\
        );

    \I__1768\ : ClkMux
    port map (
            O => \N__8749\,
            I => \N__8675\
        );

    \I__1767\ : ClkMux
    port map (
            O => \N__8748\,
            I => \N__8675\
        );

    \I__1766\ : ClkMux
    port map (
            O => \N__8747\,
            I => \N__8675\
        );

    \I__1765\ : ClkMux
    port map (
            O => \N__8746\,
            I => \N__8675\
        );

    \I__1764\ : ClkMux
    port map (
            O => \N__8745\,
            I => \N__8675\
        );

    \I__1763\ : ClkMux
    port map (
            O => \N__8744\,
            I => \N__8675\
        );

    \I__1762\ : ClkMux
    port map (
            O => \N__8743\,
            I => \N__8675\
        );

    \I__1761\ : ClkMux
    port map (
            O => \N__8742\,
            I => \N__8675\
        );

    \I__1760\ : ClkMux
    port map (
            O => \N__8741\,
            I => \N__8675\
        );

    \I__1759\ : ClkMux
    port map (
            O => \N__8740\,
            I => \N__8675\
        );

    \I__1758\ : GlobalMux
    port map (
            O => \N__8675\,
            I => \N__8672\
        );

    \I__1757\ : gio2CtrlBuf
    port map (
            O => \N__8672\,
            I => wclk_c_g
        );

    \I__1756\ : CascadeMux
    port map (
            O => \N__8669\,
            I => \N__8666\
        );

    \I__1755\ : CascadeBuf
    port map (
            O => \N__8666\,
            I => \N__8663\
        );

    \I__1754\ : CascadeMux
    port map (
            O => \N__8663\,
            I => \N__8659\
        );

    \I__1753\ : CascadeMux
    port map (
            O => \N__8662\,
            I => \N__8656\
        );

    \I__1752\ : CascadeBuf
    port map (
            O => \N__8659\,
            I => \N__8653\
        );

    \I__1751\ : CascadeBuf
    port map (
            O => \N__8656\,
            I => \N__8650\
        );

    \I__1750\ : CascadeMux
    port map (
            O => \N__8653\,
            I => \N__8647\
        );

    \I__1749\ : CascadeMux
    port map (
            O => \N__8650\,
            I => \N__8644\
        );

    \I__1748\ : CascadeBuf
    port map (
            O => \N__8647\,
            I => \N__8641\
        );

    \I__1747\ : CascadeBuf
    port map (
            O => \N__8644\,
            I => \N__8638\
        );

    \I__1746\ : CascadeMux
    port map (
            O => \N__8641\,
            I => \N__8635\
        );

    \I__1745\ : CascadeMux
    port map (
            O => \N__8638\,
            I => \N__8632\
        );

    \I__1744\ : CascadeBuf
    port map (
            O => \N__8635\,
            I => \N__8629\
        );

    \I__1743\ : CascadeBuf
    port map (
            O => \N__8632\,
            I => \N__8626\
        );

    \I__1742\ : CascadeMux
    port map (
            O => \N__8629\,
            I => \N__8623\
        );

    \I__1741\ : CascadeMux
    port map (
            O => \N__8626\,
            I => \N__8620\
        );

    \I__1740\ : CascadeBuf
    port map (
            O => \N__8623\,
            I => \N__8617\
        );

    \I__1739\ : CascadeBuf
    port map (
            O => \N__8620\,
            I => \N__8614\
        );

    \I__1738\ : CascadeMux
    port map (
            O => \N__8617\,
            I => \N__8611\
        );

    \I__1737\ : CascadeMux
    port map (
            O => \N__8614\,
            I => \N__8608\
        );

    \I__1736\ : CascadeBuf
    port map (
            O => \N__8611\,
            I => \N__8605\
        );

    \I__1735\ : CascadeBuf
    port map (
            O => \N__8608\,
            I => \N__8602\
        );

    \I__1734\ : CascadeMux
    port map (
            O => \N__8605\,
            I => \N__8599\
        );

    \I__1733\ : CascadeMux
    port map (
            O => \N__8602\,
            I => \N__8596\
        );

    \I__1732\ : CascadeBuf
    port map (
            O => \N__8599\,
            I => \N__8593\
        );

    \I__1731\ : CascadeBuf
    port map (
            O => \N__8596\,
            I => \N__8590\
        );

    \I__1730\ : CascadeMux
    port map (
            O => \N__8593\,
            I => \N__8587\
        );

    \I__1729\ : CascadeMux
    port map (
            O => \N__8590\,
            I => \N__8584\
        );

    \I__1728\ : CascadeBuf
    port map (
            O => \N__8587\,
            I => \N__8581\
        );

    \I__1727\ : CascadeBuf
    port map (
            O => \N__8584\,
            I => \N__8578\
        );

    \I__1726\ : CascadeMux
    port map (
            O => \N__8581\,
            I => \N__8575\
        );

    \I__1725\ : CascadeMux
    port map (
            O => \N__8578\,
            I => \N__8572\
        );

    \I__1724\ : CascadeBuf
    port map (
            O => \N__8575\,
            I => \N__8569\
        );

    \I__1723\ : CascadeBuf
    port map (
            O => \N__8572\,
            I => \N__8566\
        );

    \I__1722\ : CascadeMux
    port map (
            O => \N__8569\,
            I => \N__8563\
        );

    \I__1721\ : CascadeMux
    port map (
            O => \N__8566\,
            I => \N__8560\
        );

    \I__1720\ : CascadeBuf
    port map (
            O => \N__8563\,
            I => \N__8557\
        );

    \I__1719\ : CascadeBuf
    port map (
            O => \N__8560\,
            I => \N__8554\
        );

    \I__1718\ : CascadeMux
    port map (
            O => \N__8557\,
            I => \N__8551\
        );

    \I__1717\ : CascadeMux
    port map (
            O => \N__8554\,
            I => \N__8548\
        );

    \I__1716\ : CascadeBuf
    port map (
            O => \N__8551\,
            I => \N__8545\
        );

    \I__1715\ : CascadeBuf
    port map (
            O => \N__8548\,
            I => \N__8542\
        );

    \I__1714\ : CascadeMux
    port map (
            O => \N__8545\,
            I => \N__8539\
        );

    \I__1713\ : CascadeMux
    port map (
            O => \N__8542\,
            I => \N__8536\
        );

    \I__1712\ : CascadeBuf
    port map (
            O => \N__8539\,
            I => \N__8533\
        );

    \I__1711\ : CascadeBuf
    port map (
            O => \N__8536\,
            I => \N__8530\
        );

    \I__1710\ : CascadeMux
    port map (
            O => \N__8533\,
            I => \N__8527\
        );

    \I__1709\ : CascadeMux
    port map (
            O => \N__8530\,
            I => \N__8524\
        );

    \I__1708\ : CascadeBuf
    port map (
            O => \N__8527\,
            I => \N__8521\
        );

    \I__1707\ : CascadeBuf
    port map (
            O => \N__8524\,
            I => \N__8518\
        );

    \I__1706\ : CascadeMux
    port map (
            O => \N__8521\,
            I => \N__8515\
        );

    \I__1705\ : CascadeMux
    port map (
            O => \N__8518\,
            I => \N__8512\
        );

    \I__1704\ : CascadeBuf
    port map (
            O => \N__8515\,
            I => \N__8509\
        );

    \I__1703\ : CascadeBuf
    port map (
            O => \N__8512\,
            I => \N__8506\
        );

    \I__1702\ : CascadeMux
    port map (
            O => \N__8509\,
            I => \N__8503\
        );

    \I__1701\ : CascadeMux
    port map (
            O => \N__8506\,
            I => \N__8500\
        );

    \I__1700\ : CascadeBuf
    port map (
            O => \N__8503\,
            I => \N__8497\
        );

    \I__1699\ : CascadeBuf
    port map (
            O => \N__8500\,
            I => \N__8494\
        );

    \I__1698\ : CascadeMux
    port map (
            O => \N__8497\,
            I => \N__8491\
        );

    \I__1697\ : CascadeMux
    port map (
            O => \N__8494\,
            I => \N__8488\
        );

    \I__1696\ : InMux
    port map (
            O => \N__8491\,
            I => \N__8485\
        );

    \I__1695\ : CascadeBuf
    port map (
            O => \N__8488\,
            I => \N__8482\
        );

    \I__1694\ : LocalMux
    port map (
            O => \N__8485\,
            I => \N__8479\
        );

    \I__1693\ : CascadeMux
    port map (
            O => \N__8482\,
            I => \N__8476\
        );

    \I__1692\ : Span4Mux_h
    port map (
            O => \N__8479\,
            I => \N__8473\
        );

    \I__1691\ : InMux
    port map (
            O => \N__8476\,
            I => \N__8470\
        );

    \I__1690\ : Span4Mux_h
    port map (
            O => \N__8473\,
            I => \N__8467\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__8470\,
            I => \N__8464\
        );

    \I__1688\ : Sp12to4
    port map (
            O => \N__8467\,
            I => \N__8461\
        );

    \I__1687\ : Span4Mux_h
    port map (
            O => \N__8464\,
            I => \N__8458\
        );

    \I__1686\ : Span12Mux_s11_v
    port map (
            O => \N__8461\,
            I => \N__8455\
        );

    \I__1685\ : Sp12to4
    port map (
            O => \N__8458\,
            I => \N__8452\
        );

    \I__1684\ : Span12Mux_h
    port map (
            O => \N__8455\,
            I => \N__8447\
        );

    \I__1683\ : Span12Mux_s11_v
    port map (
            O => \N__8452\,
            I => \N__8447\
        );

    \I__1682\ : Odrv12
    port map (
            O => \N__8447\,
            I => raddr_c_2
        );

    \I__1681\ : CascadeMux
    port map (
            O => \N__8444\,
            I => \N__8441\
        );

    \I__1680\ : CascadeBuf
    port map (
            O => \N__8441\,
            I => \N__8438\
        );

    \I__1679\ : CascadeMux
    port map (
            O => \N__8438\,
            I => \N__8434\
        );

    \I__1678\ : CascadeMux
    port map (
            O => \N__8437\,
            I => \N__8431\
        );

    \I__1677\ : CascadeBuf
    port map (
            O => \N__8434\,
            I => \N__8428\
        );

    \I__1676\ : CascadeBuf
    port map (
            O => \N__8431\,
            I => \N__8425\
        );

    \I__1675\ : CascadeMux
    port map (
            O => \N__8428\,
            I => \N__8422\
        );

    \I__1674\ : CascadeMux
    port map (
            O => \N__8425\,
            I => \N__8419\
        );

    \I__1673\ : CascadeBuf
    port map (
            O => \N__8422\,
            I => \N__8416\
        );

    \I__1672\ : CascadeBuf
    port map (
            O => \N__8419\,
            I => \N__8413\
        );

    \I__1671\ : CascadeMux
    port map (
            O => \N__8416\,
            I => \N__8410\
        );

    \I__1670\ : CascadeMux
    port map (
            O => \N__8413\,
            I => \N__8407\
        );

    \I__1669\ : CascadeBuf
    port map (
            O => \N__8410\,
            I => \N__8404\
        );

    \I__1668\ : CascadeBuf
    port map (
            O => \N__8407\,
            I => \N__8401\
        );

    \I__1667\ : CascadeMux
    port map (
            O => \N__8404\,
            I => \N__8398\
        );

    \I__1666\ : CascadeMux
    port map (
            O => \N__8401\,
            I => \N__8395\
        );

    \I__1665\ : CascadeBuf
    port map (
            O => \N__8398\,
            I => \N__8392\
        );

    \I__1664\ : CascadeBuf
    port map (
            O => \N__8395\,
            I => \N__8389\
        );

    \I__1663\ : CascadeMux
    port map (
            O => \N__8392\,
            I => \N__8386\
        );

    \I__1662\ : CascadeMux
    port map (
            O => \N__8389\,
            I => \N__8383\
        );

    \I__1661\ : CascadeBuf
    port map (
            O => \N__8386\,
            I => \N__8380\
        );

    \I__1660\ : CascadeBuf
    port map (
            O => \N__8383\,
            I => \N__8377\
        );

    \I__1659\ : CascadeMux
    port map (
            O => \N__8380\,
            I => \N__8374\
        );

    \I__1658\ : CascadeMux
    port map (
            O => \N__8377\,
            I => \N__8371\
        );

    \I__1657\ : CascadeBuf
    port map (
            O => \N__8374\,
            I => \N__8368\
        );

    \I__1656\ : CascadeBuf
    port map (
            O => \N__8371\,
            I => \N__8365\
        );

    \I__1655\ : CascadeMux
    port map (
            O => \N__8368\,
            I => \N__8362\
        );

    \I__1654\ : CascadeMux
    port map (
            O => \N__8365\,
            I => \N__8359\
        );

    \I__1653\ : CascadeBuf
    port map (
            O => \N__8362\,
            I => \N__8356\
        );

    \I__1652\ : CascadeBuf
    port map (
            O => \N__8359\,
            I => \N__8353\
        );

    \I__1651\ : CascadeMux
    port map (
            O => \N__8356\,
            I => \N__8350\
        );

    \I__1650\ : CascadeMux
    port map (
            O => \N__8353\,
            I => \N__8347\
        );

    \I__1649\ : CascadeBuf
    port map (
            O => \N__8350\,
            I => \N__8344\
        );

    \I__1648\ : CascadeBuf
    port map (
            O => \N__8347\,
            I => \N__8341\
        );

    \I__1647\ : CascadeMux
    port map (
            O => \N__8344\,
            I => \N__8338\
        );

    \I__1646\ : CascadeMux
    port map (
            O => \N__8341\,
            I => \N__8335\
        );

    \I__1645\ : CascadeBuf
    port map (
            O => \N__8338\,
            I => \N__8332\
        );

    \I__1644\ : CascadeBuf
    port map (
            O => \N__8335\,
            I => \N__8329\
        );

    \I__1643\ : CascadeMux
    port map (
            O => \N__8332\,
            I => \N__8326\
        );

    \I__1642\ : CascadeMux
    port map (
            O => \N__8329\,
            I => \N__8323\
        );

    \I__1641\ : CascadeBuf
    port map (
            O => \N__8326\,
            I => \N__8320\
        );

    \I__1640\ : CascadeBuf
    port map (
            O => \N__8323\,
            I => \N__8317\
        );

    \I__1639\ : CascadeMux
    port map (
            O => \N__8320\,
            I => \N__8314\
        );

    \I__1638\ : CascadeMux
    port map (
            O => \N__8317\,
            I => \N__8311\
        );

    \I__1637\ : CascadeBuf
    port map (
            O => \N__8314\,
            I => \N__8308\
        );

    \I__1636\ : CascadeBuf
    port map (
            O => \N__8311\,
            I => \N__8305\
        );

    \I__1635\ : CascadeMux
    port map (
            O => \N__8308\,
            I => \N__8302\
        );

    \I__1634\ : CascadeMux
    port map (
            O => \N__8305\,
            I => \N__8299\
        );

    \I__1633\ : CascadeBuf
    port map (
            O => \N__8302\,
            I => \N__8296\
        );

    \I__1632\ : CascadeBuf
    port map (
            O => \N__8299\,
            I => \N__8293\
        );

    \I__1631\ : CascadeMux
    port map (
            O => \N__8296\,
            I => \N__8290\
        );

    \I__1630\ : CascadeMux
    port map (
            O => \N__8293\,
            I => \N__8287\
        );

    \I__1629\ : CascadeBuf
    port map (
            O => \N__8290\,
            I => \N__8284\
        );

    \I__1628\ : CascadeBuf
    port map (
            O => \N__8287\,
            I => \N__8281\
        );

    \I__1627\ : CascadeMux
    port map (
            O => \N__8284\,
            I => \N__8278\
        );

    \I__1626\ : CascadeMux
    port map (
            O => \N__8281\,
            I => \N__8275\
        );

    \I__1625\ : CascadeBuf
    port map (
            O => \N__8278\,
            I => \N__8272\
        );

    \I__1624\ : CascadeBuf
    port map (
            O => \N__8275\,
            I => \N__8269\
        );

    \I__1623\ : CascadeMux
    port map (
            O => \N__8272\,
            I => \N__8266\
        );

    \I__1622\ : CascadeMux
    port map (
            O => \N__8269\,
            I => \N__8263\
        );

    \I__1621\ : InMux
    port map (
            O => \N__8266\,
            I => \N__8260\
        );

    \I__1620\ : CascadeBuf
    port map (
            O => \N__8263\,
            I => \N__8257\
        );

    \I__1619\ : LocalMux
    port map (
            O => \N__8260\,
            I => \N__8254\
        );

    \I__1618\ : CascadeMux
    port map (
            O => \N__8257\,
            I => \N__8251\
        );

    \I__1617\ : Span4Mux_v
    port map (
            O => \N__8254\,
            I => \N__8248\
        );

    \I__1616\ : InMux
    port map (
            O => \N__8251\,
            I => \N__8245\
        );

    \I__1615\ : Sp12to4
    port map (
            O => \N__8248\,
            I => \N__8242\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__8245\,
            I => \N__8239\
        );

    \I__1613\ : Span12Mux_h
    port map (
            O => \N__8242\,
            I => \N__8236\
        );

    \I__1612\ : Span12Mux_s5_v
    port map (
            O => \N__8239\,
            I => \N__8233\
        );

    \I__1611\ : Odrv12
    port map (
            O => \N__8236\,
            I => raddr_c_7
        );

    \I__1610\ : Odrv12
    port map (
            O => \N__8233\,
            I => raddr_c_7
        );

    \I__1609\ : CascadeMux
    port map (
            O => \N__8228\,
            I => \N__8225\
        );

    \I__1608\ : CascadeBuf
    port map (
            O => \N__8225\,
            I => \N__8222\
        );

    \I__1607\ : CascadeMux
    port map (
            O => \N__8222\,
            I => \N__8219\
        );

    \I__1606\ : CascadeBuf
    port map (
            O => \N__8219\,
            I => \N__8216\
        );

    \I__1605\ : CascadeMux
    port map (
            O => \N__8216\,
            I => \N__8213\
        );

    \I__1604\ : CascadeBuf
    port map (
            O => \N__8213\,
            I => \N__8209\
        );

    \I__1603\ : CascadeMux
    port map (
            O => \N__8212\,
            I => \N__8206\
        );

    \I__1602\ : CascadeMux
    port map (
            O => \N__8209\,
            I => \N__8203\
        );

    \I__1601\ : CascadeBuf
    port map (
            O => \N__8206\,
            I => \N__8200\
        );

    \I__1600\ : CascadeBuf
    port map (
            O => \N__8203\,
            I => \N__8197\
        );

    \I__1599\ : CascadeMux
    port map (
            O => \N__8200\,
            I => \N__8194\
        );

    \I__1598\ : CascadeMux
    port map (
            O => \N__8197\,
            I => \N__8191\
        );

    \I__1597\ : CascadeBuf
    port map (
            O => \N__8194\,
            I => \N__8188\
        );

    \I__1596\ : CascadeBuf
    port map (
            O => \N__8191\,
            I => \N__8185\
        );

    \I__1595\ : CascadeMux
    port map (
            O => \N__8188\,
            I => \N__8182\
        );

    \I__1594\ : CascadeMux
    port map (
            O => \N__8185\,
            I => \N__8179\
        );

    \I__1593\ : CascadeBuf
    port map (
            O => \N__8182\,
            I => \N__8176\
        );

    \I__1592\ : CascadeBuf
    port map (
            O => \N__8179\,
            I => \N__8173\
        );

    \I__1591\ : CascadeMux
    port map (
            O => \N__8176\,
            I => \N__8170\
        );

    \I__1590\ : CascadeMux
    port map (
            O => \N__8173\,
            I => \N__8167\
        );

    \I__1589\ : CascadeBuf
    port map (
            O => \N__8170\,
            I => \N__8164\
        );

    \I__1588\ : CascadeBuf
    port map (
            O => \N__8167\,
            I => \N__8161\
        );

    \I__1587\ : CascadeMux
    port map (
            O => \N__8164\,
            I => \N__8158\
        );

    \I__1586\ : CascadeMux
    port map (
            O => \N__8161\,
            I => \N__8155\
        );

    \I__1585\ : CascadeBuf
    port map (
            O => \N__8158\,
            I => \N__8152\
        );

    \I__1584\ : CascadeBuf
    port map (
            O => \N__8155\,
            I => \N__8149\
        );

    \I__1583\ : CascadeMux
    port map (
            O => \N__8152\,
            I => \N__8146\
        );

    \I__1582\ : CascadeMux
    port map (
            O => \N__8149\,
            I => \N__8143\
        );

    \I__1581\ : CascadeBuf
    port map (
            O => \N__8146\,
            I => \N__8140\
        );

    \I__1580\ : CascadeBuf
    port map (
            O => \N__8143\,
            I => \N__8137\
        );

    \I__1579\ : CascadeMux
    port map (
            O => \N__8140\,
            I => \N__8134\
        );

    \I__1578\ : CascadeMux
    port map (
            O => \N__8137\,
            I => \N__8131\
        );

    \I__1577\ : CascadeBuf
    port map (
            O => \N__8134\,
            I => \N__8128\
        );

    \I__1576\ : CascadeBuf
    port map (
            O => \N__8131\,
            I => \N__8125\
        );

    \I__1575\ : CascadeMux
    port map (
            O => \N__8128\,
            I => \N__8122\
        );

    \I__1574\ : CascadeMux
    port map (
            O => \N__8125\,
            I => \N__8119\
        );

    \I__1573\ : CascadeBuf
    port map (
            O => \N__8122\,
            I => \N__8116\
        );

    \I__1572\ : CascadeBuf
    port map (
            O => \N__8119\,
            I => \N__8113\
        );

    \I__1571\ : CascadeMux
    port map (
            O => \N__8116\,
            I => \N__8110\
        );

    \I__1570\ : CascadeMux
    port map (
            O => \N__8113\,
            I => \N__8107\
        );

    \I__1569\ : CascadeBuf
    port map (
            O => \N__8110\,
            I => \N__8104\
        );

    \I__1568\ : CascadeBuf
    port map (
            O => \N__8107\,
            I => \N__8101\
        );

    \I__1567\ : CascadeMux
    port map (
            O => \N__8104\,
            I => \N__8098\
        );

    \I__1566\ : CascadeMux
    port map (
            O => \N__8101\,
            I => \N__8095\
        );

    \I__1565\ : CascadeBuf
    port map (
            O => \N__8098\,
            I => \N__8092\
        );

    \I__1564\ : CascadeBuf
    port map (
            O => \N__8095\,
            I => \N__8089\
        );

    \I__1563\ : CascadeMux
    port map (
            O => \N__8092\,
            I => \N__8086\
        );

    \I__1562\ : CascadeMux
    port map (
            O => \N__8089\,
            I => \N__8083\
        );

    \I__1561\ : CascadeBuf
    port map (
            O => \N__8086\,
            I => \N__8080\
        );

    \I__1560\ : CascadeBuf
    port map (
            O => \N__8083\,
            I => \N__8077\
        );

    \I__1559\ : CascadeMux
    port map (
            O => \N__8080\,
            I => \N__8074\
        );

    \I__1558\ : CascadeMux
    port map (
            O => \N__8077\,
            I => \N__8071\
        );

    \I__1557\ : CascadeBuf
    port map (
            O => \N__8074\,
            I => \N__8068\
        );

    \I__1556\ : CascadeBuf
    port map (
            O => \N__8071\,
            I => \N__8065\
        );

    \I__1555\ : CascadeMux
    port map (
            O => \N__8068\,
            I => \N__8062\
        );

    \I__1554\ : CascadeMux
    port map (
            O => \N__8065\,
            I => \N__8059\
        );

    \I__1553\ : CascadeBuf
    port map (
            O => \N__8062\,
            I => \N__8056\
        );

    \I__1552\ : InMux
    port map (
            O => \N__8059\,
            I => \N__8053\
        );

    \I__1551\ : CascadeMux
    port map (
            O => \N__8056\,
            I => \N__8050\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__8053\,
            I => \N__8047\
        );

    \I__1549\ : CascadeBuf
    port map (
            O => \N__8050\,
            I => \N__8044\
        );

    \I__1548\ : Span4Mux_s1_v
    port map (
            O => \N__8047\,
            I => \N__8041\
        );

    \I__1547\ : CascadeMux
    port map (
            O => \N__8044\,
            I => \N__8038\
        );

    \I__1546\ : Span4Mux_h
    port map (
            O => \N__8041\,
            I => \N__8035\
        );

    \I__1545\ : CascadeBuf
    port map (
            O => \N__8038\,
            I => \N__8032\
        );

    \I__1544\ : Sp12to4
    port map (
            O => \N__8035\,
            I => \N__8029\
        );

    \I__1543\ : CascadeMux
    port map (
            O => \N__8032\,
            I => \N__8026\
        );

    \I__1542\ : Span12Mux_h
    port map (
            O => \N__8029\,
            I => \N__8023\
        );

    \I__1541\ : InMux
    port map (
            O => \N__8026\,
            I => \N__8020\
        );

    \I__1540\ : Odrv12
    port map (
            O => \N__8023\,
            I => waddr_c_5
        );

    \I__1539\ : LocalMux
    port map (
            O => \N__8020\,
            I => waddr_c_5
        );

    \I__1538\ : InMux
    port map (
            O => \N__8015\,
            I => \N__8009\
        );

    \I__1537\ : InMux
    port map (
            O => \N__8014\,
            I => \N__8006\
        );

    \I__1536\ : InMux
    port map (
            O => \N__8013\,
            I => \N__7999\
        );

    \I__1535\ : InMux
    port map (
            O => \N__8012\,
            I => \N__7996\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__8009\,
            I => \N__7993\
        );

    \I__1533\ : LocalMux
    port map (
            O => \N__8006\,
            I => \N__7990\
        );

    \I__1532\ : InMux
    port map (
            O => \N__8005\,
            I => \N__7987\
        );

    \I__1531\ : InMux
    port map (
            O => \N__8004\,
            I => \N__7984\
        );

    \I__1530\ : InMux
    port map (
            O => \N__8003\,
            I => \N__7981\
        );

    \I__1529\ : InMux
    port map (
            O => \N__8002\,
            I => \N__7978\
        );

    \I__1528\ : LocalMux
    port map (
            O => \N__7999\,
            I => \N__7975\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__7996\,
            I => \N__7972\
        );

    \I__1526\ : Span12Mux_h
    port map (
            O => \N__7993\,
            I => \N__7967\
        );

    \I__1525\ : Span12Mux_h
    port map (
            O => \N__7990\,
            I => \N__7967\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__7987\,
            I => \N__7964\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__7984\,
            I => \N__7961\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__7981\,
            I => \N__7958\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__7978\,
            I => \N__7955\
        );

    \I__1520\ : Span4Mux_v
    port map (
            O => \N__7975\,
            I => \N__7952\
        );

    \I__1519\ : Span4Mux_v
    port map (
            O => \N__7972\,
            I => \N__7949\
        );

    \I__1518\ : Span12Mux_v
    port map (
            O => \N__7967\,
            I => \N__7946\
        );

    \I__1517\ : Span12Mux_h
    port map (
            O => \N__7964\,
            I => \N__7941\
        );

    \I__1516\ : Span12Mux_h
    port map (
            O => \N__7961\,
            I => \N__7941\
        );

    \I__1515\ : Span12Mux_h
    port map (
            O => \N__7958\,
            I => \N__7936\
        );

    \I__1514\ : Span12Mux_h
    port map (
            O => \N__7955\,
            I => \N__7936\
        );

    \I__1513\ : Sp12to4
    port map (
            O => \N__7952\,
            I => \N__7933\
        );

    \I__1512\ : Sp12to4
    port map (
            O => \N__7949\,
            I => \N__7930\
        );

    \I__1511\ : Span12Mux_v
    port map (
            O => \N__7946\,
            I => \N__7927\
        );

    \I__1510\ : Span12Mux_v
    port map (
            O => \N__7941\,
            I => \N__7924\
        );

    \I__1509\ : Span12Mux_v
    port map (
            O => \N__7936\,
            I => \N__7917\
        );

    \I__1508\ : Span12Mux_h
    port map (
            O => \N__7933\,
            I => \N__7917\
        );

    \I__1507\ : Span12Mux_h
    port map (
            O => \N__7930\,
            I => \N__7917\
        );

    \I__1506\ : Odrv12
    port map (
            O => \N__7927\,
            I => din_c_1
        );

    \I__1505\ : Odrv12
    port map (
            O => \N__7924\,
            I => din_c_1
        );

    \I__1504\ : Odrv12
    port map (
            O => \N__7917\,
            I => din_c_1
        );

    \I__1503\ : CascadeMux
    port map (
            O => \N__7910\,
            I => \N__7907\
        );

    \I__1502\ : CascadeBuf
    port map (
            O => \N__7907\,
            I => \N__7904\
        );

    \I__1501\ : CascadeMux
    port map (
            O => \N__7904\,
            I => \N__7900\
        );

    \I__1500\ : CascadeMux
    port map (
            O => \N__7903\,
            I => \N__7897\
        );

    \I__1499\ : CascadeBuf
    port map (
            O => \N__7900\,
            I => \N__7894\
        );

    \I__1498\ : CascadeBuf
    port map (
            O => \N__7897\,
            I => \N__7891\
        );

    \I__1497\ : CascadeMux
    port map (
            O => \N__7894\,
            I => \N__7888\
        );

    \I__1496\ : CascadeMux
    port map (
            O => \N__7891\,
            I => \N__7885\
        );

    \I__1495\ : CascadeBuf
    port map (
            O => \N__7888\,
            I => \N__7882\
        );

    \I__1494\ : CascadeBuf
    port map (
            O => \N__7885\,
            I => \N__7879\
        );

    \I__1493\ : CascadeMux
    port map (
            O => \N__7882\,
            I => \N__7876\
        );

    \I__1492\ : CascadeMux
    port map (
            O => \N__7879\,
            I => \N__7873\
        );

    \I__1491\ : CascadeBuf
    port map (
            O => \N__7876\,
            I => \N__7870\
        );

    \I__1490\ : CascadeBuf
    port map (
            O => \N__7873\,
            I => \N__7867\
        );

    \I__1489\ : CascadeMux
    port map (
            O => \N__7870\,
            I => \N__7864\
        );

    \I__1488\ : CascadeMux
    port map (
            O => \N__7867\,
            I => \N__7861\
        );

    \I__1487\ : CascadeBuf
    port map (
            O => \N__7864\,
            I => \N__7858\
        );

    \I__1486\ : CascadeBuf
    port map (
            O => \N__7861\,
            I => \N__7855\
        );

    \I__1485\ : CascadeMux
    port map (
            O => \N__7858\,
            I => \N__7852\
        );

    \I__1484\ : CascadeMux
    port map (
            O => \N__7855\,
            I => \N__7849\
        );

    \I__1483\ : CascadeBuf
    port map (
            O => \N__7852\,
            I => \N__7846\
        );

    \I__1482\ : CascadeBuf
    port map (
            O => \N__7849\,
            I => \N__7843\
        );

    \I__1481\ : CascadeMux
    port map (
            O => \N__7846\,
            I => \N__7840\
        );

    \I__1480\ : CascadeMux
    port map (
            O => \N__7843\,
            I => \N__7837\
        );

    \I__1479\ : CascadeBuf
    port map (
            O => \N__7840\,
            I => \N__7834\
        );

    \I__1478\ : CascadeBuf
    port map (
            O => \N__7837\,
            I => \N__7831\
        );

    \I__1477\ : CascadeMux
    port map (
            O => \N__7834\,
            I => \N__7828\
        );

    \I__1476\ : CascadeMux
    port map (
            O => \N__7831\,
            I => \N__7825\
        );

    \I__1475\ : CascadeBuf
    port map (
            O => \N__7828\,
            I => \N__7822\
        );

    \I__1474\ : CascadeBuf
    port map (
            O => \N__7825\,
            I => \N__7819\
        );

    \I__1473\ : CascadeMux
    port map (
            O => \N__7822\,
            I => \N__7816\
        );

    \I__1472\ : CascadeMux
    port map (
            O => \N__7819\,
            I => \N__7813\
        );

    \I__1471\ : CascadeBuf
    port map (
            O => \N__7816\,
            I => \N__7810\
        );

    \I__1470\ : CascadeBuf
    port map (
            O => \N__7813\,
            I => \N__7807\
        );

    \I__1469\ : CascadeMux
    port map (
            O => \N__7810\,
            I => \N__7804\
        );

    \I__1468\ : CascadeMux
    port map (
            O => \N__7807\,
            I => \N__7801\
        );

    \I__1467\ : CascadeBuf
    port map (
            O => \N__7804\,
            I => \N__7798\
        );

    \I__1466\ : CascadeBuf
    port map (
            O => \N__7801\,
            I => \N__7795\
        );

    \I__1465\ : CascadeMux
    port map (
            O => \N__7798\,
            I => \N__7792\
        );

    \I__1464\ : CascadeMux
    port map (
            O => \N__7795\,
            I => \N__7789\
        );

    \I__1463\ : CascadeBuf
    port map (
            O => \N__7792\,
            I => \N__7786\
        );

    \I__1462\ : CascadeBuf
    port map (
            O => \N__7789\,
            I => \N__7783\
        );

    \I__1461\ : CascadeMux
    port map (
            O => \N__7786\,
            I => \N__7780\
        );

    \I__1460\ : CascadeMux
    port map (
            O => \N__7783\,
            I => \N__7777\
        );

    \I__1459\ : CascadeBuf
    port map (
            O => \N__7780\,
            I => \N__7774\
        );

    \I__1458\ : CascadeBuf
    port map (
            O => \N__7777\,
            I => \N__7771\
        );

    \I__1457\ : CascadeMux
    port map (
            O => \N__7774\,
            I => \N__7768\
        );

    \I__1456\ : CascadeMux
    port map (
            O => \N__7771\,
            I => \N__7765\
        );

    \I__1455\ : CascadeBuf
    port map (
            O => \N__7768\,
            I => \N__7762\
        );

    \I__1454\ : CascadeBuf
    port map (
            O => \N__7765\,
            I => \N__7759\
        );

    \I__1453\ : CascadeMux
    port map (
            O => \N__7762\,
            I => \N__7756\
        );

    \I__1452\ : CascadeMux
    port map (
            O => \N__7759\,
            I => \N__7753\
        );

    \I__1451\ : CascadeBuf
    port map (
            O => \N__7756\,
            I => \N__7750\
        );

    \I__1450\ : CascadeBuf
    port map (
            O => \N__7753\,
            I => \N__7747\
        );

    \I__1449\ : CascadeMux
    port map (
            O => \N__7750\,
            I => \N__7744\
        );

    \I__1448\ : CascadeMux
    port map (
            O => \N__7747\,
            I => \N__7741\
        );

    \I__1447\ : CascadeBuf
    port map (
            O => \N__7744\,
            I => \N__7738\
        );

    \I__1446\ : CascadeBuf
    port map (
            O => \N__7741\,
            I => \N__7735\
        );

    \I__1445\ : CascadeMux
    port map (
            O => \N__7738\,
            I => \N__7732\
        );

    \I__1444\ : CascadeMux
    port map (
            O => \N__7735\,
            I => \N__7729\
        );

    \I__1443\ : InMux
    port map (
            O => \N__7732\,
            I => \N__7726\
        );

    \I__1442\ : CascadeBuf
    port map (
            O => \N__7729\,
            I => \N__7723\
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__7726\,
            I => \N__7720\
        );

    \I__1440\ : CascadeMux
    port map (
            O => \N__7723\,
            I => \N__7717\
        );

    \I__1439\ : Span4Mux_v
    port map (
            O => \N__7720\,
            I => \N__7714\
        );

    \I__1438\ : InMux
    port map (
            O => \N__7717\,
            I => \N__7711\
        );

    \I__1437\ : Span4Mux_h
    port map (
            O => \N__7714\,
            I => \N__7708\
        );

    \I__1436\ : LocalMux
    port map (
            O => \N__7711\,
            I => \N__7705\
        );

    \I__1435\ : Sp12to4
    port map (
            O => \N__7708\,
            I => \N__7702\
        );

    \I__1434\ : Span4Mux_v
    port map (
            O => \N__7705\,
            I => \N__7699\
        );

    \I__1433\ : Span12Mux_h
    port map (
            O => \N__7702\,
            I => \N__7694\
        );

    \I__1432\ : Sp12to4
    port map (
            O => \N__7699\,
            I => \N__7694\
        );

    \I__1431\ : Odrv12
    port map (
            O => \N__7694\,
            I => raddr_c_8
        );

    \I__1430\ : CascadeMux
    port map (
            O => \N__7691\,
            I => \N__7688\
        );

    \I__1429\ : CascadeBuf
    port map (
            O => \N__7688\,
            I => \N__7685\
        );

    \I__1428\ : CascadeMux
    port map (
            O => \N__7685\,
            I => \N__7682\
        );

    \I__1427\ : CascadeBuf
    port map (
            O => \N__7682\,
            I => \N__7678\
        );

    \I__1426\ : CascadeMux
    port map (
            O => \N__7681\,
            I => \N__7675\
        );

    \I__1425\ : CascadeMux
    port map (
            O => \N__7678\,
            I => \N__7672\
        );

    \I__1424\ : CascadeBuf
    port map (
            O => \N__7675\,
            I => \N__7669\
        );

    \I__1423\ : CascadeBuf
    port map (
            O => \N__7672\,
            I => \N__7666\
        );

    \I__1422\ : CascadeMux
    port map (
            O => \N__7669\,
            I => \N__7663\
        );

    \I__1421\ : CascadeMux
    port map (
            O => \N__7666\,
            I => \N__7660\
        );

    \I__1420\ : CascadeBuf
    port map (
            O => \N__7663\,
            I => \N__7657\
        );

    \I__1419\ : CascadeBuf
    port map (
            O => \N__7660\,
            I => \N__7654\
        );

    \I__1418\ : CascadeMux
    port map (
            O => \N__7657\,
            I => \N__7651\
        );

    \I__1417\ : CascadeMux
    port map (
            O => \N__7654\,
            I => \N__7648\
        );

    \I__1416\ : CascadeBuf
    port map (
            O => \N__7651\,
            I => \N__7645\
        );

    \I__1415\ : CascadeBuf
    port map (
            O => \N__7648\,
            I => \N__7642\
        );

    \I__1414\ : CascadeMux
    port map (
            O => \N__7645\,
            I => \N__7639\
        );

    \I__1413\ : CascadeMux
    port map (
            O => \N__7642\,
            I => \N__7636\
        );

    \I__1412\ : CascadeBuf
    port map (
            O => \N__7639\,
            I => \N__7633\
        );

    \I__1411\ : CascadeBuf
    port map (
            O => \N__7636\,
            I => \N__7630\
        );

    \I__1410\ : CascadeMux
    port map (
            O => \N__7633\,
            I => \N__7627\
        );

    \I__1409\ : CascadeMux
    port map (
            O => \N__7630\,
            I => \N__7624\
        );

    \I__1408\ : CascadeBuf
    port map (
            O => \N__7627\,
            I => \N__7621\
        );

    \I__1407\ : CascadeBuf
    port map (
            O => \N__7624\,
            I => \N__7618\
        );

    \I__1406\ : CascadeMux
    port map (
            O => \N__7621\,
            I => \N__7615\
        );

    \I__1405\ : CascadeMux
    port map (
            O => \N__7618\,
            I => \N__7612\
        );

    \I__1404\ : CascadeBuf
    port map (
            O => \N__7615\,
            I => \N__7609\
        );

    \I__1403\ : CascadeBuf
    port map (
            O => \N__7612\,
            I => \N__7606\
        );

    \I__1402\ : CascadeMux
    port map (
            O => \N__7609\,
            I => \N__7603\
        );

    \I__1401\ : CascadeMux
    port map (
            O => \N__7606\,
            I => \N__7600\
        );

    \I__1400\ : CascadeBuf
    port map (
            O => \N__7603\,
            I => \N__7597\
        );

    \I__1399\ : CascadeBuf
    port map (
            O => \N__7600\,
            I => \N__7594\
        );

    \I__1398\ : CascadeMux
    port map (
            O => \N__7597\,
            I => \N__7591\
        );

    \I__1397\ : CascadeMux
    port map (
            O => \N__7594\,
            I => \N__7588\
        );

    \I__1396\ : CascadeBuf
    port map (
            O => \N__7591\,
            I => \N__7585\
        );

    \I__1395\ : CascadeBuf
    port map (
            O => \N__7588\,
            I => \N__7582\
        );

    \I__1394\ : CascadeMux
    port map (
            O => \N__7585\,
            I => \N__7579\
        );

    \I__1393\ : CascadeMux
    port map (
            O => \N__7582\,
            I => \N__7576\
        );

    \I__1392\ : CascadeBuf
    port map (
            O => \N__7579\,
            I => \N__7573\
        );

    \I__1391\ : CascadeBuf
    port map (
            O => \N__7576\,
            I => \N__7570\
        );

    \I__1390\ : CascadeMux
    port map (
            O => \N__7573\,
            I => \N__7567\
        );

    \I__1389\ : CascadeMux
    port map (
            O => \N__7570\,
            I => \N__7564\
        );

    \I__1388\ : CascadeBuf
    port map (
            O => \N__7567\,
            I => \N__7561\
        );

    \I__1387\ : CascadeBuf
    port map (
            O => \N__7564\,
            I => \N__7558\
        );

    \I__1386\ : CascadeMux
    port map (
            O => \N__7561\,
            I => \N__7555\
        );

    \I__1385\ : CascadeMux
    port map (
            O => \N__7558\,
            I => \N__7552\
        );

    \I__1384\ : CascadeBuf
    port map (
            O => \N__7555\,
            I => \N__7549\
        );

    \I__1383\ : CascadeBuf
    port map (
            O => \N__7552\,
            I => \N__7546\
        );

    \I__1382\ : CascadeMux
    port map (
            O => \N__7549\,
            I => \N__7543\
        );

    \I__1381\ : CascadeMux
    port map (
            O => \N__7546\,
            I => \N__7540\
        );

    \I__1380\ : CascadeBuf
    port map (
            O => \N__7543\,
            I => \N__7537\
        );

    \I__1379\ : CascadeBuf
    port map (
            O => \N__7540\,
            I => \N__7534\
        );

    \I__1378\ : CascadeMux
    port map (
            O => \N__7537\,
            I => \N__7531\
        );

    \I__1377\ : CascadeMux
    port map (
            O => \N__7534\,
            I => \N__7528\
        );

    \I__1376\ : CascadeBuf
    port map (
            O => \N__7531\,
            I => \N__7525\
        );

    \I__1375\ : CascadeBuf
    port map (
            O => \N__7528\,
            I => \N__7522\
        );

    \I__1374\ : CascadeMux
    port map (
            O => \N__7525\,
            I => \N__7519\
        );

    \I__1373\ : CascadeMux
    port map (
            O => \N__7522\,
            I => \N__7516\
        );

    \I__1372\ : CascadeBuf
    port map (
            O => \N__7519\,
            I => \N__7513\
        );

    \I__1371\ : InMux
    port map (
            O => \N__7516\,
            I => \N__7510\
        );

    \I__1370\ : CascadeMux
    port map (
            O => \N__7513\,
            I => \N__7507\
        );

    \I__1369\ : LocalMux
    port map (
            O => \N__7510\,
            I => \N__7504\
        );

    \I__1368\ : CascadeBuf
    port map (
            O => \N__7507\,
            I => \N__7501\
        );

    \I__1367\ : Span4Mux_s3_v
    port map (
            O => \N__7504\,
            I => \N__7498\
        );

    \I__1366\ : CascadeMux
    port map (
            O => \N__7501\,
            I => \N__7495\
        );

    \I__1365\ : Sp12to4
    port map (
            O => \N__7498\,
            I => \N__7492\
        );

    \I__1364\ : InMux
    port map (
            O => \N__7495\,
            I => \N__7489\
        );

    \I__1363\ : Span12Mux_h
    port map (
            O => \N__7492\,
            I => \N__7486\
        );

    \I__1362\ : LocalMux
    port map (
            O => \N__7489\,
            I => \N__7483\
        );

    \I__1361\ : Span12Mux_h
    port map (
            O => \N__7486\,
            I => \N__7480\
        );

    \I__1360\ : Span4Mux_h
    port map (
            O => \N__7483\,
            I => \N__7477\
        );

    \I__1359\ : Odrv12
    port map (
            O => \N__7480\,
            I => waddr_c_4
        );

    \I__1358\ : Odrv4
    port map (
            O => \N__7477\,
            I => waddr_c_4
        );

    \I__1357\ : CascadeMux
    port map (
            O => \N__7472\,
            I => \N__7469\
        );

    \I__1356\ : CascadeBuf
    port map (
            O => \N__7469\,
            I => \N__7466\
        );

    \I__1355\ : CascadeMux
    port map (
            O => \N__7466\,
            I => \N__7463\
        );

    \I__1354\ : CascadeBuf
    port map (
            O => \N__7463\,
            I => \N__7459\
        );

    \I__1353\ : CascadeMux
    port map (
            O => \N__7462\,
            I => \N__7456\
        );

    \I__1352\ : CascadeMux
    port map (
            O => \N__7459\,
            I => \N__7453\
        );

    \I__1351\ : CascadeBuf
    port map (
            O => \N__7456\,
            I => \N__7450\
        );

    \I__1350\ : CascadeBuf
    port map (
            O => \N__7453\,
            I => \N__7447\
        );

    \I__1349\ : CascadeMux
    port map (
            O => \N__7450\,
            I => \N__7444\
        );

    \I__1348\ : CascadeMux
    port map (
            O => \N__7447\,
            I => \N__7441\
        );

    \I__1347\ : CascadeBuf
    port map (
            O => \N__7444\,
            I => \N__7438\
        );

    \I__1346\ : CascadeBuf
    port map (
            O => \N__7441\,
            I => \N__7435\
        );

    \I__1345\ : CascadeMux
    port map (
            O => \N__7438\,
            I => \N__7432\
        );

    \I__1344\ : CascadeMux
    port map (
            O => \N__7435\,
            I => \N__7429\
        );

    \I__1343\ : CascadeBuf
    port map (
            O => \N__7432\,
            I => \N__7426\
        );

    \I__1342\ : CascadeBuf
    port map (
            O => \N__7429\,
            I => \N__7423\
        );

    \I__1341\ : CascadeMux
    port map (
            O => \N__7426\,
            I => \N__7420\
        );

    \I__1340\ : CascadeMux
    port map (
            O => \N__7423\,
            I => \N__7417\
        );

    \I__1339\ : CascadeBuf
    port map (
            O => \N__7420\,
            I => \N__7414\
        );

    \I__1338\ : CascadeBuf
    port map (
            O => \N__7417\,
            I => \N__7411\
        );

    \I__1337\ : CascadeMux
    port map (
            O => \N__7414\,
            I => \N__7408\
        );

    \I__1336\ : CascadeMux
    port map (
            O => \N__7411\,
            I => \N__7405\
        );

    \I__1335\ : CascadeBuf
    port map (
            O => \N__7408\,
            I => \N__7402\
        );

    \I__1334\ : CascadeBuf
    port map (
            O => \N__7405\,
            I => \N__7399\
        );

    \I__1333\ : CascadeMux
    port map (
            O => \N__7402\,
            I => \N__7396\
        );

    \I__1332\ : CascadeMux
    port map (
            O => \N__7399\,
            I => \N__7393\
        );

    \I__1331\ : CascadeBuf
    port map (
            O => \N__7396\,
            I => \N__7390\
        );

    \I__1330\ : CascadeBuf
    port map (
            O => \N__7393\,
            I => \N__7387\
        );

    \I__1329\ : CascadeMux
    port map (
            O => \N__7390\,
            I => \N__7384\
        );

    \I__1328\ : CascadeMux
    port map (
            O => \N__7387\,
            I => \N__7381\
        );

    \I__1327\ : CascadeBuf
    port map (
            O => \N__7384\,
            I => \N__7378\
        );

    \I__1326\ : CascadeBuf
    port map (
            O => \N__7381\,
            I => \N__7375\
        );

    \I__1325\ : CascadeMux
    port map (
            O => \N__7378\,
            I => \N__7372\
        );

    \I__1324\ : CascadeMux
    port map (
            O => \N__7375\,
            I => \N__7369\
        );

    \I__1323\ : CascadeBuf
    port map (
            O => \N__7372\,
            I => \N__7366\
        );

    \I__1322\ : CascadeBuf
    port map (
            O => \N__7369\,
            I => \N__7363\
        );

    \I__1321\ : CascadeMux
    port map (
            O => \N__7366\,
            I => \N__7360\
        );

    \I__1320\ : CascadeMux
    port map (
            O => \N__7363\,
            I => \N__7357\
        );

    \I__1319\ : CascadeBuf
    port map (
            O => \N__7360\,
            I => \N__7354\
        );

    \I__1318\ : CascadeBuf
    port map (
            O => \N__7357\,
            I => \N__7351\
        );

    \I__1317\ : CascadeMux
    port map (
            O => \N__7354\,
            I => \N__7348\
        );

    \I__1316\ : CascadeMux
    port map (
            O => \N__7351\,
            I => \N__7345\
        );

    \I__1315\ : CascadeBuf
    port map (
            O => \N__7348\,
            I => \N__7342\
        );

    \I__1314\ : CascadeBuf
    port map (
            O => \N__7345\,
            I => \N__7339\
        );

    \I__1313\ : CascadeMux
    port map (
            O => \N__7342\,
            I => \N__7336\
        );

    \I__1312\ : CascadeMux
    port map (
            O => \N__7339\,
            I => \N__7333\
        );

    \I__1311\ : CascadeBuf
    port map (
            O => \N__7336\,
            I => \N__7330\
        );

    \I__1310\ : CascadeBuf
    port map (
            O => \N__7333\,
            I => \N__7327\
        );

    \I__1309\ : CascadeMux
    port map (
            O => \N__7330\,
            I => \N__7324\
        );

    \I__1308\ : CascadeMux
    port map (
            O => \N__7327\,
            I => \N__7321\
        );

    \I__1307\ : CascadeBuf
    port map (
            O => \N__7324\,
            I => \N__7318\
        );

    \I__1306\ : CascadeBuf
    port map (
            O => \N__7321\,
            I => \N__7315\
        );

    \I__1305\ : CascadeMux
    port map (
            O => \N__7318\,
            I => \N__7312\
        );

    \I__1304\ : CascadeMux
    port map (
            O => \N__7315\,
            I => \N__7309\
        );

    \I__1303\ : CascadeBuf
    port map (
            O => \N__7312\,
            I => \N__7306\
        );

    \I__1302\ : CascadeBuf
    port map (
            O => \N__7309\,
            I => \N__7303\
        );

    \I__1301\ : CascadeMux
    port map (
            O => \N__7306\,
            I => \N__7300\
        );

    \I__1300\ : CascadeMux
    port map (
            O => \N__7303\,
            I => \N__7297\
        );

    \I__1299\ : CascadeBuf
    port map (
            O => \N__7300\,
            I => \N__7294\
        );

    \I__1298\ : InMux
    port map (
            O => \N__7297\,
            I => \N__7291\
        );

    \I__1297\ : CascadeMux
    port map (
            O => \N__7294\,
            I => \N__7288\
        );

    \I__1296\ : LocalMux
    port map (
            O => \N__7291\,
            I => \N__7285\
        );

    \I__1295\ : CascadeBuf
    port map (
            O => \N__7288\,
            I => \N__7282\
        );

    \I__1294\ : Span4Mux_h
    port map (
            O => \N__7285\,
            I => \N__7279\
        );

    \I__1293\ : CascadeMux
    port map (
            O => \N__7282\,
            I => \N__7276\
        );

    \I__1292\ : Sp12to4
    port map (
            O => \N__7279\,
            I => \N__7273\
        );

    \I__1291\ : InMux
    port map (
            O => \N__7276\,
            I => \N__7270\
        );

    \I__1290\ : Span12Mux_s11_v
    port map (
            O => \N__7273\,
            I => \N__7267\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__7270\,
            I => \N__7264\
        );

    \I__1288\ : Span12Mux_h
    port map (
            O => \N__7267\,
            I => \N__7261\
        );

    \I__1287\ : Span12Mux_s11_v
    port map (
            O => \N__7264\,
            I => \N__7258\
        );

    \I__1286\ : Odrv12
    port map (
            O => \N__7261\,
            I => raddr_c_10
        );

    \I__1285\ : Odrv12
    port map (
            O => \N__7258\,
            I => raddr_c_10
        );

    \I__1284\ : CascadeMux
    port map (
            O => \N__7253\,
            I => \N__7250\
        );

    \I__1283\ : CascadeBuf
    port map (
            O => \N__7250\,
            I => \N__7246\
        );

    \I__1282\ : CascadeMux
    port map (
            O => \N__7249\,
            I => \N__7243\
        );

    \I__1281\ : CascadeMux
    port map (
            O => \N__7246\,
            I => \N__7240\
        );

    \I__1280\ : CascadeBuf
    port map (
            O => \N__7243\,
            I => \N__7237\
        );

    \I__1279\ : CascadeBuf
    port map (
            O => \N__7240\,
            I => \N__7234\
        );

    \I__1278\ : CascadeMux
    port map (
            O => \N__7237\,
            I => \N__7231\
        );

    \I__1277\ : CascadeMux
    port map (
            O => \N__7234\,
            I => \N__7228\
        );

    \I__1276\ : CascadeBuf
    port map (
            O => \N__7231\,
            I => \N__7225\
        );

    \I__1275\ : CascadeBuf
    port map (
            O => \N__7228\,
            I => \N__7222\
        );

    \I__1274\ : CascadeMux
    port map (
            O => \N__7225\,
            I => \N__7219\
        );

    \I__1273\ : CascadeMux
    port map (
            O => \N__7222\,
            I => \N__7216\
        );

    \I__1272\ : CascadeBuf
    port map (
            O => \N__7219\,
            I => \N__7213\
        );

    \I__1271\ : CascadeBuf
    port map (
            O => \N__7216\,
            I => \N__7210\
        );

    \I__1270\ : CascadeMux
    port map (
            O => \N__7213\,
            I => \N__7207\
        );

    \I__1269\ : CascadeMux
    port map (
            O => \N__7210\,
            I => \N__7204\
        );

    \I__1268\ : CascadeBuf
    port map (
            O => \N__7207\,
            I => \N__7201\
        );

    \I__1267\ : CascadeBuf
    port map (
            O => \N__7204\,
            I => \N__7198\
        );

    \I__1266\ : CascadeMux
    port map (
            O => \N__7201\,
            I => \N__7195\
        );

    \I__1265\ : CascadeMux
    port map (
            O => \N__7198\,
            I => \N__7192\
        );

    \I__1264\ : CascadeBuf
    port map (
            O => \N__7195\,
            I => \N__7189\
        );

    \I__1263\ : CascadeBuf
    port map (
            O => \N__7192\,
            I => \N__7186\
        );

    \I__1262\ : CascadeMux
    port map (
            O => \N__7189\,
            I => \N__7183\
        );

    \I__1261\ : CascadeMux
    port map (
            O => \N__7186\,
            I => \N__7180\
        );

    \I__1260\ : CascadeBuf
    port map (
            O => \N__7183\,
            I => \N__7177\
        );

    \I__1259\ : CascadeBuf
    port map (
            O => \N__7180\,
            I => \N__7174\
        );

    \I__1258\ : CascadeMux
    port map (
            O => \N__7177\,
            I => \N__7171\
        );

    \I__1257\ : CascadeMux
    port map (
            O => \N__7174\,
            I => \N__7168\
        );

    \I__1256\ : CascadeBuf
    port map (
            O => \N__7171\,
            I => \N__7165\
        );

    \I__1255\ : CascadeBuf
    port map (
            O => \N__7168\,
            I => \N__7162\
        );

    \I__1254\ : CascadeMux
    port map (
            O => \N__7165\,
            I => \N__7159\
        );

    \I__1253\ : CascadeMux
    port map (
            O => \N__7162\,
            I => \N__7156\
        );

    \I__1252\ : CascadeBuf
    port map (
            O => \N__7159\,
            I => \N__7153\
        );

    \I__1251\ : CascadeBuf
    port map (
            O => \N__7156\,
            I => \N__7150\
        );

    \I__1250\ : CascadeMux
    port map (
            O => \N__7153\,
            I => \N__7147\
        );

    \I__1249\ : CascadeMux
    port map (
            O => \N__7150\,
            I => \N__7144\
        );

    \I__1248\ : CascadeBuf
    port map (
            O => \N__7147\,
            I => \N__7141\
        );

    \I__1247\ : CascadeBuf
    port map (
            O => \N__7144\,
            I => \N__7138\
        );

    \I__1246\ : CascadeMux
    port map (
            O => \N__7141\,
            I => \N__7135\
        );

    \I__1245\ : CascadeMux
    port map (
            O => \N__7138\,
            I => \N__7132\
        );

    \I__1244\ : CascadeBuf
    port map (
            O => \N__7135\,
            I => \N__7129\
        );

    \I__1243\ : CascadeBuf
    port map (
            O => \N__7132\,
            I => \N__7126\
        );

    \I__1242\ : CascadeMux
    port map (
            O => \N__7129\,
            I => \N__7123\
        );

    \I__1241\ : CascadeMux
    port map (
            O => \N__7126\,
            I => \N__7120\
        );

    \I__1240\ : CascadeBuf
    port map (
            O => \N__7123\,
            I => \N__7117\
        );

    \I__1239\ : CascadeBuf
    port map (
            O => \N__7120\,
            I => \N__7114\
        );

    \I__1238\ : CascadeMux
    port map (
            O => \N__7117\,
            I => \N__7111\
        );

    \I__1237\ : CascadeMux
    port map (
            O => \N__7114\,
            I => \N__7108\
        );

    \I__1236\ : CascadeBuf
    port map (
            O => \N__7111\,
            I => \N__7105\
        );

    \I__1235\ : CascadeBuf
    port map (
            O => \N__7108\,
            I => \N__7102\
        );

    \I__1234\ : CascadeMux
    port map (
            O => \N__7105\,
            I => \N__7099\
        );

    \I__1233\ : CascadeMux
    port map (
            O => \N__7102\,
            I => \N__7096\
        );

    \I__1232\ : CascadeBuf
    port map (
            O => \N__7099\,
            I => \N__7093\
        );

    \I__1231\ : CascadeBuf
    port map (
            O => \N__7096\,
            I => \N__7090\
        );

    \I__1230\ : CascadeMux
    port map (
            O => \N__7093\,
            I => \N__7087\
        );

    \I__1229\ : CascadeMux
    port map (
            O => \N__7090\,
            I => \N__7084\
        );

    \I__1228\ : CascadeBuf
    port map (
            O => \N__7087\,
            I => \N__7081\
        );

    \I__1227\ : CascadeBuf
    port map (
            O => \N__7084\,
            I => \N__7078\
        );

    \I__1226\ : CascadeMux
    port map (
            O => \N__7081\,
            I => \N__7075\
        );

    \I__1225\ : CascadeMux
    port map (
            O => \N__7078\,
            I => \N__7072\
        );

    \I__1224\ : CascadeBuf
    port map (
            O => \N__7075\,
            I => \N__7069\
        );

    \I__1223\ : InMux
    port map (
            O => \N__7072\,
            I => \N__7066\
        );

    \I__1222\ : CascadeMux
    port map (
            O => \N__7069\,
            I => \N__7063\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__7066\,
            I => \N__7060\
        );

    \I__1220\ : InMux
    port map (
            O => \N__7063\,
            I => \N__7057\
        );

    \I__1219\ : Span4Mux_v
    port map (
            O => \N__7060\,
            I => \N__7054\
        );

    \I__1218\ : LocalMux
    port map (
            O => \N__7057\,
            I => \N__7051\
        );

    \I__1217\ : Span4Mux_h
    port map (
            O => \N__7054\,
            I => \N__7048\
        );

    \I__1216\ : Span4Mux_s2_v
    port map (
            O => \N__7051\,
            I => \N__7045\
        );

    \I__1215\ : Sp12to4
    port map (
            O => \N__7048\,
            I => \N__7042\
        );

    \I__1214\ : Span4Mux_v
    port map (
            O => \N__7045\,
            I => \N__7039\
        );

    \I__1213\ : Span12Mux_s10_v
    port map (
            O => \N__7042\,
            I => \N__7036\
        );

    \I__1212\ : Span4Mux_v
    port map (
            O => \N__7039\,
            I => \N__7033\
        );

    \I__1211\ : Span12Mux_h
    port map (
            O => \N__7036\,
            I => \N__7028\
        );

    \I__1210\ : Sp12to4
    port map (
            O => \N__7033\,
            I => \N__7028\
        );

    \I__1209\ : Odrv12
    port map (
            O => \N__7028\,
            I => raddr_c_4
        );

    \I__1208\ : CascadeMux
    port map (
            O => \N__7025\,
            I => \N__7022\
        );

    \I__1207\ : CascadeBuf
    port map (
            O => \N__7022\,
            I => \N__7019\
        );

    \I__1206\ : CascadeMux
    port map (
            O => \N__7019\,
            I => \N__7016\
        );

    \I__1205\ : CascadeBuf
    port map (
            O => \N__7016\,
            I => \N__7012\
        );

    \I__1204\ : CascadeMux
    port map (
            O => \N__7015\,
            I => \N__7009\
        );

    \I__1203\ : CascadeMux
    port map (
            O => \N__7012\,
            I => \N__7006\
        );

    \I__1202\ : CascadeBuf
    port map (
            O => \N__7009\,
            I => \N__7003\
        );

    \I__1201\ : CascadeBuf
    port map (
            O => \N__7006\,
            I => \N__7000\
        );

    \I__1200\ : CascadeMux
    port map (
            O => \N__7003\,
            I => \N__6997\
        );

    \I__1199\ : CascadeMux
    port map (
            O => \N__7000\,
            I => \N__6994\
        );

    \I__1198\ : CascadeBuf
    port map (
            O => \N__6997\,
            I => \N__6991\
        );

    \I__1197\ : CascadeBuf
    port map (
            O => \N__6994\,
            I => \N__6988\
        );

    \I__1196\ : CascadeMux
    port map (
            O => \N__6991\,
            I => \N__6985\
        );

    \I__1195\ : CascadeMux
    port map (
            O => \N__6988\,
            I => \N__6982\
        );

    \I__1194\ : CascadeBuf
    port map (
            O => \N__6985\,
            I => \N__6979\
        );

    \I__1193\ : CascadeBuf
    port map (
            O => \N__6982\,
            I => \N__6976\
        );

    \I__1192\ : CascadeMux
    port map (
            O => \N__6979\,
            I => \N__6973\
        );

    \I__1191\ : CascadeMux
    port map (
            O => \N__6976\,
            I => \N__6970\
        );

    \I__1190\ : CascadeBuf
    port map (
            O => \N__6973\,
            I => \N__6967\
        );

    \I__1189\ : CascadeBuf
    port map (
            O => \N__6970\,
            I => \N__6964\
        );

    \I__1188\ : CascadeMux
    port map (
            O => \N__6967\,
            I => \N__6961\
        );

    \I__1187\ : CascadeMux
    port map (
            O => \N__6964\,
            I => \N__6958\
        );

    \I__1186\ : CascadeBuf
    port map (
            O => \N__6961\,
            I => \N__6955\
        );

    \I__1185\ : CascadeBuf
    port map (
            O => \N__6958\,
            I => \N__6952\
        );

    \I__1184\ : CascadeMux
    port map (
            O => \N__6955\,
            I => \N__6949\
        );

    \I__1183\ : CascadeMux
    port map (
            O => \N__6952\,
            I => \N__6946\
        );

    \I__1182\ : CascadeBuf
    port map (
            O => \N__6949\,
            I => \N__6943\
        );

    \I__1181\ : CascadeBuf
    port map (
            O => \N__6946\,
            I => \N__6940\
        );

    \I__1180\ : CascadeMux
    port map (
            O => \N__6943\,
            I => \N__6937\
        );

    \I__1179\ : CascadeMux
    port map (
            O => \N__6940\,
            I => \N__6934\
        );

    \I__1178\ : CascadeBuf
    port map (
            O => \N__6937\,
            I => \N__6931\
        );

    \I__1177\ : CascadeBuf
    port map (
            O => \N__6934\,
            I => \N__6928\
        );

    \I__1176\ : CascadeMux
    port map (
            O => \N__6931\,
            I => \N__6925\
        );

    \I__1175\ : CascadeMux
    port map (
            O => \N__6928\,
            I => \N__6922\
        );

    \I__1174\ : CascadeBuf
    port map (
            O => \N__6925\,
            I => \N__6919\
        );

    \I__1173\ : CascadeBuf
    port map (
            O => \N__6922\,
            I => \N__6916\
        );

    \I__1172\ : CascadeMux
    port map (
            O => \N__6919\,
            I => \N__6913\
        );

    \I__1171\ : CascadeMux
    port map (
            O => \N__6916\,
            I => \N__6910\
        );

    \I__1170\ : CascadeBuf
    port map (
            O => \N__6913\,
            I => \N__6907\
        );

    \I__1169\ : CascadeBuf
    port map (
            O => \N__6910\,
            I => \N__6904\
        );

    \I__1168\ : CascadeMux
    port map (
            O => \N__6907\,
            I => \N__6901\
        );

    \I__1167\ : CascadeMux
    port map (
            O => \N__6904\,
            I => \N__6898\
        );

    \I__1166\ : CascadeBuf
    port map (
            O => \N__6901\,
            I => \N__6895\
        );

    \I__1165\ : CascadeBuf
    port map (
            O => \N__6898\,
            I => \N__6892\
        );

    \I__1164\ : CascadeMux
    port map (
            O => \N__6895\,
            I => \N__6889\
        );

    \I__1163\ : CascadeMux
    port map (
            O => \N__6892\,
            I => \N__6886\
        );

    \I__1162\ : CascadeBuf
    port map (
            O => \N__6889\,
            I => \N__6883\
        );

    \I__1161\ : CascadeBuf
    port map (
            O => \N__6886\,
            I => \N__6880\
        );

    \I__1160\ : CascadeMux
    port map (
            O => \N__6883\,
            I => \N__6877\
        );

    \I__1159\ : CascadeMux
    port map (
            O => \N__6880\,
            I => \N__6874\
        );

    \I__1158\ : CascadeBuf
    port map (
            O => \N__6877\,
            I => \N__6871\
        );

    \I__1157\ : CascadeBuf
    port map (
            O => \N__6874\,
            I => \N__6868\
        );

    \I__1156\ : CascadeMux
    port map (
            O => \N__6871\,
            I => \N__6865\
        );

    \I__1155\ : CascadeMux
    port map (
            O => \N__6868\,
            I => \N__6862\
        );

    \I__1154\ : CascadeBuf
    port map (
            O => \N__6865\,
            I => \N__6859\
        );

    \I__1153\ : CascadeBuf
    port map (
            O => \N__6862\,
            I => \N__6856\
        );

    \I__1152\ : CascadeMux
    port map (
            O => \N__6859\,
            I => \N__6853\
        );

    \I__1151\ : CascadeMux
    port map (
            O => \N__6856\,
            I => \N__6850\
        );

    \I__1150\ : CascadeBuf
    port map (
            O => \N__6853\,
            I => \N__6847\
        );

    \I__1149\ : InMux
    port map (
            O => \N__6850\,
            I => \N__6844\
        );

    \I__1148\ : CascadeMux
    port map (
            O => \N__6847\,
            I => \N__6841\
        );

    \I__1147\ : LocalMux
    port map (
            O => \N__6844\,
            I => \N__6838\
        );

    \I__1146\ : CascadeBuf
    port map (
            O => \N__6841\,
            I => \N__6835\
        );

    \I__1145\ : Span4Mux_h
    port map (
            O => \N__6838\,
            I => \N__6832\
        );

    \I__1144\ : CascadeMux
    port map (
            O => \N__6835\,
            I => \N__6829\
        );

    \I__1143\ : Span4Mux_h
    port map (
            O => \N__6832\,
            I => \N__6826\
        );

    \I__1142\ : InMux
    port map (
            O => \N__6829\,
            I => \N__6823\
        );

    \I__1141\ : Span4Mux_h
    port map (
            O => \N__6826\,
            I => \N__6820\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__6823\,
            I => \N__6817\
        );

    \I__1139\ : Span4Mux_h
    port map (
            O => \N__6820\,
            I => \N__6812\
        );

    \I__1138\ : Span4Mux_h
    port map (
            O => \N__6817\,
            I => \N__6812\
        );

    \I__1137\ : Odrv4
    port map (
            O => \N__6812\,
            I => waddr_c_9
        );

    \I__1136\ : CascadeMux
    port map (
            O => \N__6809\,
            I => \N__6806\
        );

    \I__1135\ : CascadeBuf
    port map (
            O => \N__6806\,
            I => \N__6803\
        );

    \I__1134\ : CascadeMux
    port map (
            O => \N__6803\,
            I => \N__6800\
        );

    \I__1133\ : CascadeBuf
    port map (
            O => \N__6800\,
            I => \N__6796\
        );

    \I__1132\ : CascadeMux
    port map (
            O => \N__6799\,
            I => \N__6793\
        );

    \I__1131\ : CascadeMux
    port map (
            O => \N__6796\,
            I => \N__6790\
        );

    \I__1130\ : CascadeBuf
    port map (
            O => \N__6793\,
            I => \N__6787\
        );

    \I__1129\ : CascadeBuf
    port map (
            O => \N__6790\,
            I => \N__6784\
        );

    \I__1128\ : CascadeMux
    port map (
            O => \N__6787\,
            I => \N__6781\
        );

    \I__1127\ : CascadeMux
    port map (
            O => \N__6784\,
            I => \N__6778\
        );

    \I__1126\ : CascadeBuf
    port map (
            O => \N__6781\,
            I => \N__6775\
        );

    \I__1125\ : CascadeBuf
    port map (
            O => \N__6778\,
            I => \N__6772\
        );

    \I__1124\ : CascadeMux
    port map (
            O => \N__6775\,
            I => \N__6769\
        );

    \I__1123\ : CascadeMux
    port map (
            O => \N__6772\,
            I => \N__6766\
        );

    \I__1122\ : CascadeBuf
    port map (
            O => \N__6769\,
            I => \N__6763\
        );

    \I__1121\ : CascadeBuf
    port map (
            O => \N__6766\,
            I => \N__6760\
        );

    \I__1120\ : CascadeMux
    port map (
            O => \N__6763\,
            I => \N__6757\
        );

    \I__1119\ : CascadeMux
    port map (
            O => \N__6760\,
            I => \N__6754\
        );

    \I__1118\ : CascadeBuf
    port map (
            O => \N__6757\,
            I => \N__6751\
        );

    \I__1117\ : CascadeBuf
    port map (
            O => \N__6754\,
            I => \N__6748\
        );

    \I__1116\ : CascadeMux
    port map (
            O => \N__6751\,
            I => \N__6745\
        );

    \I__1115\ : CascadeMux
    port map (
            O => \N__6748\,
            I => \N__6742\
        );

    \I__1114\ : CascadeBuf
    port map (
            O => \N__6745\,
            I => \N__6739\
        );

    \I__1113\ : CascadeBuf
    port map (
            O => \N__6742\,
            I => \N__6736\
        );

    \I__1112\ : CascadeMux
    port map (
            O => \N__6739\,
            I => \N__6733\
        );

    \I__1111\ : CascadeMux
    port map (
            O => \N__6736\,
            I => \N__6730\
        );

    \I__1110\ : CascadeBuf
    port map (
            O => \N__6733\,
            I => \N__6727\
        );

    \I__1109\ : CascadeBuf
    port map (
            O => \N__6730\,
            I => \N__6724\
        );

    \I__1108\ : CascadeMux
    port map (
            O => \N__6727\,
            I => \N__6721\
        );

    \I__1107\ : CascadeMux
    port map (
            O => \N__6724\,
            I => \N__6718\
        );

    \I__1106\ : CascadeBuf
    port map (
            O => \N__6721\,
            I => \N__6715\
        );

    \I__1105\ : CascadeBuf
    port map (
            O => \N__6718\,
            I => \N__6712\
        );

    \I__1104\ : CascadeMux
    port map (
            O => \N__6715\,
            I => \N__6709\
        );

    \I__1103\ : CascadeMux
    port map (
            O => \N__6712\,
            I => \N__6706\
        );

    \I__1102\ : CascadeBuf
    port map (
            O => \N__6709\,
            I => \N__6703\
        );

    \I__1101\ : CascadeBuf
    port map (
            O => \N__6706\,
            I => \N__6700\
        );

    \I__1100\ : CascadeMux
    port map (
            O => \N__6703\,
            I => \N__6697\
        );

    \I__1099\ : CascadeMux
    port map (
            O => \N__6700\,
            I => \N__6694\
        );

    \I__1098\ : CascadeBuf
    port map (
            O => \N__6697\,
            I => \N__6691\
        );

    \I__1097\ : CascadeBuf
    port map (
            O => \N__6694\,
            I => \N__6688\
        );

    \I__1096\ : CascadeMux
    port map (
            O => \N__6691\,
            I => \N__6685\
        );

    \I__1095\ : CascadeMux
    port map (
            O => \N__6688\,
            I => \N__6682\
        );

    \I__1094\ : CascadeBuf
    port map (
            O => \N__6685\,
            I => \N__6679\
        );

    \I__1093\ : CascadeBuf
    port map (
            O => \N__6682\,
            I => \N__6676\
        );

    \I__1092\ : CascadeMux
    port map (
            O => \N__6679\,
            I => \N__6673\
        );

    \I__1091\ : CascadeMux
    port map (
            O => \N__6676\,
            I => \N__6670\
        );

    \I__1090\ : CascadeBuf
    port map (
            O => \N__6673\,
            I => \N__6667\
        );

    \I__1089\ : CascadeBuf
    port map (
            O => \N__6670\,
            I => \N__6664\
        );

    \I__1088\ : CascadeMux
    port map (
            O => \N__6667\,
            I => \N__6661\
        );

    \I__1087\ : CascadeMux
    port map (
            O => \N__6664\,
            I => \N__6658\
        );

    \I__1086\ : CascadeBuf
    port map (
            O => \N__6661\,
            I => \N__6655\
        );

    \I__1085\ : CascadeBuf
    port map (
            O => \N__6658\,
            I => \N__6652\
        );

    \I__1084\ : CascadeMux
    port map (
            O => \N__6655\,
            I => \N__6649\
        );

    \I__1083\ : CascadeMux
    port map (
            O => \N__6652\,
            I => \N__6646\
        );

    \I__1082\ : CascadeBuf
    port map (
            O => \N__6649\,
            I => \N__6643\
        );

    \I__1081\ : CascadeBuf
    port map (
            O => \N__6646\,
            I => \N__6640\
        );

    \I__1080\ : CascadeMux
    port map (
            O => \N__6643\,
            I => \N__6637\
        );

    \I__1079\ : CascadeMux
    port map (
            O => \N__6640\,
            I => \N__6634\
        );

    \I__1078\ : CascadeBuf
    port map (
            O => \N__6637\,
            I => \N__6631\
        );

    \I__1077\ : InMux
    port map (
            O => \N__6634\,
            I => \N__6628\
        );

    \I__1076\ : CascadeMux
    port map (
            O => \N__6631\,
            I => \N__6625\
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__6628\,
            I => \N__6622\
        );

    \I__1074\ : CascadeBuf
    port map (
            O => \N__6625\,
            I => \N__6619\
        );

    \I__1073\ : Span4Mux_s2_v
    port map (
            O => \N__6622\,
            I => \N__6616\
        );

    \I__1072\ : CascadeMux
    port map (
            O => \N__6619\,
            I => \N__6613\
        );

    \I__1071\ : Span4Mux_h
    port map (
            O => \N__6616\,
            I => \N__6610\
        );

    \I__1070\ : InMux
    port map (
            O => \N__6613\,
            I => \N__6607\
        );

    \I__1069\ : Sp12to4
    port map (
            O => \N__6610\,
            I => \N__6604\
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__6607\,
            I => \N__6601\
        );

    \I__1067\ : Span12Mux_h
    port map (
            O => \N__6604\,
            I => \N__6596\
        );

    \I__1066\ : Span12Mux_s2_v
    port map (
            O => \N__6601\,
            I => \N__6596\
        );

    \I__1065\ : Odrv12
    port map (
            O => \N__6596\,
            I => raddr_c_9
        );

    \I__1064\ : CascadeMux
    port map (
            O => \N__6593\,
            I => \N__6590\
        );

    \I__1063\ : CascadeBuf
    port map (
            O => \N__6590\,
            I => \N__6587\
        );

    \I__1062\ : CascadeMux
    port map (
            O => \N__6587\,
            I => \N__6584\
        );

    \I__1061\ : CascadeBuf
    port map (
            O => \N__6584\,
            I => \N__6580\
        );

    \I__1060\ : CascadeMux
    port map (
            O => \N__6583\,
            I => \N__6577\
        );

    \I__1059\ : CascadeMux
    port map (
            O => \N__6580\,
            I => \N__6574\
        );

    \I__1058\ : CascadeBuf
    port map (
            O => \N__6577\,
            I => \N__6571\
        );

    \I__1057\ : CascadeBuf
    port map (
            O => \N__6574\,
            I => \N__6568\
        );

    \I__1056\ : CascadeMux
    port map (
            O => \N__6571\,
            I => \N__6565\
        );

    \I__1055\ : CascadeMux
    port map (
            O => \N__6568\,
            I => \N__6562\
        );

    \I__1054\ : CascadeBuf
    port map (
            O => \N__6565\,
            I => \N__6559\
        );

    \I__1053\ : CascadeBuf
    port map (
            O => \N__6562\,
            I => \N__6556\
        );

    \I__1052\ : CascadeMux
    port map (
            O => \N__6559\,
            I => \N__6553\
        );

    \I__1051\ : CascadeMux
    port map (
            O => \N__6556\,
            I => \N__6550\
        );

    \I__1050\ : CascadeBuf
    port map (
            O => \N__6553\,
            I => \N__6547\
        );

    \I__1049\ : CascadeBuf
    port map (
            O => \N__6550\,
            I => \N__6544\
        );

    \I__1048\ : CascadeMux
    port map (
            O => \N__6547\,
            I => \N__6541\
        );

    \I__1047\ : CascadeMux
    port map (
            O => \N__6544\,
            I => \N__6538\
        );

    \I__1046\ : CascadeBuf
    port map (
            O => \N__6541\,
            I => \N__6535\
        );

    \I__1045\ : CascadeBuf
    port map (
            O => \N__6538\,
            I => \N__6532\
        );

    \I__1044\ : CascadeMux
    port map (
            O => \N__6535\,
            I => \N__6529\
        );

    \I__1043\ : CascadeMux
    port map (
            O => \N__6532\,
            I => \N__6526\
        );

    \I__1042\ : CascadeBuf
    port map (
            O => \N__6529\,
            I => \N__6523\
        );

    \I__1041\ : CascadeBuf
    port map (
            O => \N__6526\,
            I => \N__6520\
        );

    \I__1040\ : CascadeMux
    port map (
            O => \N__6523\,
            I => \N__6517\
        );

    \I__1039\ : CascadeMux
    port map (
            O => \N__6520\,
            I => \N__6514\
        );

    \I__1038\ : CascadeBuf
    port map (
            O => \N__6517\,
            I => \N__6511\
        );

    \I__1037\ : CascadeBuf
    port map (
            O => \N__6514\,
            I => \N__6508\
        );

    \I__1036\ : CascadeMux
    port map (
            O => \N__6511\,
            I => \N__6505\
        );

    \I__1035\ : CascadeMux
    port map (
            O => \N__6508\,
            I => \N__6502\
        );

    \I__1034\ : CascadeBuf
    port map (
            O => \N__6505\,
            I => \N__6499\
        );

    \I__1033\ : CascadeBuf
    port map (
            O => \N__6502\,
            I => \N__6496\
        );

    \I__1032\ : CascadeMux
    port map (
            O => \N__6499\,
            I => \N__6493\
        );

    \I__1031\ : CascadeMux
    port map (
            O => \N__6496\,
            I => \N__6490\
        );

    \I__1030\ : CascadeBuf
    port map (
            O => \N__6493\,
            I => \N__6487\
        );

    \I__1029\ : CascadeBuf
    port map (
            O => \N__6490\,
            I => \N__6484\
        );

    \I__1028\ : CascadeMux
    port map (
            O => \N__6487\,
            I => \N__6481\
        );

    \I__1027\ : CascadeMux
    port map (
            O => \N__6484\,
            I => \N__6478\
        );

    \I__1026\ : CascadeBuf
    port map (
            O => \N__6481\,
            I => \N__6475\
        );

    \I__1025\ : CascadeBuf
    port map (
            O => \N__6478\,
            I => \N__6472\
        );

    \I__1024\ : CascadeMux
    port map (
            O => \N__6475\,
            I => \N__6469\
        );

    \I__1023\ : CascadeMux
    port map (
            O => \N__6472\,
            I => \N__6466\
        );

    \I__1022\ : CascadeBuf
    port map (
            O => \N__6469\,
            I => \N__6463\
        );

    \I__1021\ : CascadeBuf
    port map (
            O => \N__6466\,
            I => \N__6460\
        );

    \I__1020\ : CascadeMux
    port map (
            O => \N__6463\,
            I => \N__6457\
        );

    \I__1019\ : CascadeMux
    port map (
            O => \N__6460\,
            I => \N__6454\
        );

    \I__1018\ : CascadeBuf
    port map (
            O => \N__6457\,
            I => \N__6451\
        );

    \I__1017\ : CascadeBuf
    port map (
            O => \N__6454\,
            I => \N__6448\
        );

    \I__1016\ : CascadeMux
    port map (
            O => \N__6451\,
            I => \N__6445\
        );

    \I__1015\ : CascadeMux
    port map (
            O => \N__6448\,
            I => \N__6442\
        );

    \I__1014\ : CascadeBuf
    port map (
            O => \N__6445\,
            I => \N__6439\
        );

    \I__1013\ : CascadeBuf
    port map (
            O => \N__6442\,
            I => \N__6436\
        );

    \I__1012\ : CascadeMux
    port map (
            O => \N__6439\,
            I => \N__6433\
        );

    \I__1011\ : CascadeMux
    port map (
            O => \N__6436\,
            I => \N__6430\
        );

    \I__1010\ : CascadeBuf
    port map (
            O => \N__6433\,
            I => \N__6427\
        );

    \I__1009\ : CascadeBuf
    port map (
            O => \N__6430\,
            I => \N__6424\
        );

    \I__1008\ : CascadeMux
    port map (
            O => \N__6427\,
            I => \N__6421\
        );

    \I__1007\ : CascadeMux
    port map (
            O => \N__6424\,
            I => \N__6418\
        );

    \I__1006\ : CascadeBuf
    port map (
            O => \N__6421\,
            I => \N__6415\
        );

    \I__1005\ : InMux
    port map (
            O => \N__6418\,
            I => \N__6412\
        );

    \I__1004\ : CascadeMux
    port map (
            O => \N__6415\,
            I => \N__6409\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__6412\,
            I => \N__6406\
        );

    \I__1002\ : CascadeBuf
    port map (
            O => \N__6409\,
            I => \N__6403\
        );

    \I__1001\ : Span4Mux_h
    port map (
            O => \N__6406\,
            I => \N__6400\
        );

    \I__1000\ : CascadeMux
    port map (
            O => \N__6403\,
            I => \N__6397\
        );

    \I__999\ : Span4Mux_h
    port map (
            O => \N__6400\,
            I => \N__6394\
        );

    \I__998\ : InMux
    port map (
            O => \N__6397\,
            I => \N__6391\
        );

    \I__997\ : Span4Mux_h
    port map (
            O => \N__6394\,
            I => \N__6388\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__6391\,
            I => \N__6385\
        );

    \I__995\ : Span4Mux_h
    port map (
            O => \N__6388\,
            I => \N__6380\
        );

    \I__994\ : Span4Mux_h
    port map (
            O => \N__6385\,
            I => \N__6380\
        );

    \I__993\ : Odrv4
    port map (
            O => \N__6380\,
            I => waddr_c_7
        );

    \I__992\ : CascadeMux
    port map (
            O => \N__6377\,
            I => \N__6374\
        );

    \I__991\ : CascadeBuf
    port map (
            O => \N__6374\,
            I => \N__6371\
        );

    \I__990\ : CascadeMux
    port map (
            O => \N__6371\,
            I => \N__6368\
        );

    \I__989\ : CascadeBuf
    port map (
            O => \N__6368\,
            I => \N__6364\
        );

    \I__988\ : CascadeMux
    port map (
            O => \N__6367\,
            I => \N__6361\
        );

    \I__987\ : CascadeMux
    port map (
            O => \N__6364\,
            I => \N__6358\
        );

    \I__986\ : CascadeBuf
    port map (
            O => \N__6361\,
            I => \N__6355\
        );

    \I__985\ : CascadeBuf
    port map (
            O => \N__6358\,
            I => \N__6352\
        );

    \I__984\ : CascadeMux
    port map (
            O => \N__6355\,
            I => \N__6349\
        );

    \I__983\ : CascadeMux
    port map (
            O => \N__6352\,
            I => \N__6346\
        );

    \I__982\ : CascadeBuf
    port map (
            O => \N__6349\,
            I => \N__6343\
        );

    \I__981\ : CascadeBuf
    port map (
            O => \N__6346\,
            I => \N__6340\
        );

    \I__980\ : CascadeMux
    port map (
            O => \N__6343\,
            I => \N__6337\
        );

    \I__979\ : CascadeMux
    port map (
            O => \N__6340\,
            I => \N__6334\
        );

    \I__978\ : CascadeBuf
    port map (
            O => \N__6337\,
            I => \N__6331\
        );

    \I__977\ : CascadeBuf
    port map (
            O => \N__6334\,
            I => \N__6328\
        );

    \I__976\ : CascadeMux
    port map (
            O => \N__6331\,
            I => \N__6325\
        );

    \I__975\ : CascadeMux
    port map (
            O => \N__6328\,
            I => \N__6322\
        );

    \I__974\ : CascadeBuf
    port map (
            O => \N__6325\,
            I => \N__6319\
        );

    \I__973\ : CascadeBuf
    port map (
            O => \N__6322\,
            I => \N__6316\
        );

    \I__972\ : CascadeMux
    port map (
            O => \N__6319\,
            I => \N__6313\
        );

    \I__971\ : CascadeMux
    port map (
            O => \N__6316\,
            I => \N__6310\
        );

    \I__970\ : CascadeBuf
    port map (
            O => \N__6313\,
            I => \N__6307\
        );

    \I__969\ : CascadeBuf
    port map (
            O => \N__6310\,
            I => \N__6304\
        );

    \I__968\ : CascadeMux
    port map (
            O => \N__6307\,
            I => \N__6301\
        );

    \I__967\ : CascadeMux
    port map (
            O => \N__6304\,
            I => \N__6298\
        );

    \I__966\ : CascadeBuf
    port map (
            O => \N__6301\,
            I => \N__6295\
        );

    \I__965\ : CascadeBuf
    port map (
            O => \N__6298\,
            I => \N__6292\
        );

    \I__964\ : CascadeMux
    port map (
            O => \N__6295\,
            I => \N__6289\
        );

    \I__963\ : CascadeMux
    port map (
            O => \N__6292\,
            I => \N__6286\
        );

    \I__962\ : CascadeBuf
    port map (
            O => \N__6289\,
            I => \N__6283\
        );

    \I__961\ : CascadeBuf
    port map (
            O => \N__6286\,
            I => \N__6280\
        );

    \I__960\ : CascadeMux
    port map (
            O => \N__6283\,
            I => \N__6277\
        );

    \I__959\ : CascadeMux
    port map (
            O => \N__6280\,
            I => \N__6274\
        );

    \I__958\ : CascadeBuf
    port map (
            O => \N__6277\,
            I => \N__6271\
        );

    \I__957\ : CascadeBuf
    port map (
            O => \N__6274\,
            I => \N__6268\
        );

    \I__956\ : CascadeMux
    port map (
            O => \N__6271\,
            I => \N__6265\
        );

    \I__955\ : CascadeMux
    port map (
            O => \N__6268\,
            I => \N__6262\
        );

    \I__954\ : CascadeBuf
    port map (
            O => \N__6265\,
            I => \N__6259\
        );

    \I__953\ : CascadeBuf
    port map (
            O => \N__6262\,
            I => \N__6256\
        );

    \I__952\ : CascadeMux
    port map (
            O => \N__6259\,
            I => \N__6253\
        );

    \I__951\ : CascadeMux
    port map (
            O => \N__6256\,
            I => \N__6250\
        );

    \I__950\ : CascadeBuf
    port map (
            O => \N__6253\,
            I => \N__6247\
        );

    \I__949\ : CascadeBuf
    port map (
            O => \N__6250\,
            I => \N__6244\
        );

    \I__948\ : CascadeMux
    port map (
            O => \N__6247\,
            I => \N__6241\
        );

    \I__947\ : CascadeMux
    port map (
            O => \N__6244\,
            I => \N__6238\
        );

    \I__946\ : CascadeBuf
    port map (
            O => \N__6241\,
            I => \N__6235\
        );

    \I__945\ : CascadeBuf
    port map (
            O => \N__6238\,
            I => \N__6232\
        );

    \I__944\ : CascadeMux
    port map (
            O => \N__6235\,
            I => \N__6229\
        );

    \I__943\ : CascadeMux
    port map (
            O => \N__6232\,
            I => \N__6226\
        );

    \I__942\ : CascadeBuf
    port map (
            O => \N__6229\,
            I => \N__6223\
        );

    \I__941\ : CascadeBuf
    port map (
            O => \N__6226\,
            I => \N__6220\
        );

    \I__940\ : CascadeMux
    port map (
            O => \N__6223\,
            I => \N__6217\
        );

    \I__939\ : CascadeMux
    port map (
            O => \N__6220\,
            I => \N__6214\
        );

    \I__938\ : CascadeBuf
    port map (
            O => \N__6217\,
            I => \N__6211\
        );

    \I__937\ : CascadeBuf
    port map (
            O => \N__6214\,
            I => \N__6208\
        );

    \I__936\ : CascadeMux
    port map (
            O => \N__6211\,
            I => \N__6205\
        );

    \I__935\ : CascadeMux
    port map (
            O => \N__6208\,
            I => \N__6202\
        );

    \I__934\ : CascadeBuf
    port map (
            O => \N__6205\,
            I => \N__6199\
        );

    \I__933\ : InMux
    port map (
            O => \N__6202\,
            I => \N__6196\
        );

    \I__932\ : CascadeMux
    port map (
            O => \N__6199\,
            I => \N__6193\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__6196\,
            I => \N__6190\
        );

    \I__930\ : CascadeBuf
    port map (
            O => \N__6193\,
            I => \N__6187\
        );

    \I__929\ : Span4Mux_v
    port map (
            O => \N__6190\,
            I => \N__6184\
        );

    \I__928\ : CascadeMux
    port map (
            O => \N__6187\,
            I => \N__6181\
        );

    \I__927\ : Sp12to4
    port map (
            O => \N__6184\,
            I => \N__6178\
        );

    \I__926\ : InMux
    port map (
            O => \N__6181\,
            I => \N__6175\
        );

    \I__925\ : Span12Mux_h
    port map (
            O => \N__6178\,
            I => \N__6172\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__6175\,
            I => \N__6169\
        );

    \I__923\ : Span12Mux_v
    port map (
            O => \N__6172\,
            I => \N__6166\
        );

    \I__922\ : Span12Mux_v
    port map (
            O => \N__6169\,
            I => \N__6163\
        );

    \I__921\ : Odrv12
    port map (
            O => \N__6166\,
            I => raddr_c_0
        );

    \I__920\ : Odrv12
    port map (
            O => \N__6163\,
            I => raddr_c_0
        );

    \I__919\ : CascadeMux
    port map (
            O => \N__6158\,
            I => \N__6155\
        );

    \I__918\ : CascadeBuf
    port map (
            O => \N__6155\,
            I => \N__6152\
        );

    \I__917\ : CascadeMux
    port map (
            O => \N__6152\,
            I => \N__6149\
        );

    \I__916\ : CascadeBuf
    port map (
            O => \N__6149\,
            I => \N__6146\
        );

    \I__915\ : CascadeMux
    port map (
            O => \N__6146\,
            I => \N__6142\
        );

    \I__914\ : CascadeMux
    port map (
            O => \N__6145\,
            I => \N__6139\
        );

    \I__913\ : CascadeBuf
    port map (
            O => \N__6142\,
            I => \N__6136\
        );

    \I__912\ : CascadeBuf
    port map (
            O => \N__6139\,
            I => \N__6133\
        );

    \I__911\ : CascadeMux
    port map (
            O => \N__6136\,
            I => \N__6130\
        );

    \I__910\ : CascadeMux
    port map (
            O => \N__6133\,
            I => \N__6127\
        );

    \I__909\ : CascadeBuf
    port map (
            O => \N__6130\,
            I => \N__6124\
        );

    \I__908\ : CascadeBuf
    port map (
            O => \N__6127\,
            I => \N__6121\
        );

    \I__907\ : CascadeMux
    port map (
            O => \N__6124\,
            I => \N__6118\
        );

    \I__906\ : CascadeMux
    port map (
            O => \N__6121\,
            I => \N__6115\
        );

    \I__905\ : CascadeBuf
    port map (
            O => \N__6118\,
            I => \N__6112\
        );

    \I__904\ : CascadeBuf
    port map (
            O => \N__6115\,
            I => \N__6109\
        );

    \I__903\ : CascadeMux
    port map (
            O => \N__6112\,
            I => \N__6106\
        );

    \I__902\ : CascadeMux
    port map (
            O => \N__6109\,
            I => \N__6103\
        );

    \I__901\ : CascadeBuf
    port map (
            O => \N__6106\,
            I => \N__6100\
        );

    \I__900\ : CascadeBuf
    port map (
            O => \N__6103\,
            I => \N__6097\
        );

    \I__899\ : CascadeMux
    port map (
            O => \N__6100\,
            I => \N__6094\
        );

    \I__898\ : CascadeMux
    port map (
            O => \N__6097\,
            I => \N__6091\
        );

    \I__897\ : CascadeBuf
    port map (
            O => \N__6094\,
            I => \N__6088\
        );

    \I__896\ : CascadeBuf
    port map (
            O => \N__6091\,
            I => \N__6085\
        );

    \I__895\ : CascadeMux
    port map (
            O => \N__6088\,
            I => \N__6082\
        );

    \I__894\ : CascadeMux
    port map (
            O => \N__6085\,
            I => \N__6079\
        );

    \I__893\ : CascadeBuf
    port map (
            O => \N__6082\,
            I => \N__6076\
        );

    \I__892\ : CascadeBuf
    port map (
            O => \N__6079\,
            I => \N__6073\
        );

    \I__891\ : CascadeMux
    port map (
            O => \N__6076\,
            I => \N__6070\
        );

    \I__890\ : CascadeMux
    port map (
            O => \N__6073\,
            I => \N__6067\
        );

    \I__889\ : CascadeBuf
    port map (
            O => \N__6070\,
            I => \N__6064\
        );

    \I__888\ : CascadeBuf
    port map (
            O => \N__6067\,
            I => \N__6061\
        );

    \I__887\ : CascadeMux
    port map (
            O => \N__6064\,
            I => \N__6058\
        );

    \I__886\ : CascadeMux
    port map (
            O => \N__6061\,
            I => \N__6055\
        );

    \I__885\ : CascadeBuf
    port map (
            O => \N__6058\,
            I => \N__6052\
        );

    \I__884\ : CascadeBuf
    port map (
            O => \N__6055\,
            I => \N__6049\
        );

    \I__883\ : CascadeMux
    port map (
            O => \N__6052\,
            I => \N__6046\
        );

    \I__882\ : CascadeMux
    port map (
            O => \N__6049\,
            I => \N__6043\
        );

    \I__881\ : CascadeBuf
    port map (
            O => \N__6046\,
            I => \N__6040\
        );

    \I__880\ : CascadeBuf
    port map (
            O => \N__6043\,
            I => \N__6037\
        );

    \I__879\ : CascadeMux
    port map (
            O => \N__6040\,
            I => \N__6034\
        );

    \I__878\ : CascadeMux
    port map (
            O => \N__6037\,
            I => \N__6031\
        );

    \I__877\ : CascadeBuf
    port map (
            O => \N__6034\,
            I => \N__6028\
        );

    \I__876\ : CascadeBuf
    port map (
            O => \N__6031\,
            I => \N__6025\
        );

    \I__875\ : CascadeMux
    port map (
            O => \N__6028\,
            I => \N__6022\
        );

    \I__874\ : CascadeMux
    port map (
            O => \N__6025\,
            I => \N__6019\
        );

    \I__873\ : CascadeBuf
    port map (
            O => \N__6022\,
            I => \N__6016\
        );

    \I__872\ : CascadeBuf
    port map (
            O => \N__6019\,
            I => \N__6013\
        );

    \I__871\ : CascadeMux
    port map (
            O => \N__6016\,
            I => \N__6010\
        );

    \I__870\ : CascadeMux
    port map (
            O => \N__6013\,
            I => \N__6007\
        );

    \I__869\ : CascadeBuf
    port map (
            O => \N__6010\,
            I => \N__6004\
        );

    \I__868\ : CascadeBuf
    port map (
            O => \N__6007\,
            I => \N__6001\
        );

    \I__867\ : CascadeMux
    port map (
            O => \N__6004\,
            I => \N__5998\
        );

    \I__866\ : CascadeMux
    port map (
            O => \N__6001\,
            I => \N__5995\
        );

    \I__865\ : CascadeBuf
    port map (
            O => \N__5998\,
            I => \N__5992\
        );

    \I__864\ : CascadeBuf
    port map (
            O => \N__5995\,
            I => \N__5989\
        );

    \I__863\ : CascadeMux
    port map (
            O => \N__5992\,
            I => \N__5986\
        );

    \I__862\ : CascadeMux
    port map (
            O => \N__5989\,
            I => \N__5983\
        );

    \I__861\ : InMux
    port map (
            O => \N__5986\,
            I => \N__5980\
        );

    \I__860\ : CascadeBuf
    port map (
            O => \N__5983\,
            I => \N__5977\
        );

    \I__859\ : LocalMux
    port map (
            O => \N__5980\,
            I => \N__5974\
        );

    \I__858\ : CascadeMux
    port map (
            O => \N__5977\,
            I => \N__5971\
        );

    \I__857\ : Span4Mux_h
    port map (
            O => \N__5974\,
            I => \N__5968\
        );

    \I__856\ : CascadeBuf
    port map (
            O => \N__5971\,
            I => \N__5965\
        );

    \I__855\ : Span4Mux_h
    port map (
            O => \N__5968\,
            I => \N__5962\
        );

    \I__854\ : CascadeMux
    port map (
            O => \N__5965\,
            I => \N__5959\
        );

    \I__853\ : Span4Mux_h
    port map (
            O => \N__5962\,
            I => \N__5956\
        );

    \I__852\ : InMux
    port map (
            O => \N__5959\,
            I => \N__5953\
        );

    \I__851\ : Span4Mux_h
    port map (
            O => \N__5956\,
            I => \N__5948\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__5953\,
            I => \N__5948\
        );

    \I__849\ : Span4Mux_h
    port map (
            O => \N__5948\,
            I => \N__5945\
        );

    \I__848\ : Span4Mux_h
    port map (
            O => \N__5945\,
            I => \N__5942\
        );

    \I__847\ : Odrv4
    port map (
            O => \N__5942\,
            I => waddr_c_10
        );

    \I__846\ : CascadeMux
    port map (
            O => \N__5939\,
            I => \N__5936\
        );

    \I__845\ : CascadeBuf
    port map (
            O => \N__5936\,
            I => \N__5933\
        );

    \I__844\ : CascadeMux
    port map (
            O => \N__5933\,
            I => \N__5930\
        );

    \I__843\ : CascadeBuf
    port map (
            O => \N__5930\,
            I => \N__5926\
        );

    \I__842\ : CascadeMux
    port map (
            O => \N__5929\,
            I => \N__5923\
        );

    \I__841\ : CascadeMux
    port map (
            O => \N__5926\,
            I => \N__5920\
        );

    \I__840\ : CascadeBuf
    port map (
            O => \N__5923\,
            I => \N__5917\
        );

    \I__839\ : CascadeBuf
    port map (
            O => \N__5920\,
            I => \N__5914\
        );

    \I__838\ : CascadeMux
    port map (
            O => \N__5917\,
            I => \N__5911\
        );

    \I__837\ : CascadeMux
    port map (
            O => \N__5914\,
            I => \N__5908\
        );

    \I__836\ : CascadeBuf
    port map (
            O => \N__5911\,
            I => \N__5905\
        );

    \I__835\ : CascadeBuf
    port map (
            O => \N__5908\,
            I => \N__5902\
        );

    \I__834\ : CascadeMux
    port map (
            O => \N__5905\,
            I => \N__5899\
        );

    \I__833\ : CascadeMux
    port map (
            O => \N__5902\,
            I => \N__5896\
        );

    \I__832\ : CascadeBuf
    port map (
            O => \N__5899\,
            I => \N__5893\
        );

    \I__831\ : CascadeBuf
    port map (
            O => \N__5896\,
            I => \N__5890\
        );

    \I__830\ : CascadeMux
    port map (
            O => \N__5893\,
            I => \N__5887\
        );

    \I__829\ : CascadeMux
    port map (
            O => \N__5890\,
            I => \N__5884\
        );

    \I__828\ : CascadeBuf
    port map (
            O => \N__5887\,
            I => \N__5881\
        );

    \I__827\ : CascadeBuf
    port map (
            O => \N__5884\,
            I => \N__5878\
        );

    \I__826\ : CascadeMux
    port map (
            O => \N__5881\,
            I => \N__5875\
        );

    \I__825\ : CascadeMux
    port map (
            O => \N__5878\,
            I => \N__5872\
        );

    \I__824\ : CascadeBuf
    port map (
            O => \N__5875\,
            I => \N__5869\
        );

    \I__823\ : CascadeBuf
    port map (
            O => \N__5872\,
            I => \N__5866\
        );

    \I__822\ : CascadeMux
    port map (
            O => \N__5869\,
            I => \N__5863\
        );

    \I__821\ : CascadeMux
    port map (
            O => \N__5866\,
            I => \N__5860\
        );

    \I__820\ : CascadeBuf
    port map (
            O => \N__5863\,
            I => \N__5857\
        );

    \I__819\ : CascadeBuf
    port map (
            O => \N__5860\,
            I => \N__5854\
        );

    \I__818\ : CascadeMux
    port map (
            O => \N__5857\,
            I => \N__5851\
        );

    \I__817\ : CascadeMux
    port map (
            O => \N__5854\,
            I => \N__5848\
        );

    \I__816\ : CascadeBuf
    port map (
            O => \N__5851\,
            I => \N__5845\
        );

    \I__815\ : CascadeBuf
    port map (
            O => \N__5848\,
            I => \N__5842\
        );

    \I__814\ : CascadeMux
    port map (
            O => \N__5845\,
            I => \N__5839\
        );

    \I__813\ : CascadeMux
    port map (
            O => \N__5842\,
            I => \N__5836\
        );

    \I__812\ : CascadeBuf
    port map (
            O => \N__5839\,
            I => \N__5833\
        );

    \I__811\ : CascadeBuf
    port map (
            O => \N__5836\,
            I => \N__5830\
        );

    \I__810\ : CascadeMux
    port map (
            O => \N__5833\,
            I => \N__5827\
        );

    \I__809\ : CascadeMux
    port map (
            O => \N__5830\,
            I => \N__5824\
        );

    \I__808\ : CascadeBuf
    port map (
            O => \N__5827\,
            I => \N__5821\
        );

    \I__807\ : CascadeBuf
    port map (
            O => \N__5824\,
            I => \N__5818\
        );

    \I__806\ : CascadeMux
    port map (
            O => \N__5821\,
            I => \N__5815\
        );

    \I__805\ : CascadeMux
    port map (
            O => \N__5818\,
            I => \N__5812\
        );

    \I__804\ : CascadeBuf
    port map (
            O => \N__5815\,
            I => \N__5809\
        );

    \I__803\ : CascadeBuf
    port map (
            O => \N__5812\,
            I => \N__5806\
        );

    \I__802\ : CascadeMux
    port map (
            O => \N__5809\,
            I => \N__5803\
        );

    \I__801\ : CascadeMux
    port map (
            O => \N__5806\,
            I => \N__5800\
        );

    \I__800\ : CascadeBuf
    port map (
            O => \N__5803\,
            I => \N__5797\
        );

    \I__799\ : CascadeBuf
    port map (
            O => \N__5800\,
            I => \N__5794\
        );

    \I__798\ : CascadeMux
    port map (
            O => \N__5797\,
            I => \N__5791\
        );

    \I__797\ : CascadeMux
    port map (
            O => \N__5794\,
            I => \N__5788\
        );

    \I__796\ : CascadeBuf
    port map (
            O => \N__5791\,
            I => \N__5785\
        );

    \I__795\ : CascadeBuf
    port map (
            O => \N__5788\,
            I => \N__5782\
        );

    \I__794\ : CascadeMux
    port map (
            O => \N__5785\,
            I => \N__5779\
        );

    \I__793\ : CascadeMux
    port map (
            O => \N__5782\,
            I => \N__5776\
        );

    \I__792\ : CascadeBuf
    port map (
            O => \N__5779\,
            I => \N__5773\
        );

    \I__791\ : CascadeBuf
    port map (
            O => \N__5776\,
            I => \N__5770\
        );

    \I__790\ : CascadeMux
    port map (
            O => \N__5773\,
            I => \N__5767\
        );

    \I__789\ : CascadeMux
    port map (
            O => \N__5770\,
            I => \N__5764\
        );

    \I__788\ : CascadeBuf
    port map (
            O => \N__5767\,
            I => \N__5761\
        );

    \I__787\ : InMux
    port map (
            O => \N__5764\,
            I => \N__5758\
        );

    \I__786\ : CascadeMux
    port map (
            O => \N__5761\,
            I => \N__5755\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__5758\,
            I => \N__5752\
        );

    \I__784\ : CascadeBuf
    port map (
            O => \N__5755\,
            I => \N__5749\
        );

    \I__783\ : Span4Mux_h
    port map (
            O => \N__5752\,
            I => \N__5746\
        );

    \I__782\ : CascadeMux
    port map (
            O => \N__5749\,
            I => \N__5743\
        );

    \I__781\ : Span4Mux_h
    port map (
            O => \N__5746\,
            I => \N__5740\
        );

    \I__780\ : InMux
    port map (
            O => \N__5743\,
            I => \N__5737\
        );

    \I__779\ : Span4Mux_h
    port map (
            O => \N__5740\,
            I => \N__5734\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__5737\,
            I => \N__5731\
        );

    \I__777\ : Span4Mux_h
    port map (
            O => \N__5734\,
            I => \N__5726\
        );

    \I__776\ : Span4Mux_h
    port map (
            O => \N__5731\,
            I => \N__5726\
        );

    \I__775\ : Odrv4
    port map (
            O => \N__5726\,
            I => waddr_c_8
        );

    \I__774\ : CascadeMux
    port map (
            O => \N__5723\,
            I => \N__5720\
        );

    \I__773\ : CascadeBuf
    port map (
            O => \N__5720\,
            I => \N__5716\
        );

    \I__772\ : CascadeMux
    port map (
            O => \N__5719\,
            I => \N__5713\
        );

    \I__771\ : CascadeMux
    port map (
            O => \N__5716\,
            I => \N__5710\
        );

    \I__770\ : CascadeBuf
    port map (
            O => \N__5713\,
            I => \N__5707\
        );

    \I__769\ : CascadeBuf
    port map (
            O => \N__5710\,
            I => \N__5704\
        );

    \I__768\ : CascadeMux
    port map (
            O => \N__5707\,
            I => \N__5701\
        );

    \I__767\ : CascadeMux
    port map (
            O => \N__5704\,
            I => \N__5698\
        );

    \I__766\ : CascadeBuf
    port map (
            O => \N__5701\,
            I => \N__5695\
        );

    \I__765\ : CascadeBuf
    port map (
            O => \N__5698\,
            I => \N__5692\
        );

    \I__764\ : CascadeMux
    port map (
            O => \N__5695\,
            I => \N__5689\
        );

    \I__763\ : CascadeMux
    port map (
            O => \N__5692\,
            I => \N__5686\
        );

    \I__762\ : CascadeBuf
    port map (
            O => \N__5689\,
            I => \N__5683\
        );

    \I__761\ : CascadeBuf
    port map (
            O => \N__5686\,
            I => \N__5680\
        );

    \I__760\ : CascadeMux
    port map (
            O => \N__5683\,
            I => \N__5677\
        );

    \I__759\ : CascadeMux
    port map (
            O => \N__5680\,
            I => \N__5674\
        );

    \I__758\ : CascadeBuf
    port map (
            O => \N__5677\,
            I => \N__5671\
        );

    \I__757\ : CascadeBuf
    port map (
            O => \N__5674\,
            I => \N__5668\
        );

    \I__756\ : CascadeMux
    port map (
            O => \N__5671\,
            I => \N__5665\
        );

    \I__755\ : CascadeMux
    port map (
            O => \N__5668\,
            I => \N__5662\
        );

    \I__754\ : CascadeBuf
    port map (
            O => \N__5665\,
            I => \N__5659\
        );

    \I__753\ : CascadeBuf
    port map (
            O => \N__5662\,
            I => \N__5656\
        );

    \I__752\ : CascadeMux
    port map (
            O => \N__5659\,
            I => \N__5653\
        );

    \I__751\ : CascadeMux
    port map (
            O => \N__5656\,
            I => \N__5650\
        );

    \I__750\ : CascadeBuf
    port map (
            O => \N__5653\,
            I => \N__5647\
        );

    \I__749\ : CascadeBuf
    port map (
            O => \N__5650\,
            I => \N__5644\
        );

    \I__748\ : CascadeMux
    port map (
            O => \N__5647\,
            I => \N__5641\
        );

    \I__747\ : CascadeMux
    port map (
            O => \N__5644\,
            I => \N__5638\
        );

    \I__746\ : CascadeBuf
    port map (
            O => \N__5641\,
            I => \N__5635\
        );

    \I__745\ : CascadeBuf
    port map (
            O => \N__5638\,
            I => \N__5632\
        );

    \I__744\ : CascadeMux
    port map (
            O => \N__5635\,
            I => \N__5629\
        );

    \I__743\ : CascadeMux
    port map (
            O => \N__5632\,
            I => \N__5626\
        );

    \I__742\ : CascadeBuf
    port map (
            O => \N__5629\,
            I => \N__5623\
        );

    \I__741\ : CascadeBuf
    port map (
            O => \N__5626\,
            I => \N__5620\
        );

    \I__740\ : CascadeMux
    port map (
            O => \N__5623\,
            I => \N__5617\
        );

    \I__739\ : CascadeMux
    port map (
            O => \N__5620\,
            I => \N__5614\
        );

    \I__738\ : CascadeBuf
    port map (
            O => \N__5617\,
            I => \N__5611\
        );

    \I__737\ : CascadeBuf
    port map (
            O => \N__5614\,
            I => \N__5608\
        );

    \I__736\ : CascadeMux
    port map (
            O => \N__5611\,
            I => \N__5605\
        );

    \I__735\ : CascadeMux
    port map (
            O => \N__5608\,
            I => \N__5602\
        );

    \I__734\ : CascadeBuf
    port map (
            O => \N__5605\,
            I => \N__5599\
        );

    \I__733\ : CascadeBuf
    port map (
            O => \N__5602\,
            I => \N__5596\
        );

    \I__732\ : CascadeMux
    port map (
            O => \N__5599\,
            I => \N__5593\
        );

    \I__731\ : CascadeMux
    port map (
            O => \N__5596\,
            I => \N__5590\
        );

    \I__730\ : CascadeBuf
    port map (
            O => \N__5593\,
            I => \N__5587\
        );

    \I__729\ : CascadeBuf
    port map (
            O => \N__5590\,
            I => \N__5584\
        );

    \I__728\ : CascadeMux
    port map (
            O => \N__5587\,
            I => \N__5581\
        );

    \I__727\ : CascadeMux
    port map (
            O => \N__5584\,
            I => \N__5578\
        );

    \I__726\ : CascadeBuf
    port map (
            O => \N__5581\,
            I => \N__5575\
        );

    \I__725\ : CascadeBuf
    port map (
            O => \N__5578\,
            I => \N__5572\
        );

    \I__724\ : CascadeMux
    port map (
            O => \N__5575\,
            I => \N__5569\
        );

    \I__723\ : CascadeMux
    port map (
            O => \N__5572\,
            I => \N__5566\
        );

    \I__722\ : CascadeBuf
    port map (
            O => \N__5569\,
            I => \N__5563\
        );

    \I__721\ : CascadeBuf
    port map (
            O => \N__5566\,
            I => \N__5560\
        );

    \I__720\ : CascadeMux
    port map (
            O => \N__5563\,
            I => \N__5557\
        );

    \I__719\ : CascadeMux
    port map (
            O => \N__5560\,
            I => \N__5554\
        );

    \I__718\ : CascadeBuf
    port map (
            O => \N__5557\,
            I => \N__5551\
        );

    \I__717\ : CascadeBuf
    port map (
            O => \N__5554\,
            I => \N__5548\
        );

    \I__716\ : CascadeMux
    port map (
            O => \N__5551\,
            I => \N__5545\
        );

    \I__715\ : CascadeMux
    port map (
            O => \N__5548\,
            I => \N__5542\
        );

    \I__714\ : CascadeBuf
    port map (
            O => \N__5545\,
            I => \N__5539\
        );

    \I__713\ : InMux
    port map (
            O => \N__5542\,
            I => \N__5536\
        );

    \I__712\ : CascadeMux
    port map (
            O => \N__5539\,
            I => \N__5533\
        );

    \I__711\ : LocalMux
    port map (
            O => \N__5536\,
            I => \N__5530\
        );

    \I__710\ : InMux
    port map (
            O => \N__5533\,
            I => \N__5527\
        );

    \I__709\ : Span4Mux_v
    port map (
            O => \N__5530\,
            I => \N__5524\
        );

    \I__708\ : LocalMux
    port map (
            O => \N__5527\,
            I => \N__5521\
        );

    \I__707\ : Span4Mux_h
    port map (
            O => \N__5524\,
            I => \N__5518\
        );

    \I__706\ : Span4Mux_v
    port map (
            O => \N__5521\,
            I => \N__5515\
        );

    \I__705\ : Sp12to4
    port map (
            O => \N__5518\,
            I => \N__5512\
        );

    \I__704\ : Span4Mux_v
    port map (
            O => \N__5515\,
            I => \N__5509\
        );

    \I__703\ : Span12Mux_v
    port map (
            O => \N__5512\,
            I => \N__5506\
        );

    \I__702\ : Span4Mux_v
    port map (
            O => \N__5509\,
            I => \N__5503\
        );

    \I__701\ : Span12Mux_h
    port map (
            O => \N__5506\,
            I => \N__5498\
        );

    \I__700\ : Sp12to4
    port map (
            O => \N__5503\,
            I => \N__5498\
        );

    \I__699\ : Odrv12
    port map (
            O => \N__5498\,
            I => raddr_c_1
        );

    \I__698\ : CascadeMux
    port map (
            O => \N__5495\,
            I => \N__5492\
        );

    \I__697\ : CascadeBuf
    port map (
            O => \N__5492\,
            I => \N__5488\
        );

    \I__696\ : CascadeMux
    port map (
            O => \N__5491\,
            I => \N__5485\
        );

    \I__695\ : CascadeMux
    port map (
            O => \N__5488\,
            I => \N__5482\
        );

    \I__694\ : CascadeBuf
    port map (
            O => \N__5485\,
            I => \N__5479\
        );

    \I__693\ : CascadeBuf
    port map (
            O => \N__5482\,
            I => \N__5476\
        );

    \I__692\ : CascadeMux
    port map (
            O => \N__5479\,
            I => \N__5473\
        );

    \I__691\ : CascadeMux
    port map (
            O => \N__5476\,
            I => \N__5470\
        );

    \I__690\ : CascadeBuf
    port map (
            O => \N__5473\,
            I => \N__5467\
        );

    \I__689\ : CascadeBuf
    port map (
            O => \N__5470\,
            I => \N__5464\
        );

    \I__688\ : CascadeMux
    port map (
            O => \N__5467\,
            I => \N__5461\
        );

    \I__687\ : CascadeMux
    port map (
            O => \N__5464\,
            I => \N__5458\
        );

    \I__686\ : CascadeBuf
    port map (
            O => \N__5461\,
            I => \N__5455\
        );

    \I__685\ : CascadeBuf
    port map (
            O => \N__5458\,
            I => \N__5452\
        );

    \I__684\ : CascadeMux
    port map (
            O => \N__5455\,
            I => \N__5449\
        );

    \I__683\ : CascadeMux
    port map (
            O => \N__5452\,
            I => \N__5446\
        );

    \I__682\ : CascadeBuf
    port map (
            O => \N__5449\,
            I => \N__5443\
        );

    \I__681\ : CascadeBuf
    port map (
            O => \N__5446\,
            I => \N__5440\
        );

    \I__680\ : CascadeMux
    port map (
            O => \N__5443\,
            I => \N__5437\
        );

    \I__679\ : CascadeMux
    port map (
            O => \N__5440\,
            I => \N__5434\
        );

    \I__678\ : CascadeBuf
    port map (
            O => \N__5437\,
            I => \N__5431\
        );

    \I__677\ : CascadeBuf
    port map (
            O => \N__5434\,
            I => \N__5428\
        );

    \I__676\ : CascadeMux
    port map (
            O => \N__5431\,
            I => \N__5425\
        );

    \I__675\ : CascadeMux
    port map (
            O => \N__5428\,
            I => \N__5422\
        );

    \I__674\ : CascadeBuf
    port map (
            O => \N__5425\,
            I => \N__5419\
        );

    \I__673\ : CascadeBuf
    port map (
            O => \N__5422\,
            I => \N__5416\
        );

    \I__672\ : CascadeMux
    port map (
            O => \N__5419\,
            I => \N__5413\
        );

    \I__671\ : CascadeMux
    port map (
            O => \N__5416\,
            I => \N__5410\
        );

    \I__670\ : CascadeBuf
    port map (
            O => \N__5413\,
            I => \N__5407\
        );

    \I__669\ : CascadeBuf
    port map (
            O => \N__5410\,
            I => \N__5404\
        );

    \I__668\ : CascadeMux
    port map (
            O => \N__5407\,
            I => \N__5401\
        );

    \I__667\ : CascadeMux
    port map (
            O => \N__5404\,
            I => \N__5398\
        );

    \I__666\ : CascadeBuf
    port map (
            O => \N__5401\,
            I => \N__5395\
        );

    \I__665\ : CascadeBuf
    port map (
            O => \N__5398\,
            I => \N__5392\
        );

    \I__664\ : CascadeMux
    port map (
            O => \N__5395\,
            I => \N__5389\
        );

    \I__663\ : CascadeMux
    port map (
            O => \N__5392\,
            I => \N__5386\
        );

    \I__662\ : CascadeBuf
    port map (
            O => \N__5389\,
            I => \N__5383\
        );

    \I__661\ : CascadeBuf
    port map (
            O => \N__5386\,
            I => \N__5380\
        );

    \I__660\ : CascadeMux
    port map (
            O => \N__5383\,
            I => \N__5377\
        );

    \I__659\ : CascadeMux
    port map (
            O => \N__5380\,
            I => \N__5374\
        );

    \I__658\ : CascadeBuf
    port map (
            O => \N__5377\,
            I => \N__5371\
        );

    \I__657\ : CascadeBuf
    port map (
            O => \N__5374\,
            I => \N__5368\
        );

    \I__656\ : CascadeMux
    port map (
            O => \N__5371\,
            I => \N__5365\
        );

    \I__655\ : CascadeMux
    port map (
            O => \N__5368\,
            I => \N__5362\
        );

    \I__654\ : CascadeBuf
    port map (
            O => \N__5365\,
            I => \N__5359\
        );

    \I__653\ : CascadeBuf
    port map (
            O => \N__5362\,
            I => \N__5356\
        );

    \I__652\ : CascadeMux
    port map (
            O => \N__5359\,
            I => \N__5353\
        );

    \I__651\ : CascadeMux
    port map (
            O => \N__5356\,
            I => \N__5350\
        );

    \I__650\ : CascadeBuf
    port map (
            O => \N__5353\,
            I => \N__5347\
        );

    \I__649\ : CascadeBuf
    port map (
            O => \N__5350\,
            I => \N__5344\
        );

    \I__648\ : CascadeMux
    port map (
            O => \N__5347\,
            I => \N__5341\
        );

    \I__647\ : CascadeMux
    port map (
            O => \N__5344\,
            I => \N__5338\
        );

    \I__646\ : CascadeBuf
    port map (
            O => \N__5341\,
            I => \N__5335\
        );

    \I__645\ : CascadeBuf
    port map (
            O => \N__5338\,
            I => \N__5332\
        );

    \I__644\ : CascadeMux
    port map (
            O => \N__5335\,
            I => \N__5329\
        );

    \I__643\ : CascadeMux
    port map (
            O => \N__5332\,
            I => \N__5326\
        );

    \I__642\ : CascadeBuf
    port map (
            O => \N__5329\,
            I => \N__5323\
        );

    \I__641\ : CascadeBuf
    port map (
            O => \N__5326\,
            I => \N__5320\
        );

    \I__640\ : CascadeMux
    port map (
            O => \N__5323\,
            I => \N__5317\
        );

    \I__639\ : CascadeMux
    port map (
            O => \N__5320\,
            I => \N__5314\
        );

    \I__638\ : CascadeBuf
    port map (
            O => \N__5317\,
            I => \N__5311\
        );

    \I__637\ : InMux
    port map (
            O => \N__5314\,
            I => \N__5308\
        );

    \I__636\ : CascadeMux
    port map (
            O => \N__5311\,
            I => \N__5305\
        );

    \I__635\ : LocalMux
    port map (
            O => \N__5308\,
            I => \N__5302\
        );

    \I__634\ : InMux
    port map (
            O => \N__5305\,
            I => \N__5299\
        );

    \I__633\ : Span4Mux_h
    port map (
            O => \N__5302\,
            I => \N__5296\
        );

    \I__632\ : LocalMux
    port map (
            O => \N__5299\,
            I => \N__5293\
        );

    \I__631\ : Sp12to4
    port map (
            O => \N__5296\,
            I => \N__5290\
        );

    \I__630\ : Span4Mux_s3_v
    port map (
            O => \N__5293\,
            I => \N__5287\
        );

    \I__629\ : Span12Mux_s7_v
    port map (
            O => \N__5290\,
            I => \N__5284\
        );

    \I__628\ : Span4Mux_h
    port map (
            O => \N__5287\,
            I => \N__5281\
        );

    \I__627\ : Span12Mux_h
    port map (
            O => \N__5284\,
            I => \N__5278\
        );

    \I__626\ : Span4Mux_v
    port map (
            O => \N__5281\,
            I => \N__5275\
        );

    \I__625\ : Odrv12
    port map (
            O => \N__5278\,
            I => raddr_c_6
        );

    \I__624\ : Odrv4
    port map (
            O => \N__5275\,
            I => raddr_c_6
        );

    \I__623\ : CascadeMux
    port map (
            O => \N__5270\,
            I => \N__5267\
        );

    \I__622\ : CascadeBuf
    port map (
            O => \N__5267\,
            I => \N__5264\
        );

    \I__621\ : CascadeMux
    port map (
            O => \N__5264\,
            I => \N__5261\
        );

    \I__620\ : CascadeBuf
    port map (
            O => \N__5261\,
            I => \N__5258\
        );

    \I__619\ : CascadeMux
    port map (
            O => \N__5258\,
            I => \N__5254\
        );

    \I__618\ : CascadeMux
    port map (
            O => \N__5257\,
            I => \N__5251\
        );

    \I__617\ : CascadeBuf
    port map (
            O => \N__5254\,
            I => \N__5248\
        );

    \I__616\ : CascadeBuf
    port map (
            O => \N__5251\,
            I => \N__5245\
        );

    \I__615\ : CascadeMux
    port map (
            O => \N__5248\,
            I => \N__5242\
        );

    \I__614\ : CascadeMux
    port map (
            O => \N__5245\,
            I => \N__5239\
        );

    \I__613\ : CascadeBuf
    port map (
            O => \N__5242\,
            I => \N__5236\
        );

    \I__612\ : CascadeBuf
    port map (
            O => \N__5239\,
            I => \N__5233\
        );

    \I__611\ : CascadeMux
    port map (
            O => \N__5236\,
            I => \N__5230\
        );

    \I__610\ : CascadeMux
    port map (
            O => \N__5233\,
            I => \N__5227\
        );

    \I__609\ : CascadeBuf
    port map (
            O => \N__5230\,
            I => \N__5224\
        );

    \I__608\ : CascadeBuf
    port map (
            O => \N__5227\,
            I => \N__5221\
        );

    \I__607\ : CascadeMux
    port map (
            O => \N__5224\,
            I => \N__5218\
        );

    \I__606\ : CascadeMux
    port map (
            O => \N__5221\,
            I => \N__5215\
        );

    \I__605\ : CascadeBuf
    port map (
            O => \N__5218\,
            I => \N__5212\
        );

    \I__604\ : CascadeBuf
    port map (
            O => \N__5215\,
            I => \N__5209\
        );

    \I__603\ : CascadeMux
    port map (
            O => \N__5212\,
            I => \N__5206\
        );

    \I__602\ : CascadeMux
    port map (
            O => \N__5209\,
            I => \N__5203\
        );

    \I__601\ : CascadeBuf
    port map (
            O => \N__5206\,
            I => \N__5200\
        );

    \I__600\ : CascadeBuf
    port map (
            O => \N__5203\,
            I => \N__5197\
        );

    \I__599\ : CascadeMux
    port map (
            O => \N__5200\,
            I => \N__5194\
        );

    \I__598\ : CascadeMux
    port map (
            O => \N__5197\,
            I => \N__5191\
        );

    \I__597\ : CascadeBuf
    port map (
            O => \N__5194\,
            I => \N__5188\
        );

    \I__596\ : CascadeBuf
    port map (
            O => \N__5191\,
            I => \N__5185\
        );

    \I__595\ : CascadeMux
    port map (
            O => \N__5188\,
            I => \N__5182\
        );

    \I__594\ : CascadeMux
    port map (
            O => \N__5185\,
            I => \N__5179\
        );

    \I__593\ : CascadeBuf
    port map (
            O => \N__5182\,
            I => \N__5176\
        );

    \I__592\ : CascadeBuf
    port map (
            O => \N__5179\,
            I => \N__5173\
        );

    \I__591\ : CascadeMux
    port map (
            O => \N__5176\,
            I => \N__5170\
        );

    \I__590\ : CascadeMux
    port map (
            O => \N__5173\,
            I => \N__5167\
        );

    \I__589\ : CascadeBuf
    port map (
            O => \N__5170\,
            I => \N__5164\
        );

    \I__588\ : CascadeBuf
    port map (
            O => \N__5167\,
            I => \N__5161\
        );

    \I__587\ : CascadeMux
    port map (
            O => \N__5164\,
            I => \N__5158\
        );

    \I__586\ : CascadeMux
    port map (
            O => \N__5161\,
            I => \N__5155\
        );

    \I__585\ : CascadeBuf
    port map (
            O => \N__5158\,
            I => \N__5152\
        );

    \I__584\ : CascadeBuf
    port map (
            O => \N__5155\,
            I => \N__5149\
        );

    \I__583\ : CascadeMux
    port map (
            O => \N__5152\,
            I => \N__5146\
        );

    \I__582\ : CascadeMux
    port map (
            O => \N__5149\,
            I => \N__5143\
        );

    \I__581\ : CascadeBuf
    port map (
            O => \N__5146\,
            I => \N__5140\
        );

    \I__580\ : CascadeBuf
    port map (
            O => \N__5143\,
            I => \N__5137\
        );

    \I__579\ : CascadeMux
    port map (
            O => \N__5140\,
            I => \N__5134\
        );

    \I__578\ : CascadeMux
    port map (
            O => \N__5137\,
            I => \N__5131\
        );

    \I__577\ : CascadeBuf
    port map (
            O => \N__5134\,
            I => \N__5128\
        );

    \I__576\ : CascadeBuf
    port map (
            O => \N__5131\,
            I => \N__5125\
        );

    \I__575\ : CascadeMux
    port map (
            O => \N__5128\,
            I => \N__5122\
        );

    \I__574\ : CascadeMux
    port map (
            O => \N__5125\,
            I => \N__5119\
        );

    \I__573\ : CascadeBuf
    port map (
            O => \N__5122\,
            I => \N__5116\
        );

    \I__572\ : CascadeBuf
    port map (
            O => \N__5119\,
            I => \N__5113\
        );

    \I__571\ : CascadeMux
    port map (
            O => \N__5116\,
            I => \N__5110\
        );

    \I__570\ : CascadeMux
    port map (
            O => \N__5113\,
            I => \N__5107\
        );

    \I__569\ : CascadeBuf
    port map (
            O => \N__5110\,
            I => \N__5104\
        );

    \I__568\ : CascadeBuf
    port map (
            O => \N__5107\,
            I => \N__5101\
        );

    \I__567\ : CascadeMux
    port map (
            O => \N__5104\,
            I => \N__5098\
        );

    \I__566\ : CascadeMux
    port map (
            O => \N__5101\,
            I => \N__5095\
        );

    \I__565\ : InMux
    port map (
            O => \N__5098\,
            I => \N__5092\
        );

    \I__564\ : CascadeBuf
    port map (
            O => \N__5095\,
            I => \N__5089\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__5092\,
            I => \N__5086\
        );

    \I__562\ : CascadeMux
    port map (
            O => \N__5089\,
            I => \N__5083\
        );

    \I__561\ : Span4Mux_h
    port map (
            O => \N__5086\,
            I => \N__5080\
        );

    \I__560\ : CascadeBuf
    port map (
            O => \N__5083\,
            I => \N__5077\
        );

    \I__559\ : Span4Mux_h
    port map (
            O => \N__5080\,
            I => \N__5074\
        );

    \I__558\ : CascadeMux
    port map (
            O => \N__5077\,
            I => \N__5071\
        );

    \I__557\ : Span4Mux_h
    port map (
            O => \N__5074\,
            I => \N__5068\
        );

    \I__556\ : InMux
    port map (
            O => \N__5071\,
            I => \N__5065\
        );

    \I__555\ : Span4Mux_h
    port map (
            O => \N__5068\,
            I => \N__5060\
        );

    \I__554\ : LocalMux
    port map (
            O => \N__5065\,
            I => \N__5060\
        );

    \I__553\ : Span4Mux_h
    port map (
            O => \N__5060\,
            I => \N__5057\
        );

    \I__552\ : IoSpan4Mux
    port map (
            O => \N__5057\,
            I => \N__5054\
        );

    \I__551\ : Odrv4
    port map (
            O => \N__5054\,
            I => waddr_c_2
        );

    \I__550\ : InMux
    port map (
            O => \N__5051\,
            I => \N__5047\
        );

    \I__549\ : InMux
    port map (
            O => \N__5050\,
            I => \N__5044\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__5047\,
            I => \N__5041\
        );

    \I__547\ : LocalMux
    port map (
            O => \N__5044\,
            I => \N__5037\
        );

    \I__546\ : Span4Mux_s2_v
    port map (
            O => \N__5041\,
            I => \N__5033\
        );

    \I__545\ : InMux
    port map (
            O => \N__5040\,
            I => \N__5030\
        );

    \I__544\ : Span4Mux_h
    port map (
            O => \N__5037\,
            I => \N__5027\
        );

    \I__543\ : InMux
    port map (
            O => \N__5036\,
            I => \N__5024\
        );

    \I__542\ : Span4Mux_v
    port map (
            O => \N__5033\,
            I => \N__5019\
        );

    \I__541\ : LocalMux
    port map (
            O => \N__5030\,
            I => \N__5019\
        );

    \I__540\ : Span4Mux_v
    port map (
            O => \N__5027\,
            I => \N__5015\
        );

    \I__539\ : LocalMux
    port map (
            O => \N__5024\,
            I => \N__5012\
        );

    \I__538\ : Span4Mux_v
    port map (
            O => \N__5019\,
            I => \N__5008\
        );

    \I__537\ : InMux
    port map (
            O => \N__5018\,
            I => \N__5005\
        );

    \I__536\ : Span4Mux_v
    port map (
            O => \N__5015\,
            I => \N__5000\
        );

    \I__535\ : Span4Mux_h
    port map (
            O => \N__5012\,
            I => \N__5000\
        );

    \I__534\ : InMux
    port map (
            O => \N__5011\,
            I => \N__4997\
        );

    \I__533\ : Span4Mux_v
    port map (
            O => \N__5008\,
            I => \N__4992\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__5005\,
            I => \N__4992\
        );

    \I__531\ : Span4Mux_v
    port map (
            O => \N__5000\,
            I => \N__4988\
        );

    \I__530\ : LocalMux
    port map (
            O => \N__4997\,
            I => \N__4985\
        );

    \I__529\ : Span4Mux_v
    port map (
            O => \N__4992\,
            I => \N__4981\
        );

    \I__528\ : InMux
    port map (
            O => \N__4991\,
            I => \N__4978\
        );

    \I__527\ : Span4Mux_v
    port map (
            O => \N__4988\,
            I => \N__4973\
        );

    \I__526\ : Span4Mux_h
    port map (
            O => \N__4985\,
            I => \N__4973\
        );

    \I__525\ : InMux
    port map (
            O => \N__4984\,
            I => \N__4970\
        );

    \I__524\ : Span4Mux_v
    port map (
            O => \N__4981\,
            I => \N__4965\
        );

    \I__523\ : LocalMux
    port map (
            O => \N__4978\,
            I => \N__4965\
        );

    \I__522\ : Span4Mux_v
    port map (
            O => \N__4973\,
            I => \N__4962\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__4970\,
            I => \N__4959\
        );

    \I__520\ : Span4Mux_v
    port map (
            O => \N__4965\,
            I => \N__4956\
        );

    \I__519\ : Span4Mux_v
    port map (
            O => \N__4962\,
            I => \N__4951\
        );

    \I__518\ : Span4Mux_h
    port map (
            O => \N__4959\,
            I => \N__4951\
        );

    \I__517\ : Sp12to4
    port map (
            O => \N__4956\,
            I => \N__4948\
        );

    \I__516\ : Span4Mux_v
    port map (
            O => \N__4951\,
            I => \N__4945\
        );

    \I__515\ : Span12Mux_h
    port map (
            O => \N__4948\,
            I => \N__4942\
        );

    \I__514\ : Span4Mux_h
    port map (
            O => \N__4945\,
            I => \N__4939\
        );

    \I__513\ : Odrv12
    port map (
            O => \N__4942\,
            I => din_c_0
        );

    \I__512\ : Odrv4
    port map (
            O => \N__4939\,
            I => din_c_0
        );

    \I__511\ : ClkMux
    port map (
            O => \N__4934\,
            I => \N__4829\
        );

    \I__510\ : ClkMux
    port map (
            O => \N__4933\,
            I => \N__4829\
        );

    \I__509\ : ClkMux
    port map (
            O => \N__4932\,
            I => \N__4829\
        );

    \I__508\ : ClkMux
    port map (
            O => \N__4931\,
            I => \N__4829\
        );

    \I__507\ : ClkMux
    port map (
            O => \N__4930\,
            I => \N__4829\
        );

    \I__506\ : ClkMux
    port map (
            O => \N__4929\,
            I => \N__4829\
        );

    \I__505\ : ClkMux
    port map (
            O => \N__4928\,
            I => \N__4829\
        );

    \I__504\ : ClkMux
    port map (
            O => \N__4927\,
            I => \N__4829\
        );

    \I__503\ : ClkMux
    port map (
            O => \N__4926\,
            I => \N__4829\
        );

    \I__502\ : ClkMux
    port map (
            O => \N__4925\,
            I => \N__4829\
        );

    \I__501\ : ClkMux
    port map (
            O => \N__4924\,
            I => \N__4829\
        );

    \I__500\ : ClkMux
    port map (
            O => \N__4923\,
            I => \N__4829\
        );

    \I__499\ : ClkMux
    port map (
            O => \N__4922\,
            I => \N__4829\
        );

    \I__498\ : ClkMux
    port map (
            O => \N__4921\,
            I => \N__4829\
        );

    \I__497\ : ClkMux
    port map (
            O => \N__4920\,
            I => \N__4829\
        );

    \I__496\ : ClkMux
    port map (
            O => \N__4919\,
            I => \N__4829\
        );

    \I__495\ : ClkMux
    port map (
            O => \N__4918\,
            I => \N__4829\
        );

    \I__494\ : ClkMux
    port map (
            O => \N__4917\,
            I => \N__4829\
        );

    \I__493\ : ClkMux
    port map (
            O => \N__4916\,
            I => \N__4829\
        );

    \I__492\ : ClkMux
    port map (
            O => \N__4915\,
            I => \N__4829\
        );

    \I__491\ : ClkMux
    port map (
            O => \N__4914\,
            I => \N__4829\
        );

    \I__490\ : ClkMux
    port map (
            O => \N__4913\,
            I => \N__4829\
        );

    \I__489\ : ClkMux
    port map (
            O => \N__4912\,
            I => \N__4829\
        );

    \I__488\ : ClkMux
    port map (
            O => \N__4911\,
            I => \N__4829\
        );

    \I__487\ : ClkMux
    port map (
            O => \N__4910\,
            I => \N__4829\
        );

    \I__486\ : ClkMux
    port map (
            O => \N__4909\,
            I => \N__4829\
        );

    \I__485\ : ClkMux
    port map (
            O => \N__4908\,
            I => \N__4829\
        );

    \I__484\ : ClkMux
    port map (
            O => \N__4907\,
            I => \N__4829\
        );

    \I__483\ : ClkMux
    port map (
            O => \N__4906\,
            I => \N__4829\
        );

    \I__482\ : ClkMux
    port map (
            O => \N__4905\,
            I => \N__4829\
        );

    \I__481\ : ClkMux
    port map (
            O => \N__4904\,
            I => \N__4829\
        );

    \I__480\ : ClkMux
    port map (
            O => \N__4903\,
            I => \N__4829\
        );

    \I__479\ : ClkMux
    port map (
            O => \N__4902\,
            I => \N__4829\
        );

    \I__478\ : ClkMux
    port map (
            O => \N__4901\,
            I => \N__4829\
        );

    \I__477\ : ClkMux
    port map (
            O => \N__4900\,
            I => \N__4829\
        );

    \I__476\ : GlobalMux
    port map (
            O => \N__4829\,
            I => \N__4826\
        );

    \I__475\ : gio2CtrlBuf
    port map (
            O => \N__4826\,
            I => rclk_c_g
        );

    \I__474\ : CascadeMux
    port map (
            O => \N__4823\,
            I => \N__4820\
        );

    \I__473\ : CascadeBuf
    port map (
            O => \N__4820\,
            I => \N__4817\
        );

    \I__472\ : CascadeMux
    port map (
            O => \N__4817\,
            I => \N__4814\
        );

    \I__471\ : CascadeBuf
    port map (
            O => \N__4814\,
            I => \N__4811\
        );

    \I__470\ : CascadeMux
    port map (
            O => \N__4811\,
            I => \N__4807\
        );

    \I__469\ : CascadeMux
    port map (
            O => \N__4810\,
            I => \N__4804\
        );

    \I__468\ : CascadeBuf
    port map (
            O => \N__4807\,
            I => \N__4801\
        );

    \I__467\ : CascadeBuf
    port map (
            O => \N__4804\,
            I => \N__4798\
        );

    \I__466\ : CascadeMux
    port map (
            O => \N__4801\,
            I => \N__4795\
        );

    \I__465\ : CascadeMux
    port map (
            O => \N__4798\,
            I => \N__4792\
        );

    \I__464\ : CascadeBuf
    port map (
            O => \N__4795\,
            I => \N__4789\
        );

    \I__463\ : CascadeBuf
    port map (
            O => \N__4792\,
            I => \N__4786\
        );

    \I__462\ : CascadeMux
    port map (
            O => \N__4789\,
            I => \N__4783\
        );

    \I__461\ : CascadeMux
    port map (
            O => \N__4786\,
            I => \N__4780\
        );

    \I__460\ : CascadeBuf
    port map (
            O => \N__4783\,
            I => \N__4777\
        );

    \I__459\ : CascadeBuf
    port map (
            O => \N__4780\,
            I => \N__4774\
        );

    \I__458\ : CascadeMux
    port map (
            O => \N__4777\,
            I => \N__4771\
        );

    \I__457\ : CascadeMux
    port map (
            O => \N__4774\,
            I => \N__4768\
        );

    \I__456\ : CascadeBuf
    port map (
            O => \N__4771\,
            I => \N__4765\
        );

    \I__455\ : CascadeBuf
    port map (
            O => \N__4768\,
            I => \N__4762\
        );

    \I__454\ : CascadeMux
    port map (
            O => \N__4765\,
            I => \N__4759\
        );

    \I__453\ : CascadeMux
    port map (
            O => \N__4762\,
            I => \N__4756\
        );

    \I__452\ : CascadeBuf
    port map (
            O => \N__4759\,
            I => \N__4753\
        );

    \I__451\ : CascadeBuf
    port map (
            O => \N__4756\,
            I => \N__4750\
        );

    \I__450\ : CascadeMux
    port map (
            O => \N__4753\,
            I => \N__4747\
        );

    \I__449\ : CascadeMux
    port map (
            O => \N__4750\,
            I => \N__4744\
        );

    \I__448\ : CascadeBuf
    port map (
            O => \N__4747\,
            I => \N__4741\
        );

    \I__447\ : CascadeBuf
    port map (
            O => \N__4744\,
            I => \N__4738\
        );

    \I__446\ : CascadeMux
    port map (
            O => \N__4741\,
            I => \N__4735\
        );

    \I__445\ : CascadeMux
    port map (
            O => \N__4738\,
            I => \N__4732\
        );

    \I__444\ : CascadeBuf
    port map (
            O => \N__4735\,
            I => \N__4729\
        );

    \I__443\ : CascadeBuf
    port map (
            O => \N__4732\,
            I => \N__4726\
        );

    \I__442\ : CascadeMux
    port map (
            O => \N__4729\,
            I => \N__4723\
        );

    \I__441\ : CascadeMux
    port map (
            O => \N__4726\,
            I => \N__4720\
        );

    \I__440\ : CascadeBuf
    port map (
            O => \N__4723\,
            I => \N__4717\
        );

    \I__439\ : CascadeBuf
    port map (
            O => \N__4720\,
            I => \N__4714\
        );

    \I__438\ : CascadeMux
    port map (
            O => \N__4717\,
            I => \N__4711\
        );

    \I__437\ : CascadeMux
    port map (
            O => \N__4714\,
            I => \N__4708\
        );

    \I__436\ : CascadeBuf
    port map (
            O => \N__4711\,
            I => \N__4705\
        );

    \I__435\ : CascadeBuf
    port map (
            O => \N__4708\,
            I => \N__4702\
        );

    \I__434\ : CascadeMux
    port map (
            O => \N__4705\,
            I => \N__4699\
        );

    \I__433\ : CascadeMux
    port map (
            O => \N__4702\,
            I => \N__4696\
        );

    \I__432\ : CascadeBuf
    port map (
            O => \N__4699\,
            I => \N__4693\
        );

    \I__431\ : CascadeBuf
    port map (
            O => \N__4696\,
            I => \N__4690\
        );

    \I__430\ : CascadeMux
    port map (
            O => \N__4693\,
            I => \N__4687\
        );

    \I__429\ : CascadeMux
    port map (
            O => \N__4690\,
            I => \N__4684\
        );

    \I__428\ : CascadeBuf
    port map (
            O => \N__4687\,
            I => \N__4681\
        );

    \I__427\ : CascadeBuf
    port map (
            O => \N__4684\,
            I => \N__4678\
        );

    \I__426\ : CascadeMux
    port map (
            O => \N__4681\,
            I => \N__4675\
        );

    \I__425\ : CascadeMux
    port map (
            O => \N__4678\,
            I => \N__4672\
        );

    \I__424\ : CascadeBuf
    port map (
            O => \N__4675\,
            I => \N__4669\
        );

    \I__423\ : CascadeBuf
    port map (
            O => \N__4672\,
            I => \N__4666\
        );

    \I__422\ : CascadeMux
    port map (
            O => \N__4669\,
            I => \N__4663\
        );

    \I__421\ : CascadeMux
    port map (
            O => \N__4666\,
            I => \N__4660\
        );

    \I__420\ : CascadeBuf
    port map (
            O => \N__4663\,
            I => \N__4657\
        );

    \I__419\ : CascadeBuf
    port map (
            O => \N__4660\,
            I => \N__4654\
        );

    \I__418\ : CascadeMux
    port map (
            O => \N__4657\,
            I => \N__4651\
        );

    \I__417\ : CascadeMux
    port map (
            O => \N__4654\,
            I => \N__4648\
        );

    \I__416\ : InMux
    port map (
            O => \N__4651\,
            I => \N__4645\
        );

    \I__415\ : CascadeBuf
    port map (
            O => \N__4648\,
            I => \N__4642\
        );

    \I__414\ : LocalMux
    port map (
            O => \N__4645\,
            I => \N__4639\
        );

    \I__413\ : CascadeMux
    port map (
            O => \N__4642\,
            I => \N__4636\
        );

    \I__412\ : Span4Mux_s2_v
    port map (
            O => \N__4639\,
            I => \N__4633\
        );

    \I__411\ : CascadeBuf
    port map (
            O => \N__4636\,
            I => \N__4630\
        );

    \I__410\ : Span4Mux_h
    port map (
            O => \N__4633\,
            I => \N__4627\
        );

    \I__409\ : CascadeMux
    port map (
            O => \N__4630\,
            I => \N__4624\
        );

    \I__408\ : Span4Mux_v
    port map (
            O => \N__4627\,
            I => \N__4621\
        );

    \I__407\ : InMux
    port map (
            O => \N__4624\,
            I => \N__4618\
        );

    \I__406\ : Span4Mux_v
    port map (
            O => \N__4621\,
            I => \N__4615\
        );

    \I__405\ : LocalMux
    port map (
            O => \N__4618\,
            I => \N__4612\
        );

    \I__404\ : Sp12to4
    port map (
            O => \N__4615\,
            I => \N__4609\
        );

    \I__403\ : Sp12to4
    port map (
            O => \N__4612\,
            I => \N__4606\
        );

    \I__402\ : Span12Mux_h
    port map (
            O => \N__4609\,
            I => \N__4601\
        );

    \I__401\ : Span12Mux_s10_v
    port map (
            O => \N__4606\,
            I => \N__4601\
        );

    \I__400\ : Odrv12
    port map (
            O => \N__4601\,
            I => raddr_c_3
        );

    \I__399\ : CascadeMux
    port map (
            O => \N__4598\,
            I => \N__4595\
        );

    \I__398\ : CascadeBuf
    port map (
            O => \N__4595\,
            I => \N__4592\
        );

    \I__397\ : CascadeMux
    port map (
            O => \N__4592\,
            I => \N__4589\
        );

    \I__396\ : CascadeBuf
    port map (
            O => \N__4589\,
            I => \N__4586\
        );

    \I__395\ : CascadeMux
    port map (
            O => \N__4586\,
            I => \N__4582\
        );

    \I__394\ : CascadeMux
    port map (
            O => \N__4585\,
            I => \N__4579\
        );

    \I__393\ : CascadeBuf
    port map (
            O => \N__4582\,
            I => \N__4576\
        );

    \I__392\ : CascadeBuf
    port map (
            O => \N__4579\,
            I => \N__4573\
        );

    \I__391\ : CascadeMux
    port map (
            O => \N__4576\,
            I => \N__4570\
        );

    \I__390\ : CascadeMux
    port map (
            O => \N__4573\,
            I => \N__4567\
        );

    \I__389\ : CascadeBuf
    port map (
            O => \N__4570\,
            I => \N__4564\
        );

    \I__388\ : CascadeBuf
    port map (
            O => \N__4567\,
            I => \N__4561\
        );

    \I__387\ : CascadeMux
    port map (
            O => \N__4564\,
            I => \N__4558\
        );

    \I__386\ : CascadeMux
    port map (
            O => \N__4561\,
            I => \N__4555\
        );

    \I__385\ : CascadeBuf
    port map (
            O => \N__4558\,
            I => \N__4552\
        );

    \I__384\ : CascadeBuf
    port map (
            O => \N__4555\,
            I => \N__4549\
        );

    \I__383\ : CascadeMux
    port map (
            O => \N__4552\,
            I => \N__4546\
        );

    \I__382\ : CascadeMux
    port map (
            O => \N__4549\,
            I => \N__4543\
        );

    \I__381\ : CascadeBuf
    port map (
            O => \N__4546\,
            I => \N__4540\
        );

    \I__380\ : CascadeBuf
    port map (
            O => \N__4543\,
            I => \N__4537\
        );

    \I__379\ : CascadeMux
    port map (
            O => \N__4540\,
            I => \N__4534\
        );

    \I__378\ : CascadeMux
    port map (
            O => \N__4537\,
            I => \N__4531\
        );

    \I__377\ : CascadeBuf
    port map (
            O => \N__4534\,
            I => \N__4528\
        );

    \I__376\ : CascadeBuf
    port map (
            O => \N__4531\,
            I => \N__4525\
        );

    \I__375\ : CascadeMux
    port map (
            O => \N__4528\,
            I => \N__4522\
        );

    \I__374\ : CascadeMux
    port map (
            O => \N__4525\,
            I => \N__4519\
        );

    \I__373\ : CascadeBuf
    port map (
            O => \N__4522\,
            I => \N__4516\
        );

    \I__372\ : CascadeBuf
    port map (
            O => \N__4519\,
            I => \N__4513\
        );

    \I__371\ : CascadeMux
    port map (
            O => \N__4516\,
            I => \N__4510\
        );

    \I__370\ : CascadeMux
    port map (
            O => \N__4513\,
            I => \N__4507\
        );

    \I__369\ : CascadeBuf
    port map (
            O => \N__4510\,
            I => \N__4504\
        );

    \I__368\ : CascadeBuf
    port map (
            O => \N__4507\,
            I => \N__4501\
        );

    \I__367\ : CascadeMux
    port map (
            O => \N__4504\,
            I => \N__4498\
        );

    \I__366\ : CascadeMux
    port map (
            O => \N__4501\,
            I => \N__4495\
        );

    \I__365\ : CascadeBuf
    port map (
            O => \N__4498\,
            I => \N__4492\
        );

    \I__364\ : CascadeBuf
    port map (
            O => \N__4495\,
            I => \N__4489\
        );

    \I__363\ : CascadeMux
    port map (
            O => \N__4492\,
            I => \N__4486\
        );

    \I__362\ : CascadeMux
    port map (
            O => \N__4489\,
            I => \N__4483\
        );

    \I__361\ : CascadeBuf
    port map (
            O => \N__4486\,
            I => \N__4480\
        );

    \I__360\ : CascadeBuf
    port map (
            O => \N__4483\,
            I => \N__4477\
        );

    \I__359\ : CascadeMux
    port map (
            O => \N__4480\,
            I => \N__4474\
        );

    \I__358\ : CascadeMux
    port map (
            O => \N__4477\,
            I => \N__4471\
        );

    \I__357\ : CascadeBuf
    port map (
            O => \N__4474\,
            I => \N__4468\
        );

    \I__356\ : CascadeBuf
    port map (
            O => \N__4471\,
            I => \N__4465\
        );

    \I__355\ : CascadeMux
    port map (
            O => \N__4468\,
            I => \N__4462\
        );

    \I__354\ : CascadeMux
    port map (
            O => \N__4465\,
            I => \N__4459\
        );

    \I__353\ : CascadeBuf
    port map (
            O => \N__4462\,
            I => \N__4456\
        );

    \I__352\ : CascadeBuf
    port map (
            O => \N__4459\,
            I => \N__4453\
        );

    \I__351\ : CascadeMux
    port map (
            O => \N__4456\,
            I => \N__4450\
        );

    \I__350\ : CascadeMux
    port map (
            O => \N__4453\,
            I => \N__4447\
        );

    \I__349\ : CascadeBuf
    port map (
            O => \N__4450\,
            I => \N__4444\
        );

    \I__348\ : CascadeBuf
    port map (
            O => \N__4447\,
            I => \N__4441\
        );

    \I__347\ : CascadeMux
    port map (
            O => \N__4444\,
            I => \N__4438\
        );

    \I__346\ : CascadeMux
    port map (
            O => \N__4441\,
            I => \N__4435\
        );

    \I__345\ : CascadeBuf
    port map (
            O => \N__4438\,
            I => \N__4432\
        );

    \I__344\ : CascadeBuf
    port map (
            O => \N__4435\,
            I => \N__4429\
        );

    \I__343\ : CascadeMux
    port map (
            O => \N__4432\,
            I => \N__4426\
        );

    \I__342\ : CascadeMux
    port map (
            O => \N__4429\,
            I => \N__4423\
        );

    \I__341\ : InMux
    port map (
            O => \N__4426\,
            I => \N__4420\
        );

    \I__340\ : CascadeBuf
    port map (
            O => \N__4423\,
            I => \N__4417\
        );

    \I__339\ : LocalMux
    port map (
            O => \N__4420\,
            I => \N__4414\
        );

    \I__338\ : CascadeMux
    port map (
            O => \N__4417\,
            I => \N__4411\
        );

    \I__337\ : IoSpan4Mux
    port map (
            O => \N__4414\,
            I => \N__4408\
        );

    \I__336\ : CascadeBuf
    port map (
            O => \N__4411\,
            I => \N__4405\
        );

    \I__335\ : IoSpan4Mux
    port map (
            O => \N__4408\,
            I => \N__4402\
        );

    \I__334\ : CascadeMux
    port map (
            O => \N__4405\,
            I => \N__4399\
        );

    \I__333\ : IoSpan4Mux
    port map (
            O => \N__4402\,
            I => \N__4396\
        );

    \I__332\ : InMux
    port map (
            O => \N__4399\,
            I => \N__4393\
        );

    \I__331\ : IoSpan4Mux
    port map (
            O => \N__4396\,
            I => \N__4390\
        );

    \I__330\ : LocalMux
    port map (
            O => \N__4393\,
            I => \N__4387\
        );

    \I__329\ : IoSpan4Mux
    port map (
            O => \N__4390\,
            I => \N__4382\
        );

    \I__328\ : IoSpan4Mux
    port map (
            O => \N__4387\,
            I => \N__4382\
        );

    \I__327\ : IoSpan4Mux
    port map (
            O => \N__4382\,
            I => \N__4379\
        );

    \I__326\ : Odrv4
    port map (
            O => \N__4379\,
            I => waddr_c_1
        );

    \I__325\ : InMux
    port map (
            O => \N__4376\,
            I => \N__4373\
        );

    \I__324\ : LocalMux
    port map (
            O => \N__4373\,
            I => \N__4369\
        );

    \I__323\ : InMux
    port map (
            O => \N__4372\,
            I => \N__4365\
        );

    \I__322\ : Span4Mux_v
    port map (
            O => \N__4369\,
            I => \N__4362\
        );

    \I__321\ : InMux
    port map (
            O => \N__4368\,
            I => \N__4359\
        );

    \I__320\ : LocalMux
    port map (
            O => \N__4365\,
            I => \N__4356\
        );

    \I__319\ : Span4Mux_v
    port map (
            O => \N__4362\,
            I => \N__4350\
        );

    \I__318\ : LocalMux
    port map (
            O => \N__4359\,
            I => \N__4350\
        );

    \I__317\ : Span4Mux_h
    port map (
            O => \N__4356\,
            I => \N__4346\
        );

    \I__316\ : InMux
    port map (
            O => \N__4355\,
            I => \N__4343\
        );

    \I__315\ : Span4Mux_v
    port map (
            O => \N__4350\,
            I => \N__4340\
        );

    \I__314\ : InMux
    port map (
            O => \N__4349\,
            I => \N__4337\
        );

    \I__313\ : Span4Mux_v
    port map (
            O => \N__4346\,
            I => \N__4334\
        );

    \I__312\ : LocalMux
    port map (
            O => \N__4343\,
            I => \N__4331\
        );

    \I__311\ : Span4Mux_v
    port map (
            O => \N__4340\,
            I => \N__4325\
        );

    \I__310\ : LocalMux
    port map (
            O => \N__4337\,
            I => \N__4325\
        );

    \I__309\ : Span4Mux_v
    port map (
            O => \N__4334\,
            I => \N__4319\
        );

    \I__308\ : Span4Mux_h
    port map (
            O => \N__4331\,
            I => \N__4319\
        );

    \I__307\ : InMux
    port map (
            O => \N__4330\,
            I => \N__4316\
        );

    \I__306\ : Span4Mux_v
    port map (
            O => \N__4325\,
            I => \N__4313\
        );

    \I__305\ : InMux
    port map (
            O => \N__4324\,
            I => \N__4310\
        );

    \I__304\ : Span4Mux_v
    port map (
            O => \N__4319\,
            I => \N__4307\
        );

    \I__303\ : LocalMux
    port map (
            O => \N__4316\,
            I => \N__4304\
        );

    \I__302\ : Span4Mux_v
    port map (
            O => \N__4313\,
            I => \N__4298\
        );

    \I__301\ : LocalMux
    port map (
            O => \N__4310\,
            I => \N__4298\
        );

    \I__300\ : Span4Mux_v
    port map (
            O => \N__4307\,
            I => \N__4293\
        );

    \I__299\ : Span4Mux_h
    port map (
            O => \N__4304\,
            I => \N__4293\
        );

    \I__298\ : InMux
    port map (
            O => \N__4303\,
            I => \N__4290\
        );

    \I__297\ : Span4Mux_v
    port map (
            O => \N__4298\,
            I => \N__4287\
        );

    \I__296\ : Span4Mux_v
    port map (
            O => \N__4293\,
            I => \N__4284\
        );

    \I__295\ : LocalMux
    port map (
            O => \N__4290\,
            I => \N__4281\
        );

    \I__294\ : Sp12to4
    port map (
            O => \N__4287\,
            I => \N__4278\
        );

    \I__293\ : Span4Mux_v
    port map (
            O => \N__4284\,
            I => \N__4273\
        );

    \I__292\ : Span4Mux_h
    port map (
            O => \N__4281\,
            I => \N__4273\
        );

    \I__291\ : Span12Mux_h
    port map (
            O => \N__4278\,
            I => \N__4270\
        );

    \I__290\ : IoSpan4Mux
    port map (
            O => \N__4273\,
            I => \N__4267\
        );

    \I__289\ : Odrv12
    port map (
            O => \N__4270\,
            I => din_c_4
        );

    \I__288\ : Odrv4
    port map (
            O => \N__4267\,
            I => din_c_4
        );

    \I__287\ : InMux
    port map (
            O => \N__4262\,
            I => \N__4258\
        );

    \I__286\ : InMux
    port map (
            O => \N__4261\,
            I => \N__4255\
        );

    \I__285\ : LocalMux
    port map (
            O => \N__4258\,
            I => \N__4252\
        );

    \I__284\ : LocalMux
    port map (
            O => \N__4255\,
            I => \N__4248\
        );

    \I__283\ : Span4Mux_v
    port map (
            O => \N__4252\,
            I => \N__4244\
        );

    \I__282\ : InMux
    port map (
            O => \N__4251\,
            I => \N__4241\
        );

    \I__281\ : Span4Mux_v
    port map (
            O => \N__4248\,
            I => \N__4237\
        );

    \I__280\ : InMux
    port map (
            O => \N__4247\,
            I => \N__4234\
        );

    \I__279\ : Span4Mux_v
    port map (
            O => \N__4244\,
            I => \N__4229\
        );

    \I__278\ : LocalMux
    port map (
            O => \N__4241\,
            I => \N__4229\
        );

    \I__277\ : InMux
    port map (
            O => \N__4240\,
            I => \N__4225\
        );

    \I__276\ : Span4Mux_v
    port map (
            O => \N__4237\,
            I => \N__4220\
        );

    \I__275\ : LocalMux
    port map (
            O => \N__4234\,
            I => \N__4220\
        );

    \I__274\ : Span4Mux_v
    port map (
            O => \N__4229\,
            I => \N__4216\
        );

    \I__273\ : InMux
    port map (
            O => \N__4228\,
            I => \N__4213\
        );

    \I__272\ : LocalMux
    port map (
            O => \N__4225\,
            I => \N__4210\
        );

    \I__271\ : Span4Mux_v
    port map (
            O => \N__4220\,
            I => \N__4207\
        );

    \I__270\ : InMux
    port map (
            O => \N__4219\,
            I => \N__4204\
        );

    \I__269\ : Span4Mux_v
    port map (
            O => \N__4216\,
            I => \N__4199\
        );

    \I__268\ : LocalMux
    port map (
            O => \N__4213\,
            I => \N__4199\
        );

    \I__267\ : Span4Mux_s1_v
    port map (
            O => \N__4210\,
            I => \N__4196\
        );

    \I__266\ : Span4Mux_v
    port map (
            O => \N__4207\,
            I => \N__4191\
        );

    \I__265\ : LocalMux
    port map (
            O => \N__4204\,
            I => \N__4191\
        );

    \I__264\ : Span4Mux_v
    port map (
            O => \N__4199\,
            I => \N__4185\
        );

    \I__263\ : Span4Mux_v
    port map (
            O => \N__4196\,
            I => \N__4185\
        );

    \I__262\ : Span4Mux_v
    port map (
            O => \N__4191\,
            I => \N__4182\
        );

    \I__261\ : InMux
    port map (
            O => \N__4190\,
            I => \N__4179\
        );

    \I__260\ : Sp12to4
    port map (
            O => \N__4185\,
            I => \N__4176\
        );

    \I__259\ : Span4Mux_v
    port map (
            O => \N__4182\,
            I => \N__4171\
        );

    \I__258\ : LocalMux
    port map (
            O => \N__4179\,
            I => \N__4171\
        );

    \I__257\ : Span12Mux_h
    port map (
            O => \N__4176\,
            I => \N__4168\
        );

    \I__256\ : IoSpan4Mux
    port map (
            O => \N__4171\,
            I => \N__4165\
        );

    \I__255\ : Span12Mux_h
    port map (
            O => \N__4168\,
            I => \N__4162\
        );

    \I__254\ : IoSpan4Mux
    port map (
            O => \N__4165\,
            I => \N__4159\
        );

    \I__253\ : Odrv12
    port map (
            O => \N__4162\,
            I => din_c_6
        );

    \I__252\ : Odrv4
    port map (
            O => \N__4159\,
            I => din_c_6
        );

    \I__251\ : InMux
    port map (
            O => \N__4154\,
            I => \N__4151\
        );

    \I__250\ : LocalMux
    port map (
            O => \N__4151\,
            I => \N__4148\
        );

    \I__249\ : Span4Mux_v
    port map (
            O => \N__4148\,
            I => \N__4141\
        );

    \I__248\ : InMux
    port map (
            O => \N__4147\,
            I => \N__4138\
        );

    \I__247\ : InMux
    port map (
            O => \N__4146\,
            I => \N__4135\
        );

    \I__246\ : InMux
    port map (
            O => \N__4145\,
            I => \N__4132\
        );

    \I__245\ : InMux
    port map (
            O => \N__4144\,
            I => \N__4128\
        );

    \I__244\ : Span4Mux_v
    port map (
            O => \N__4141\,
            I => \N__4123\
        );

    \I__243\ : LocalMux
    port map (
            O => \N__4138\,
            I => \N__4123\
        );

    \I__242\ : LocalMux
    port map (
            O => \N__4135\,
            I => \N__4119\
        );

    \I__241\ : LocalMux
    port map (
            O => \N__4132\,
            I => \N__4116\
        );

    \I__240\ : InMux
    port map (
            O => \N__4131\,
            I => \N__4113\
        );

    \I__239\ : LocalMux
    port map (
            O => \N__4128\,
            I => \N__4110\
        );

    \I__238\ : Span4Mux_v
    port map (
            O => \N__4123\,
            I => \N__4107\
        );

    \I__237\ : InMux
    port map (
            O => \N__4122\,
            I => \N__4104\
        );

    \I__236\ : Span12Mux_v
    port map (
            O => \N__4119\,
            I => \N__4100\
        );

    \I__235\ : Sp12to4
    port map (
            O => \N__4116\,
            I => \N__4095\
        );

    \I__234\ : LocalMux
    port map (
            O => \N__4113\,
            I => \N__4095\
        );

    \I__233\ : Sp12to4
    port map (
            O => \N__4110\,
            I => \N__4092\
        );

    \I__232\ : Span4Mux_v
    port map (
            O => \N__4107\,
            I => \N__4087\
        );

    \I__231\ : LocalMux
    port map (
            O => \N__4104\,
            I => \N__4087\
        );

    \I__230\ : InMux
    port map (
            O => \N__4103\,
            I => \N__4084\
        );

    \I__229\ : Span12Mux_h
    port map (
            O => \N__4100\,
            I => \N__4081\
        );

    \I__228\ : Span12Mux_v
    port map (
            O => \N__4095\,
            I => \N__4076\
        );

    \I__227\ : Span12Mux_s4_v
    port map (
            O => \N__4092\,
            I => \N__4076\
        );

    \I__226\ : Span4Mux_v
    port map (
            O => \N__4087\,
            I => \N__4073\
        );

    \I__225\ : LocalMux
    port map (
            O => \N__4084\,
            I => \N__4070\
        );

    \I__224\ : Span12Mux_h
    port map (
            O => \N__4081\,
            I => \N__4067\
        );

    \I__223\ : Span12Mux_h
    port map (
            O => \N__4076\,
            I => \N__4064\
        );

    \I__222\ : Span4Mux_v
    port map (
            O => \N__4073\,
            I => \N__4059\
        );

    \I__221\ : Span4Mux_v
    port map (
            O => \N__4070\,
            I => \N__4059\
        );

    \I__220\ : Span12Mux_v
    port map (
            O => \N__4067\,
            I => \N__4054\
        );

    \I__219\ : Span12Mux_h
    port map (
            O => \N__4064\,
            I => \N__4054\
        );

    \I__218\ : Span4Mux_h
    port map (
            O => \N__4059\,
            I => \N__4051\
        );

    \I__217\ : Odrv12
    port map (
            O => \N__4054\,
            I => din_c_7
        );

    \I__216\ : Odrv4
    port map (
            O => \N__4051\,
            I => din_c_7
        );

    \I__215\ : InMux
    port map (
            O => \N__4046\,
            I => \N__4043\
        );

    \I__214\ : LocalMux
    port map (
            O => \N__4043\,
            I => \N__4040\
        );

    \I__213\ : Span4Mux_v
    port map (
            O => \N__4040\,
            I => \N__4036\
        );

    \I__212\ : InMux
    port map (
            O => \N__4039\,
            I => \N__4033\
        );

    \I__211\ : Span4Mux_v
    port map (
            O => \N__4036\,
            I => \N__4028\
        );

    \I__210\ : LocalMux
    port map (
            O => \N__4033\,
            I => \N__4028\
        );

    \I__209\ : Span4Mux_v
    port map (
            O => \N__4028\,
            I => \N__4024\
        );

    \I__208\ : InMux
    port map (
            O => \N__4027\,
            I => \N__4021\
        );

    \I__207\ : Span4Mux_v
    port map (
            O => \N__4024\,
            I => \N__4016\
        );

    \I__206\ : LocalMux
    port map (
            O => \N__4021\,
            I => \N__4016\
        );

    \I__205\ : Span4Mux_v
    port map (
            O => \N__4016\,
            I => \N__4011\
        );

    \I__204\ : InMux
    port map (
            O => \N__4015\,
            I => \N__4008\
        );

    \I__203\ : InMux
    port map (
            O => \N__4014\,
            I => \N__4004\
        );

    \I__202\ : Span4Mux_v
    port map (
            O => \N__4011\,
            I => \N__3999\
        );

    \I__201\ : LocalMux
    port map (
            O => \N__4008\,
            I => \N__3999\
        );

    \I__200\ : InMux
    port map (
            O => \N__4007\,
            I => \N__3995\
        );

    \I__199\ : LocalMux
    port map (
            O => \N__4004\,
            I => \N__3992\
        );

    \I__198\ : Span4Mux_v
    port map (
            O => \N__3999\,
            I => \N__3989\
        );

    \I__197\ : InMux
    port map (
            O => \N__3998\,
            I => \N__3986\
        );

    \I__196\ : LocalMux
    port map (
            O => \N__3995\,
            I => \N__3983\
        );

    \I__195\ : Sp12to4
    port map (
            O => \N__3992\,
            I => \N__3979\
        );

    \I__194\ : Span4Mux_h
    port map (
            O => \N__3989\,
            I => \N__3976\
        );

    \I__193\ : LocalMux
    port map (
            O => \N__3986\,
            I => \N__3973\
        );

    \I__192\ : Span4Mux_v
    port map (
            O => \N__3983\,
            I => \N__3970\
        );

    \I__191\ : InMux
    port map (
            O => \N__3982\,
            I => \N__3967\
        );

    \I__190\ : Span12Mux_v
    port map (
            O => \N__3979\,
            I => \N__3964\
        );

    \I__189\ : Sp12to4
    port map (
            O => \N__3976\,
            I => \N__3961\
        );

    \I__188\ : Sp12to4
    port map (
            O => \N__3973\,
            I => \N__3958\
        );

    \I__187\ : Span4Mux_v
    port map (
            O => \N__3970\,
            I => \N__3953\
        );

    \I__186\ : LocalMux
    port map (
            O => \N__3967\,
            I => \N__3953\
        );

    \I__185\ : Span12Mux_v
    port map (
            O => \N__3964\,
            I => \N__3950\
        );

    \I__184\ : Span12Mux_h
    port map (
            O => \N__3961\,
            I => \N__3947\
        );

    \I__183\ : Span12Mux_v
    port map (
            O => \N__3958\,
            I => \N__3944\
        );

    \I__182\ : Span4Mux_v
    port map (
            O => \N__3953\,
            I => \N__3941\
        );

    \I__181\ : Odrv12
    port map (
            O => \N__3950\,
            I => din_c_3
        );

    \I__180\ : Odrv12
    port map (
            O => \N__3947\,
            I => din_c_3
        );

    \I__179\ : Odrv12
    port map (
            O => \N__3944\,
            I => din_c_3
        );

    \I__178\ : Odrv4
    port map (
            O => \N__3941\,
            I => din_c_3
        );

    \I__177\ : InMux
    port map (
            O => \N__3932\,
            I => \N__3929\
        );

    \I__176\ : LocalMux
    port map (
            O => \N__3929\,
            I => \N__3926\
        );

    \I__175\ : Span4Mux_v
    port map (
            O => \N__3926\,
            I => \N__3922\
        );

    \I__174\ : InMux
    port map (
            O => \N__3925\,
            I => \N__3919\
        );

    \I__173\ : Span4Mux_v
    port map (
            O => \N__3922\,
            I => \N__3914\
        );

    \I__172\ : LocalMux
    port map (
            O => \N__3919\,
            I => \N__3914\
        );

    \I__171\ : Span4Mux_v
    port map (
            O => \N__3914\,
            I => \N__3910\
        );

    \I__170\ : InMux
    port map (
            O => \N__3913\,
            I => \N__3907\
        );

    \I__169\ : Span4Mux_v
    port map (
            O => \N__3910\,
            I => \N__3901\
        );

    \I__168\ : LocalMux
    port map (
            O => \N__3907\,
            I => \N__3901\
        );

    \I__167\ : InMux
    port map (
            O => \N__3906\,
            I => \N__3898\
        );

    \I__166\ : Span4Mux_v
    port map (
            O => \N__3901\,
            I => \N__3895\
        );

    \I__165\ : LocalMux
    port map (
            O => \N__3898\,
            I => \N__3892\
        );

    \I__164\ : Span4Mux_v
    port map (
            O => \N__3895\,
            I => \N__3885\
        );

    \I__163\ : Span4Mux_v
    port map (
            O => \N__3892\,
            I => \N__3885\
        );

    \I__162\ : InMux
    port map (
            O => \N__3891\,
            I => \N__3882\
        );

    \I__161\ : InMux
    port map (
            O => \N__3890\,
            I => \N__3878\
        );

    \I__160\ : Span4Mux_h
    port map (
            O => \N__3885\,
            I => \N__3875\
        );

    \I__159\ : LocalMux
    port map (
            O => \N__3882\,
            I => \N__3872\
        );

    \I__158\ : InMux
    port map (
            O => \N__3881\,
            I => \N__3869\
        );

    \I__157\ : LocalMux
    port map (
            O => \N__3878\,
            I => \N__3865\
        );

    \I__156\ : Sp12to4
    port map (
            O => \N__3875\,
            I => \N__3862\
        );

    \I__155\ : Span12Mux_v
    port map (
            O => \N__3872\,
            I => \N__3857\
        );

    \I__154\ : LocalMux
    port map (
            O => \N__3869\,
            I => \N__3857\
        );

    \I__153\ : InMux
    port map (
            O => \N__3868\,
            I => \N__3854\
        );

    \I__152\ : Span12Mux_v
    port map (
            O => \N__3865\,
            I => \N__3851\
        );

    \I__151\ : Span12Mux_h
    port map (
            O => \N__3862\,
            I => \N__3844\
        );

    \I__150\ : Span12Mux_v
    port map (
            O => \N__3857\,
            I => \N__3844\
        );

    \I__149\ : LocalMux
    port map (
            O => \N__3854\,
            I => \N__3844\
        );

    \I__148\ : Odrv12
    port map (
            O => \N__3851\,
            I => din_c_2
        );

    \I__147\ : Odrv12
    port map (
            O => \N__3844\,
            I => din_c_2
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \waddr_ibuf_RNIO66O1_0_11_LC_7_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__10057\,
            in1 => \N__10093\,
            in2 => \N__9977\,
            in3 => \N__10009\,
            lcout => \mem_WE_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \waddr_ibuf_RNIO66O1_11_LC_7_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__10094\,
            in1 => \N__10058\,
            in2 => \N__10025\,
            in3 => \N__9964\,
            lcout => \mem_WE_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \waddr_ibuf_RNIO66O1_1_11_LC_7_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__10059\,
            in1 => \N__10095\,
            in2 => \N__9978\,
            in3 => \N__10013\,
            lcout => \mem_WE_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \waddr_ibuf_RNIO66O1_2_11_LC_7_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__10096\,
            in1 => \N__10060\,
            in2 => \N__10026\,
            in3 => \N__9968\,
            lcout => \mem_WE_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \waddr_ibuf_RNIO66O1_3_11_LC_7_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__10061\,
            in1 => \N__10097\,
            in2 => \N__9979\,
            in3 => \N__10017\,
            lcout => \mem_WE_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \waddr_ibuf_RNIO66O1_4_11_LC_7_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__10098\,
            in1 => \N__10062\,
            in2 => \N__10027\,
            in3 => \N__9972\,
            lcout => \mem_WE_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \waddr_ibuf_RNIO66O1_5_11_LC_7_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__10063\,
            in1 => \N__10099\,
            in2 => \N__9980\,
            in3 => \N__10021\,
            lcout => \mem_WE_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \waddr_ibuf_RNIO66O1_6_11_LC_7_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__10100\,
            in1 => \N__10064\,
            in2 => \N__10028\,
            in3 => \N__9976\,
            lcout => \mem_WE_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_4_0_LC_10_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9896\,
            in1 => \N__12430\,
            in2 => \_gnd_net_\,
            in3 => \N__9878\,
            lcout => \dout_obuf_RNO_4Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_4_1_LC_10_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__9866\,
            in1 => \N__12431\,
            in2 => \_gnd_net_\,
            in3 => \N__9851\,
            lcout => \dout_obuf_RNO_4Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_4_7_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__9842\,
            in1 => \_gnd_net_\,
            in2 => \N__12364\,
            in3 => \N__9833\,
            lcout => \dout_obuf_RNO_4Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_4_6_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__11030\,
            in1 => \N__12345\,
            in2 => \_gnd_net_\,
            in3 => \N__11012\,
            lcout => \dout_obuf_RNO_4Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_2_1_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__10439\,
            in1 => \N__12414\,
            in2 => \_gnd_net_\,
            in3 => \N__10430\,
            lcout => \dout_obuf_RNO_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_2_0_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__10415\,
            in1 => \N__12413\,
            in2 => \_gnd_net_\,
            in3 => \N__10403\,
            lcout => \dout_obuf_RNO_2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_1_1_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__11414\,
            in1 => \N__12755\,
            in2 => \_gnd_net_\,
            in3 => \N__10385\,
            lcout => OPEN,
            ltout => \mem_N_162_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_1_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__11162\,
            in1 => \_gnd_net_\,
            in2 => \N__10373\,
            in3 => \N__12584\,
            lcout => dout_c_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_1_0_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__12751\,
            in1 => \N__11372\,
            in2 => \_gnd_net_\,
            in3 => \N__10358\,
            lcout => OPEN,
            ltout => \mem_N_156_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_0_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12559\,
            in2 => \N__10346\,
            in3 => \N__11147\,
            lcout => dout_c_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_0_1_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__12011\,
            in1 => \N__12750\,
            in2 => \_gnd_net_\,
            in3 => \N__11171\,
            lcout => \mem_N_160\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_0_0_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__11156\,
            in1 => \N__12749\,
            in2 => \_gnd_net_\,
            in3 => \N__11303\,
            lcout => \mem_N_154\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_2_2_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__11141\,
            in1 => \N__12328\,
            in2 => \_gnd_net_\,
            in3 => \N__11129\,
            lcout => \dout_obuf_RNO_2Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_0_2_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__11261\,
            in1 => \N__12730\,
            in2 => \_gnd_net_\,
            in3 => \N__11111\,
            lcout => OPEN,
            ltout => \mem_N_166_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_2_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12580\,
            in2 => \N__11105\,
            in3 => \N__11795\,
            lcout => dout_c_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_1_7_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__12715\,
            in1 => \N__12047\,
            in2 => \_gnd_net_\,
            in3 => \N__11093\,
            lcout => \mem_N_150\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_2_7_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__11084\,
            in1 => \N__12321\,
            in2 => \_gnd_net_\,
            in3 => \N__11075\,
            lcout => OPEN,
            ltout => \dout_obuf_RNO_2Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_0_7_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12714\,
            in2 => \N__11060\,
            in3 => \N__11924\,
            lcout => OPEN,
            ltout => \mem_N_149_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_7_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__11057\,
            in1 => \_gnd_net_\,
            in2 => \N__11051\,
            in3 => \N__12560\,
            lcout => dout_c_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_5_1_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__11438\,
            in1 => \_gnd_net_\,
            in2 => \N__12400\,
            in3 => \N__11423\,
            lcout => \dout_obuf_RNO_5Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_5_0_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__11402\,
            in1 => \N__12384\,
            in2 => \_gnd_net_\,
            in3 => \N__11390\,
            lcout => \dout_obuf_RNO_5Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_5_3_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__11363\,
            in1 => \_gnd_net_\,
            in2 => \N__12401\,
            in3 => \N__11351\,
            lcout => \dout_obuf_RNO_5Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_3_0_LC_10_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__11333\,
            in1 => \N__12358\,
            in2 => \_gnd_net_\,
            in3 => \N__11321\,
            lcout => \dout_obuf_RNO_3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_3_2_LC_10_27_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__11291\,
            in1 => \N__12278\,
            in2 => \_gnd_net_\,
            in3 => \N__11279\,
            lcout => \dout_obuf_RNO_3Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_3_3_LC_10_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__11246\,
            in1 => \N__12279\,
            in2 => \_gnd_net_\,
            in3 => \N__11237\,
            lcout => \dout_obuf_RNO_3Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_4_2_LC_11_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__11222\,
            in1 => \N__12349\,
            in2 => \_gnd_net_\,
            in3 => \N__11210\,
            lcout => \dout_obuf_RNO_4Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_4_3_LC_11_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__11192\,
            in1 => \N__12350\,
            in2 => \_gnd_net_\,
            in3 => \N__11183\,
            lcout => \dout_obuf_RNO_4Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_4_5_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__11618\,
            in1 => \N__12424\,
            in2 => \_gnd_net_\,
            in3 => \N__11609\,
            lcout => \dout_obuf_RNO_4Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_4_4_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__11597\,
            in1 => \N__12423\,
            in2 => \_gnd_net_\,
            in3 => \N__11579\,
            lcout => \dout_obuf_RNO_4Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_1_4_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__11669\,
            in1 => \N__12728\,
            in2 => \_gnd_net_\,
            in3 => \N__11567\,
            lcout => OPEN,
            ltout => \mem_N_180_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_4_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__12578\,
            in1 => \_gnd_net_\,
            in2 => \N__11555\,
            in3 => \N__11756\,
            lcout => dout_c_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_1_6_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__12729\,
            in1 => \N__12080\,
            in2 => \_gnd_net_\,
            in3 => \N__11534\,
            lcout => OPEN,
            ltout => \mem_N_145_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_6_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__12579\,
            in1 => \_gnd_net_\,
            in2 => \N__11525\,
            in3 => \N__11711\,
            lcout => dout_c_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_1_3_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__12748\,
            in1 => \N__11504\,
            in2 => \_gnd_net_\,
            in3 => \N__11492\,
            lcout => \mem_N_174\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_2_3_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__11480\,
            in1 => \N__12327\,
            in2 => \_gnd_net_\,
            in3 => \N__11471\,
            lcout => OPEN,
            ltout => \dout_obuf_RNO_2Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_0_3_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__11456\,
            in1 => \_gnd_net_\,
            in2 => \N__11441\,
            in3 => \N__12747\,
            lcout => OPEN,
            ltout => \mem_N_172_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_3_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__11828\,
            in1 => \_gnd_net_\,
            in2 => \N__11822\,
            in3 => \N__12558\,
            lcout => dout_c_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_1_2_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__12712\,
            in1 => \N__11627\,
            in2 => \_gnd_net_\,
            in3 => \N__11807\,
            lcout => \mem_N_168\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_2_4_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__11789\,
            in1 => \N__12402\,
            in2 => \_gnd_net_\,
            in3 => \N__11771\,
            lcout => OPEN,
            ltout => \dout_obuf_RNO_2Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_0_4_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__12711\,
            in1 => \_gnd_net_\,
            in2 => \N__11759\,
            in3 => \N__11966\,
            lcout => \mem_N_178\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_2_6_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__11744\,
            in1 => \N__12320\,
            in2 => \_gnd_net_\,
            in3 => \N__11726\,
            lcout => OPEN,
            ltout => \dout_obuf_RNO_2Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_0_6_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__12713\,
            in1 => \_gnd_net_\,
            in2 => \N__11714\,
            in3 => \N__11879\,
            lcout => \mem_N_144\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_5_4_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__12314\,
            in1 => \N__11699\,
            in2 => \_gnd_net_\,
            in3 => \N__11687\,
            lcout => \dout_obuf_RNO_5Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_5_2_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__11657\,
            in1 => \N__12313\,
            in2 => \_gnd_net_\,
            in3 => \N__11639\,
            lcout => \dout_obuf_RNO_5Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_5_6_LC_11_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__12289\,
            in1 => \N__12110\,
            in2 => \_gnd_net_\,
            in3 => \N__12098\,
            lcout => \dout_obuf_RNO_5Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_5_7_LC_11_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__12290\,
            in1 => \N__12068\,
            in2 => \_gnd_net_\,
            in3 => \N__12059\,
            lcout => \dout_obuf_RNO_5Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_3_1_LC_11_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__12032\,
            in1 => \N__12357\,
            in2 => \_gnd_net_\,
            in3 => \N__12023\,
            lcout => \dout_obuf_RNO_3Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_3_4_LC_11_29_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__12335\,
            in1 => \N__11996\,
            in2 => \_gnd_net_\,
            in3 => \N__11984\,
            lcout => \dout_obuf_RNO_3Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_3_7_LC_11_31_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__12264\,
            in1 => \N__11945\,
            in2 => \_gnd_net_\,
            in3 => \N__11936\,
            lcout => \dout_obuf_RNO_3Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_3_6_LC_11_31_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__11909\,
            in1 => \N__12263\,
            in2 => \_gnd_net_\,
            in3 => \N__11897\,
            lcout => \dout_obuf_RNO_3Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_1_5_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__12440\,
            in1 => \N__12684\,
            in2 => \_gnd_net_\,
            in3 => \N__11861\,
            lcout => \mem_N_140\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_2_5_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__11849\,
            in1 => \N__12399\,
            in2 => \_gnd_net_\,
            in3 => \N__11837\,
            lcout => OPEN,
            ltout => \dout_obuf_RNO_2Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_0_5_LC_13_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__12683\,
            in1 => \_gnd_net_\,
            in2 => \N__12593\,
            in3 => \N__12122\,
            lcout => \mem_N_139\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_5_LC_13_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__12590\,
            in1 => \N__12566\,
            in2 => \_gnd_net_\,
            in3 => \N__12488\,
            lcout => dout_c_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_5_5_LC_13_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__12365\,
            in1 => \N__12461\,
            in2 => \_gnd_net_\,
            in3 => \N__12452\,
            lcout => \dout_obuf_RNO_5Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dout_obuf_RNO_3_5_LC_13_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__12329\,
            in1 => \N__12143\,
            in2 => \_gnd_net_\,
            in3 => \N__12134\,
            lcout => \dout_obuf_RNO_3Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
