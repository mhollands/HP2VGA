// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     Sep 29 2018 12:24:33

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "main" view "INTERFACE"

module main (
    TVP_VIDEO,
    ADV_B,
    ADV_G,
    ADV_R,
    DEBUG,
    TVP_CLK,
    ADV_CLK,
    TVP_HSYNC,
    ADV_HSYNC,
    TVP_VSYNC,
    ADV_VSYNC,
    ADV_BLANK_N,
    LED,
    ADV_SYNC_N);

    input [9:0] TVP_VIDEO;
    output [7:0] ADV_B;
    output [7:0] ADV_G;
    output [7:0] ADV_R;
    inout [7:0] DEBUG;
    input TVP_CLK;
    output ADV_CLK;
    input TVP_HSYNC;
    output ADV_HSYNC;
    input TVP_VSYNC;
    output ADV_VSYNC;
    output ADV_BLANK_N;
    output LED;
    output ADV_SYNC_N;

    wire N__24121;
    wire N__24120;
    wire N__24119;
    wire N__24110;
    wire N__24109;
    wire N__24108;
    wire N__24101;
    wire N__24100;
    wire N__24099;
    wire N__24092;
    wire N__24091;
    wire N__24090;
    wire N__24083;
    wire N__24082;
    wire N__24081;
    wire N__24074;
    wire N__24073;
    wire N__24072;
    wire N__24065;
    wire N__24064;
    wire N__24063;
    wire N__24056;
    wire N__24055;
    wire N__24054;
    wire N__24047;
    wire N__24046;
    wire N__24045;
    wire N__24038;
    wire N__24037;
    wire N__24036;
    wire N__24029;
    wire N__24028;
    wire N__24027;
    wire N__24020;
    wire N__24019;
    wire N__24018;
    wire N__24011;
    wire N__24010;
    wire N__24009;
    wire N__24002;
    wire N__24001;
    wire N__24000;
    wire N__23993;
    wire N__23992;
    wire N__23991;
    wire N__23984;
    wire N__23983;
    wire N__23982;
    wire N__23975;
    wire N__23974;
    wire N__23973;
    wire N__23966;
    wire N__23965;
    wire N__23964;
    wire N__23957;
    wire N__23956;
    wire N__23955;
    wire N__23948;
    wire N__23947;
    wire N__23946;
    wire N__23939;
    wire N__23938;
    wire N__23937;
    wire N__23930;
    wire N__23929;
    wire N__23928;
    wire N__23921;
    wire N__23920;
    wire N__23919;
    wire N__23912;
    wire N__23911;
    wire N__23910;
    wire N__23903;
    wire N__23902;
    wire N__23901;
    wire N__23894;
    wire N__23893;
    wire N__23892;
    wire N__23885;
    wire N__23884;
    wire N__23883;
    wire N__23876;
    wire N__23875;
    wire N__23874;
    wire N__23867;
    wire N__23866;
    wire N__23865;
    wire N__23858;
    wire N__23857;
    wire N__23856;
    wire N__23849;
    wire N__23848;
    wire N__23847;
    wire N__23840;
    wire N__23839;
    wire N__23838;
    wire N__23831;
    wire N__23830;
    wire N__23829;
    wire N__23822;
    wire N__23821;
    wire N__23820;
    wire N__23813;
    wire N__23812;
    wire N__23811;
    wire N__23804;
    wire N__23803;
    wire N__23802;
    wire N__23795;
    wire N__23794;
    wire N__23793;
    wire N__23786;
    wire N__23785;
    wire N__23784;
    wire N__23777;
    wire N__23776;
    wire N__23775;
    wire N__23768;
    wire N__23767;
    wire N__23766;
    wire N__23759;
    wire N__23758;
    wire N__23757;
    wire N__23750;
    wire N__23749;
    wire N__23748;
    wire N__23741;
    wire N__23740;
    wire N__23739;
    wire N__23732;
    wire N__23731;
    wire N__23730;
    wire N__23723;
    wire N__23722;
    wire N__23721;
    wire N__23714;
    wire N__23713;
    wire N__23712;
    wire N__23705;
    wire N__23704;
    wire N__23703;
    wire N__23696;
    wire N__23695;
    wire N__23694;
    wire N__23687;
    wire N__23686;
    wire N__23685;
    wire N__23668;
    wire N__23667;
    wire N__23666;
    wire N__23665;
    wire N__23664;
    wire N__23663;
    wire N__23660;
    wire N__23659;
    wire N__23656;
    wire N__23655;
    wire N__23654;
    wire N__23653;
    wire N__23650;
    wire N__23649;
    wire N__23648;
    wire N__23647;
    wire N__23644;
    wire N__23641;
    wire N__23640;
    wire N__23639;
    wire N__23638;
    wire N__23637;
    wire N__23634;
    wire N__23631;
    wire N__23630;
    wire N__23629;
    wire N__23626;
    wire N__23623;
    wire N__23620;
    wire N__23617;
    wire N__23614;
    wire N__23609;
    wire N__23606;
    wire N__23603;
    wire N__23602;
    wire N__23601;
    wire N__23596;
    wire N__23593;
    wire N__23590;
    wire N__23587;
    wire N__23584;
    wire N__23581;
    wire N__23578;
    wire N__23575;
    wire N__23574;
    wire N__23571;
    wire N__23564;
    wire N__23561;
    wire N__23554;
    wire N__23551;
    wire N__23548;
    wire N__23545;
    wire N__23544;
    wire N__23543;
    wire N__23536;
    wire N__23529;
    wire N__23524;
    wire N__23521;
    wire N__23516;
    wire N__23507;
    wire N__23504;
    wire N__23501;
    wire N__23498;
    wire N__23489;
    wire N__23484;
    wire N__23473;
    wire N__23470;
    wire N__23467;
    wire N__23464;
    wire N__23461;
    wire N__23458;
    wire N__23455;
    wire N__23452;
    wire N__23449;
    wire N__23446;
    wire N__23443;
    wire N__23440;
    wire N__23437;
    wire N__23434;
    wire N__23431;
    wire N__23428;
    wire N__23425;
    wire N__23424;
    wire N__23421;
    wire N__23418;
    wire N__23417;
    wire N__23412;
    wire N__23409;
    wire N__23406;
    wire N__23403;
    wire N__23400;
    wire N__23397;
    wire N__23394;
    wire N__23391;
    wire N__23388;
    wire N__23385;
    wire N__23382;
    wire N__23379;
    wire N__23374;
    wire N__23371;
    wire N__23368;
    wire N__23365;
    wire N__23364;
    wire N__23361;
    wire N__23358;
    wire N__23357;
    wire N__23354;
    wire N__23351;
    wire N__23348;
    wire N__23345;
    wire N__23342;
    wire N__23339;
    wire N__23336;
    wire N__23333;
    wire N__23330;
    wire N__23327;
    wire N__23324;
    wire N__23321;
    wire N__23318;
    wire N__23315;
    wire N__23312;
    wire N__23305;
    wire N__23302;
    wire N__23301;
    wire N__23298;
    wire N__23295;
    wire N__23294;
    wire N__23293;
    wire N__23292;
    wire N__23289;
    wire N__23286;
    wire N__23283;
    wire N__23280;
    wire N__23279;
    wire N__23278;
    wire N__23275;
    wire N__23274;
    wire N__23273;
    wire N__23272;
    wire N__23271;
    wire N__23270;
    wire N__23269;
    wire N__23268;
    wire N__23261;
    wire N__23258;
    wire N__23255;
    wire N__23252;
    wire N__23251;
    wire N__23248;
    wire N__23245;
    wire N__23242;
    wire N__23239;
    wire N__23236;
    wire N__23235;
    wire N__23232;
    wire N__23229;
    wire N__23226;
    wire N__23225;
    wire N__23224;
    wire N__23217;
    wire N__23214;
    wire N__23211;
    wire N__23204;
    wire N__23203;
    wire N__23202;
    wire N__23201;
    wire N__23200;
    wire N__23199;
    wire N__23194;
    wire N__23191;
    wire N__23190;
    wire N__23189;
    wire N__23182;
    wire N__23179;
    wire N__23176;
    wire N__23175;
    wire N__23174;
    wire N__23167;
    wire N__23164;
    wire N__23161;
    wire N__23160;
    wire N__23159;
    wire N__23156;
    wire N__23153;
    wire N__23152;
    wire N__23151;
    wire N__23148;
    wire N__23145;
    wire N__23144;
    wire N__23143;
    wire N__23138;
    wire N__23135;
    wire N__23134;
    wire N__23131;
    wire N__23130;
    wire N__23125;
    wire N__23122;
    wire N__23119;
    wire N__23116;
    wire N__23113;
    wire N__23108;
    wire N__23107;
    wire N__23106;
    wire N__23105;
    wire N__23102;
    wire N__23101;
    wire N__23100;
    wire N__23097;
    wire N__23096;
    wire N__23091;
    wire N__23088;
    wire N__23087;
    wire N__23086;
    wire N__23083;
    wire N__23082;
    wire N__23081;
    wire N__23080;
    wire N__23079;
    wire N__23078;
    wire N__23077;
    wire N__23074;
    wire N__23073;
    wire N__23070;
    wire N__23067;
    wire N__23064;
    wire N__23059;
    wire N__23056;
    wire N__23055;
    wire N__23052;
    wire N__23049;
    wire N__23042;
    wire N__23039;
    wire N__23034;
    wire N__23031;
    wire N__23028;
    wire N__23027;
    wire N__23026;
    wire N__23023;
    wire N__23020;
    wire N__23017;
    wire N__23014;
    wire N__23011;
    wire N__23008;
    wire N__23005;
    wire N__23002;
    wire N__22999;
    wire N__22998;
    wire N__22997;
    wire N__22996;
    wire N__22995;
    wire N__22994;
    wire N__22991;
    wire N__22990;
    wire N__22989;
    wire N__22986;
    wire N__22983;
    wire N__22982;
    wire N__22981;
    wire N__22980;
    wire N__22979;
    wire N__22976;
    wire N__22973;
    wire N__22972;
    wire N__22969;
    wire N__22968;
    wire N__22965;
    wire N__22962;
    wire N__22961;
    wire N__22958;
    wire N__22955;
    wire N__22948;
    wire N__22947;
    wire N__22942;
    wire N__22939;
    wire N__22938;
    wire N__22933;
    wire N__22932;
    wire N__22923;
    wire N__22920;
    wire N__22917;
    wire N__22914;
    wire N__22913;
    wire N__22912;
    wire N__22909;
    wire N__22902;
    wire N__22897;
    wire N__22890;
    wire N__22887;
    wire N__22884;
    wire N__22883;
    wire N__22882;
    wire N__22879;
    wire N__22876;
    wire N__22873;
    wire N__22872;
    wire N__22869;
    wire N__22866;
    wire N__22863;
    wire N__22858;
    wire N__22855;
    wire N__22854;
    wire N__22853;
    wire N__22850;
    wire N__22847;
    wire N__22844;
    wire N__22843;
    wire N__22840;
    wire N__22837;
    wire N__22834;
    wire N__22833;
    wire N__22832;
    wire N__22829;
    wire N__22826;
    wire N__22825;
    wire N__22824;
    wire N__22821;
    wire N__22818;
    wire N__22815;
    wire N__22810;
    wire N__22809;
    wire N__22806;
    wire N__22803;
    wire N__22800;
    wire N__22797;
    wire N__22794;
    wire N__22791;
    wire N__22788;
    wire N__22785;
    wire N__22780;
    wire N__22777;
    wire N__22774;
    wire N__22771;
    wire N__22770;
    wire N__22765;
    wire N__22758;
    wire N__22755;
    wire N__22752;
    wire N__22751;
    wire N__22748;
    wire N__22747;
    wire N__22746;
    wire N__22743;
    wire N__22738;
    wire N__22735;
    wire N__22728;
    wire N__22723;
    wire N__22720;
    wire N__22717;
    wire N__22714;
    wire N__22711;
    wire N__22708;
    wire N__22705;
    wire N__22698;
    wire N__22695;
    wire N__22694;
    wire N__22691;
    wire N__22690;
    wire N__22685;
    wire N__22682;
    wire N__22679;
    wire N__22670;
    wire N__22667;
    wire N__22662;
    wire N__22651;
    wire N__22650;
    wire N__22649;
    wire N__22646;
    wire N__22639;
    wire N__22636;
    wire N__22633;
    wire N__22632;
    wire N__22623;
    wire N__22620;
    wire N__22617;
    wire N__22614;
    wire N__22611;
    wire N__22610;
    wire N__22603;
    wire N__22594;
    wire N__22585;
    wire N__22580;
    wire N__22577;
    wire N__22574;
    wire N__22571;
    wire N__22566;
    wire N__22559;
    wire N__22558;
    wire N__22557;
    wire N__22552;
    wire N__22549;
    wire N__22546;
    wire N__22545;
    wire N__22542;
    wire N__22535;
    wire N__22532;
    wire N__22531;
    wire N__22530;
    wire N__22525;
    wire N__22520;
    wire N__22517;
    wire N__22514;
    wire N__22503;
    wire N__22498;
    wire N__22497;
    wire N__22492;
    wire N__22489;
    wire N__22486;
    wire N__22483;
    wire N__22480;
    wire N__22477;
    wire N__22474;
    wire N__22471;
    wire N__22468;
    wire N__22465;
    wire N__22462;
    wire N__22461;
    wire N__22458;
    wire N__22453;
    wire N__22450;
    wire N__22447;
    wire N__22442;
    wire N__22439;
    wire N__22434;
    wire N__22431;
    wire N__22426;
    wire N__22423;
    wire N__22420;
    wire N__22415;
    wire N__22412;
    wire N__22409;
    wire N__22406;
    wire N__22403;
    wire N__22400;
    wire N__22395;
    wire N__22392;
    wire N__22389;
    wire N__22384;
    wire N__22381;
    wire N__22376;
    wire N__22369;
    wire N__22366;
    wire N__22363;
    wire N__22358;
    wire N__22355;
    wire N__22350;
    wire N__22347;
    wire N__22340;
    wire N__22327;
    wire N__22326;
    wire N__22323;
    wire N__22322;
    wire N__22321;
    wire N__22320;
    wire N__22319;
    wire N__22316;
    wire N__22315;
    wire N__22312;
    wire N__22309;
    wire N__22306;
    wire N__22303;
    wire N__22300;
    wire N__22297;
    wire N__22294;
    wire N__22289;
    wire N__22286;
    wire N__22283;
    wire N__22280;
    wire N__22275;
    wire N__22272;
    wire N__22267;
    wire N__22264;
    wire N__22261;
    wire N__22252;
    wire N__22249;
    wire N__22246;
    wire N__22243;
    wire N__22240;
    wire N__22237;
    wire N__22236;
    wire N__22235;
    wire N__22234;
    wire N__22233;
    wire N__22232;
    wire N__22231;
    wire N__22228;
    wire N__22227;
    wire N__22226;
    wire N__22225;
    wire N__22222;
    wire N__22219;
    wire N__22218;
    wire N__22217;
    wire N__22216;
    wire N__22215;
    wire N__22212;
    wire N__22209;
    wire N__22206;
    wire N__22203;
    wire N__22200;
    wire N__22199;
    wire N__22190;
    wire N__22187;
    wire N__22186;
    wire N__22183;
    wire N__22180;
    wire N__22179;
    wire N__22178;
    wire N__22175;
    wire N__22174;
    wire N__22173;
    wire N__22172;
    wire N__22169;
    wire N__22166;
    wire N__22163;
    wire N__22160;
    wire N__22155;
    wire N__22152;
    wire N__22149;
    wire N__22146;
    wire N__22143;
    wire N__22140;
    wire N__22137;
    wire N__22134;
    wire N__22129;
    wire N__22126;
    wire N__22125;
    wire N__22124;
    wire N__22123;
    wire N__22122;
    wire N__22119;
    wire N__22116;
    wire N__22107;
    wire N__22104;
    wire N__22097;
    wire N__22092;
    wire N__22089;
    wire N__22086;
    wire N__22083;
    wire N__22080;
    wire N__22077;
    wire N__22074;
    wire N__22069;
    wire N__22066;
    wire N__22057;
    wire N__22052;
    wire N__22045;
    wire N__22030;
    wire N__22027;
    wire N__22024;
    wire N__22021;
    wire N__22018;
    wire N__22015;
    wire N__22012;
    wire N__22009;
    wire N__22006;
    wire N__22003;
    wire N__22000;
    wire N__21997;
    wire N__21994;
    wire N__21991;
    wire N__21990;
    wire N__21989;
    wire N__21986;
    wire N__21983;
    wire N__21980;
    wire N__21979;
    wire N__21976;
    wire N__21973;
    wire N__21970;
    wire N__21967;
    wire N__21962;
    wire N__21957;
    wire N__21956;
    wire N__21951;
    wire N__21948;
    wire N__21947;
    wire N__21946;
    wire N__21943;
    wire N__21940;
    wire N__21937;
    wire N__21934;
    wire N__21933;
    wire N__21926;
    wire N__21923;
    wire N__21920;
    wire N__21917;
    wire N__21914;
    wire N__21911;
    wire N__21904;
    wire N__21901;
    wire N__21898;
    wire N__21895;
    wire N__21892;
    wire N__21889;
    wire N__21886;
    wire N__21883;
    wire N__21880;
    wire N__21877;
    wire N__21874;
    wire N__21871;
    wire N__21868;
    wire N__21865;
    wire N__21862;
    wire N__21859;
    wire N__21856;
    wire N__21853;
    wire N__21850;
    wire N__21847;
    wire N__21844;
    wire N__21841;
    wire N__21838;
    wire N__21835;
    wire N__21832;
    wire N__21829;
    wire N__21826;
    wire N__21823;
    wire N__21820;
    wire N__21817;
    wire N__21814;
    wire N__21811;
    wire N__21808;
    wire N__21805;
    wire N__21802;
    wire N__21799;
    wire N__21796;
    wire N__21793;
    wire N__21790;
    wire N__21787;
    wire N__21784;
    wire N__21781;
    wire N__21778;
    wire N__21775;
    wire N__21772;
    wire N__21769;
    wire N__21766;
    wire N__21763;
    wire N__21760;
    wire N__21757;
    wire N__21754;
    wire N__21751;
    wire N__21748;
    wire N__21745;
    wire N__21742;
    wire N__21739;
    wire N__21736;
    wire N__21733;
    wire N__21730;
    wire N__21727;
    wire N__21724;
    wire N__21721;
    wire N__21718;
    wire N__21715;
    wire N__21712;
    wire N__21709;
    wire N__21706;
    wire N__21703;
    wire N__21700;
    wire N__21697;
    wire N__21694;
    wire N__21693;
    wire N__21692;
    wire N__21691;
    wire N__21688;
    wire N__21685;
    wire N__21684;
    wire N__21683;
    wire N__21682;
    wire N__21679;
    wire N__21676;
    wire N__21675;
    wire N__21674;
    wire N__21671;
    wire N__21668;
    wire N__21665;
    wire N__21662;
    wire N__21661;
    wire N__21658;
    wire N__21653;
    wire N__21652;
    wire N__21649;
    wire N__21646;
    wire N__21645;
    wire N__21644;
    wire N__21641;
    wire N__21636;
    wire N__21633;
    wire N__21628;
    wire N__21625;
    wire N__21622;
    wire N__21617;
    wire N__21614;
    wire N__21611;
    wire N__21606;
    wire N__21603;
    wire N__21594;
    wire N__21591;
    wire N__21580;
    wire N__21577;
    wire N__21574;
    wire N__21571;
    wire N__21568;
    wire N__21565;
    wire N__21562;
    wire N__21559;
    wire N__21558;
    wire N__21555;
    wire N__21552;
    wire N__21549;
    wire N__21546;
    wire N__21545;
    wire N__21542;
    wire N__21539;
    wire N__21536;
    wire N__21533;
    wire N__21530;
    wire N__21527;
    wire N__21522;
    wire N__21519;
    wire N__21516;
    wire N__21513;
    wire N__21510;
    wire N__21507;
    wire N__21502;
    wire N__21499;
    wire N__21496;
    wire N__21493;
    wire N__21490;
    wire N__21489;
    wire N__21488;
    wire N__21485;
    wire N__21484;
    wire N__21483;
    wire N__21482;
    wire N__21479;
    wire N__21478;
    wire N__21475;
    wire N__21474;
    wire N__21471;
    wire N__21468;
    wire N__21465;
    wire N__21462;
    wire N__21461;
    wire N__21460;
    wire N__21459;
    wire N__21458;
    wire N__21457;
    wire N__21454;
    wire N__21453;
    wire N__21450;
    wire N__21449;
    wire N__21446;
    wire N__21443;
    wire N__21438;
    wire N__21433;
    wire N__21430;
    wire N__21427;
    wire N__21424;
    wire N__21421;
    wire N__21418;
    wire N__21415;
    wire N__21412;
    wire N__21409;
    wire N__21406;
    wire N__21403;
    wire N__21400;
    wire N__21393;
    wire N__21390;
    wire N__21387;
    wire N__21382;
    wire N__21377;
    wire N__21368;
    wire N__21359;
    wire N__21352;
    wire N__21351;
    wire N__21350;
    wire N__21349;
    wire N__21348;
    wire N__21347;
    wire N__21344;
    wire N__21341;
    wire N__21338;
    wire N__21335;
    wire N__21332;
    wire N__21331;
    wire N__21330;
    wire N__21329;
    wire N__21326;
    wire N__21325;
    wire N__21324;
    wire N__21321;
    wire N__21320;
    wire N__21319;
    wire N__21318;
    wire N__21315;
    wire N__21308;
    wire N__21305;
    wire N__21304;
    wire N__21303;
    wire N__21302;
    wire N__21301;
    wire N__21300;
    wire N__21297;
    wire N__21294;
    wire N__21291;
    wire N__21288;
    wire N__21285;
    wire N__21284;
    wire N__21283;
    wire N__21282;
    wire N__21281;
    wire N__21280;
    wire N__21277;
    wire N__21276;
    wire N__21275;
    wire N__21272;
    wire N__21269;
    wire N__21268;
    wire N__21267;
    wire N__21266;
    wire N__21265;
    wire N__21262;
    wire N__21261;
    wire N__21260;
    wire N__21259;
    wire N__21258;
    wire N__21251;
    wire N__21248;
    wire N__21245;
    wire N__21242;
    wire N__21239;
    wire N__21236;
    wire N__21235;
    wire N__21234;
    wire N__21233;
    wire N__21230;
    wire N__21221;
    wire N__21218;
    wire N__21215;
    wire N__21212;
    wire N__21209;
    wire N__21206;
    wire N__21205;
    wire N__21202;
    wire N__21199;
    wire N__21196;
    wire N__21195;
    wire N__21192;
    wire N__21189;
    wire N__21186;
    wire N__21185;
    wire N__21182;
    wire N__21179;
    wire N__21178;
    wire N__21175;
    wire N__21172;
    wire N__21171;
    wire N__21168;
    wire N__21167;
    wire N__21166;
    wire N__21163;
    wire N__21160;
    wire N__21157;
    wire N__21152;
    wire N__21145;
    wire N__21142;
    wire N__21139;
    wire N__21138;
    wire N__21135;
    wire N__21132;
    wire N__21131;
    wire N__21124;
    wire N__21121;
    wire N__21120;
    wire N__21119;
    wire N__21118;
    wire N__21117;
    wire N__21114;
    wire N__21111;
    wire N__21108;
    wire N__21105;
    wire N__21102;
    wire N__21097;
    wire N__21094;
    wire N__21089;
    wire N__21086;
    wire N__21083;
    wire N__21080;
    wire N__21077;
    wire N__21072;
    wire N__21069;
    wire N__21066;
    wire N__21063;
    wire N__21060;
    wire N__21059;
    wire N__21056;
    wire N__21055;
    wire N__21054;
    wire N__21053;
    wire N__21052;
    wire N__21051;
    wire N__21050;
    wire N__21049;
    wire N__21048;
    wire N__21045;
    wire N__21040;
    wire N__21037;
    wire N__21030;
    wire N__21027;
    wire N__21020;
    wire N__21017;
    wire N__21014;
    wire N__21009;
    wire N__21006;
    wire N__21005;
    wire N__21004;
    wire N__21003;
    wire N__21002;
    wire N__20999;
    wire N__20992;
    wire N__20989;
    wire N__20982;
    wire N__20977;
    wire N__20974;
    wire N__20969;
    wire N__20966;
    wire N__20963;
    wire N__20960;
    wire N__20957;
    wire N__20952;
    wire N__20945;
    wire N__20942;
    wire N__20937;
    wire N__20934;
    wire N__20931;
    wire N__20928;
    wire N__20925;
    wire N__20918;
    wire N__20915;
    wire N__20908;
    wire N__20903;
    wire N__20898;
    wire N__20893;
    wire N__20886;
    wire N__20873;
    wire N__20864;
    wire N__20833;
    wire N__20830;
    wire N__20827;
    wire N__20824;
    wire N__20821;
    wire N__20818;
    wire N__20815;
    wire N__20812;
    wire N__20809;
    wire N__20806;
    wire N__20803;
    wire N__20800;
    wire N__20797;
    wire N__20794;
    wire N__20791;
    wire N__20788;
    wire N__20785;
    wire N__20782;
    wire N__20779;
    wire N__20776;
    wire N__20773;
    wire N__20770;
    wire N__20767;
    wire N__20764;
    wire N__20761;
    wire N__20758;
    wire N__20755;
    wire N__20752;
    wire N__20749;
    wire N__20746;
    wire N__20743;
    wire N__20740;
    wire N__20737;
    wire N__20734;
    wire N__20731;
    wire N__20728;
    wire N__20725;
    wire N__20722;
    wire N__20719;
    wire N__20716;
    wire N__20713;
    wire N__20710;
    wire N__20707;
    wire N__20704;
    wire N__20701;
    wire N__20698;
    wire N__20697;
    wire N__20696;
    wire N__20695;
    wire N__20694;
    wire N__20693;
    wire N__20680;
    wire N__20679;
    wire N__20678;
    wire N__20675;
    wire N__20674;
    wire N__20673;
    wire N__20672;
    wire N__20669;
    wire N__20666;
    wire N__20663;
    wire N__20658;
    wire N__20655;
    wire N__20652;
    wire N__20647;
    wire N__20644;
    wire N__20637;
    wire N__20636;
    wire N__20635;
    wire N__20634;
    wire N__20633;
    wire N__20632;
    wire N__20631;
    wire N__20630;
    wire N__20629;
    wire N__20628;
    wire N__20625;
    wire N__20622;
    wire N__20617;
    wire N__20614;
    wire N__20611;
    wire N__20608;
    wire N__20599;
    wire N__20584;
    wire N__20581;
    wire N__20578;
    wire N__20575;
    wire N__20572;
    wire N__20569;
    wire N__20568;
    wire N__20567;
    wire N__20566;
    wire N__20565;
    wire N__20564;
    wire N__20561;
    wire N__20558;
    wire N__20557;
    wire N__20554;
    wire N__20551;
    wire N__20546;
    wire N__20537;
    wire N__20536;
    wire N__20535;
    wire N__20534;
    wire N__20531;
    wire N__20528;
    wire N__20525;
    wire N__20522;
    wire N__20521;
    wire N__20518;
    wire N__20515;
    wire N__20512;
    wire N__20507;
    wire N__20504;
    wire N__20503;
    wire N__20498;
    wire N__20495;
    wire N__20492;
    wire N__20487;
    wire N__20484;
    wire N__20483;
    wire N__20480;
    wire N__20477;
    wire N__20472;
    wire N__20469;
    wire N__20466;
    wire N__20465;
    wire N__20464;
    wire N__20463;
    wire N__20462;
    wire N__20459;
    wire N__20456;
    wire N__20449;
    wire N__20446;
    wire N__20439;
    wire N__20436;
    wire N__20427;
    wire N__20422;
    wire N__20421;
    wire N__20418;
    wire N__20415;
    wire N__20412;
    wire N__20409;
    wire N__20406;
    wire N__20403;
    wire N__20400;
    wire N__20397;
    wire N__20394;
    wire N__20391;
    wire N__20388;
    wire N__20385;
    wire N__20382;
    wire N__20379;
    wire N__20376;
    wire N__20373;
    wire N__20370;
    wire N__20367;
    wire N__20364;
    wire N__20361;
    wire N__20358;
    wire N__20355;
    wire N__20352;
    wire N__20349;
    wire N__20346;
    wire N__20343;
    wire N__20340;
    wire N__20337;
    wire N__20334;
    wire N__20331;
    wire N__20328;
    wire N__20325;
    wire N__20322;
    wire N__20319;
    wire N__20316;
    wire N__20313;
    wire N__20310;
    wire N__20307;
    wire N__20304;
    wire N__20301;
    wire N__20298;
    wire N__20295;
    wire N__20292;
    wire N__20289;
    wire N__20286;
    wire N__20283;
    wire N__20280;
    wire N__20277;
    wire N__20274;
    wire N__20271;
    wire N__20268;
    wire N__20265;
    wire N__20262;
    wire N__20259;
    wire N__20256;
    wire N__20253;
    wire N__20250;
    wire N__20247;
    wire N__20244;
    wire N__20241;
    wire N__20240;
    wire N__20237;
    wire N__20234;
    wire N__20231;
    wire N__20228;
    wire N__20225;
    wire N__20222;
    wire N__20219;
    wire N__20216;
    wire N__20213;
    wire N__20210;
    wire N__20209;
    wire N__20206;
    wire N__20203;
    wire N__20200;
    wire N__20197;
    wire N__20194;
    wire N__20189;
    wire N__20182;
    wire N__20179;
    wire N__20178;
    wire N__20177;
    wire N__20176;
    wire N__20175;
    wire N__20174;
    wire N__20173;
    wire N__20172;
    wire N__20171;
    wire N__20170;
    wire N__20167;
    wire N__20166;
    wire N__20165;
    wire N__20164;
    wire N__20163;
    wire N__20162;
    wire N__20161;
    wire N__20160;
    wire N__20159;
    wire N__20158;
    wire N__20157;
    wire N__20156;
    wire N__20155;
    wire N__20154;
    wire N__20153;
    wire N__20152;
    wire N__20151;
    wire N__20150;
    wire N__20149;
    wire N__20148;
    wire N__20147;
    wire N__20146;
    wire N__20145;
    wire N__20144;
    wire N__20143;
    wire N__20142;
    wire N__20141;
    wire N__20140;
    wire N__20139;
    wire N__20138;
    wire N__20137;
    wire N__20136;
    wire N__20135;
    wire N__20134;
    wire N__20133;
    wire N__20132;
    wire N__20131;
    wire N__20130;
    wire N__20129;
    wire N__20128;
    wire N__20029;
    wire N__20026;
    wire N__20023;
    wire N__20020;
    wire N__20017;
    wire N__20014;
    wire N__20011;
    wire N__20008;
    wire N__20005;
    wire N__20002;
    wire N__19999;
    wire N__19996;
    wire N__19993;
    wire N__19990;
    wire N__19987;
    wire N__19984;
    wire N__19981;
    wire N__19978;
    wire N__19975;
    wire N__19972;
    wire N__19969;
    wire N__19966;
    wire N__19963;
    wire N__19960;
    wire N__19957;
    wire N__19954;
    wire N__19951;
    wire N__19948;
    wire N__19945;
    wire N__19942;
    wire N__19939;
    wire N__19936;
    wire N__19933;
    wire N__19930;
    wire N__19927;
    wire N__19924;
    wire N__19921;
    wire N__19918;
    wire N__19915;
    wire N__19912;
    wire N__19909;
    wire N__19906;
    wire N__19905;
    wire N__19902;
    wire N__19899;
    wire N__19898;
    wire N__19895;
    wire N__19892;
    wire N__19889;
    wire N__19886;
    wire N__19883;
    wire N__19880;
    wire N__19877;
    wire N__19874;
    wire N__19871;
    wire N__19866;
    wire N__19863;
    wire N__19860;
    wire N__19855;
    wire N__19852;
    wire N__19851;
    wire N__19850;
    wire N__19847;
    wire N__19844;
    wire N__19843;
    wire N__19840;
    wire N__19839;
    wire N__19838;
    wire N__19833;
    wire N__19830;
    wire N__19829;
    wire N__19826;
    wire N__19823;
    wire N__19820;
    wire N__19819;
    wire N__19818;
    wire N__19813;
    wire N__19810;
    wire N__19809;
    wire N__19808;
    wire N__19807;
    wire N__19802;
    wire N__19799;
    wire N__19796;
    wire N__19793;
    wire N__19792;
    wire N__19791;
    wire N__19786;
    wire N__19783;
    wire N__19780;
    wire N__19777;
    wire N__19776;
    wire N__19769;
    wire N__19766;
    wire N__19763;
    wire N__19760;
    wire N__19759;
    wire N__19758;
    wire N__19757;
    wire N__19752;
    wire N__19747;
    wire N__19744;
    wire N__19743;
    wire N__19742;
    wire N__19739;
    wire N__19734;
    wire N__19731;
    wire N__19728;
    wire N__19725;
    wire N__19724;
    wire N__19723;
    wire N__19720;
    wire N__19719;
    wire N__19718;
    wire N__19715;
    wire N__19712;
    wire N__19709;
    wire N__19706;
    wire N__19705;
    wire N__19704;
    wire N__19701;
    wire N__19700;
    wire N__19699;
    wire N__19690;
    wire N__19687;
    wire N__19684;
    wire N__19681;
    wire N__19680;
    wire N__19677;
    wire N__19674;
    wire N__19671;
    wire N__19668;
    wire N__19661;
    wire N__19658;
    wire N__19657;
    wire N__19656;
    wire N__19653;
    wire N__19652;
    wire N__19649;
    wire N__19646;
    wire N__19643;
    wire N__19636;
    wire N__19633;
    wire N__19630;
    wire N__19629;
    wire N__19622;
    wire N__19615;
    wire N__19612;
    wire N__19609;
    wire N__19606;
    wire N__19603;
    wire N__19602;
    wire N__19595;
    wire N__19588;
    wire N__19585;
    wire N__19580;
    wire N__19575;
    wire N__19572;
    wire N__19569;
    wire N__19566;
    wire N__19563;
    wire N__19558;
    wire N__19555;
    wire N__19552;
    wire N__19547;
    wire N__19544;
    wire N__19539;
    wire N__19534;
    wire N__19529;
    wire N__19526;
    wire N__19519;
    wire N__19516;
    wire N__19513;
    wire N__19510;
    wire N__19507;
    wire N__19504;
    wire N__19501;
    wire N__19498;
    wire N__19495;
    wire N__19492;
    wire N__19489;
    wire N__19486;
    wire N__19483;
    wire N__19480;
    wire N__19477;
    wire N__19474;
    wire N__19471;
    wire N__19468;
    wire N__19465;
    wire N__19462;
    wire N__19459;
    wire N__19456;
    wire N__19453;
    wire N__19450;
    wire N__19447;
    wire N__19444;
    wire N__19441;
    wire N__19438;
    wire N__19435;
    wire N__19432;
    wire N__19429;
    wire N__19426;
    wire N__19423;
    wire N__19420;
    wire N__19417;
    wire N__19414;
    wire N__19411;
    wire N__19408;
    wire N__19405;
    wire N__19402;
    wire N__19399;
    wire N__19396;
    wire N__19393;
    wire N__19390;
    wire N__19387;
    wire N__19384;
    wire N__19381;
    wire N__19378;
    wire N__19375;
    wire N__19372;
    wire N__19369;
    wire N__19366;
    wire N__19363;
    wire N__19360;
    wire N__19357;
    wire N__19354;
    wire N__19351;
    wire N__19348;
    wire N__19345;
    wire N__19342;
    wire N__19339;
    wire N__19338;
    wire N__19337;
    wire N__19334;
    wire N__19329;
    wire N__19324;
    wire N__19321;
    wire N__19320;
    wire N__19319;
    wire N__19316;
    wire N__19311;
    wire N__19306;
    wire N__19303;
    wire N__19302;
    wire N__19301;
    wire N__19298;
    wire N__19293;
    wire N__19288;
    wire N__19285;
    wire N__19284;
    wire N__19283;
    wire N__19280;
    wire N__19275;
    wire N__19270;
    wire N__19267;
    wire N__19266;
    wire N__19263;
    wire N__19260;
    wire N__19255;
    wire N__19252;
    wire N__19249;
    wire N__19248;
    wire N__19245;
    wire N__19242;
    wire N__19239;
    wire N__19234;
    wire N__19233;
    wire N__19230;
    wire N__19227;
    wire N__19224;
    wire N__19221;
    wire N__19218;
    wire N__19213;
    wire N__19210;
    wire N__19207;
    wire N__19204;
    wire N__19201;
    wire N__19198;
    wire N__19195;
    wire N__19192;
    wire N__19189;
    wire N__19186;
    wire N__19183;
    wire N__19180;
    wire N__19177;
    wire N__19174;
    wire N__19171;
    wire N__19168;
    wire N__19165;
    wire N__19162;
    wire N__19159;
    wire N__19156;
    wire N__19153;
    wire N__19150;
    wire N__19147;
    wire N__19144;
    wire N__19141;
    wire N__19138;
    wire N__19135;
    wire N__19132;
    wire N__19129;
    wire N__19126;
    wire N__19123;
    wire N__19120;
    wire N__19117;
    wire N__19114;
    wire N__19113;
    wire N__19110;
    wire N__19109;
    wire N__19106;
    wire N__19103;
    wire N__19100;
    wire N__19099;
    wire N__19098;
    wire N__19097;
    wire N__19094;
    wire N__19093;
    wire N__19090;
    wire N__19087;
    wire N__19086;
    wire N__19083;
    wire N__19082;
    wire N__19081;
    wire N__19080;
    wire N__19079;
    wire N__19078;
    wire N__19077;
    wire N__19072;
    wire N__19069;
    wire N__19068;
    wire N__19067;
    wire N__19066;
    wire N__19065;
    wire N__19064;
    wire N__19061;
    wire N__19060;
    wire N__19059;
    wire N__19054;
    wire N__19051;
    wire N__19048;
    wire N__19043;
    wire N__19034;
    wire N__19031;
    wire N__19028;
    wire N__19025;
    wire N__19024;
    wire N__19023;
    wire N__19022;
    wire N__19019;
    wire N__19014;
    wire N__19011;
    wire N__19008;
    wire N__19003;
    wire N__18998;
    wire N__18993;
    wire N__18990;
    wire N__18989;
    wire N__18988;
    wire N__18987;
    wire N__18982;
    wire N__18979;
    wire N__18976;
    wire N__18971;
    wire N__18966;
    wire N__18957;
    wire N__18954;
    wire N__18951;
    wire N__18948;
    wire N__18943;
    wire N__18940;
    wire N__18929;
    wire N__18916;
    wire N__18913;
    wire N__18912;
    wire N__18909;
    wire N__18906;
    wire N__18903;
    wire N__18898;
    wire N__18895;
    wire N__18892;
    wire N__18889;
    wire N__18886;
    wire N__18885;
    wire N__18882;
    wire N__18879;
    wire N__18876;
    wire N__18873;
    wire N__18870;
    wire N__18867;
    wire N__18864;
    wire N__18861;
    wire N__18858;
    wire N__18855;
    wire N__18852;
    wire N__18849;
    wire N__18846;
    wire N__18843;
    wire N__18840;
    wire N__18837;
    wire N__18834;
    wire N__18831;
    wire N__18828;
    wire N__18825;
    wire N__18822;
    wire N__18819;
    wire N__18816;
    wire N__18813;
    wire N__18810;
    wire N__18807;
    wire N__18804;
    wire N__18801;
    wire N__18798;
    wire N__18795;
    wire N__18792;
    wire N__18789;
    wire N__18786;
    wire N__18783;
    wire N__18780;
    wire N__18777;
    wire N__18774;
    wire N__18771;
    wire N__18768;
    wire N__18765;
    wire N__18762;
    wire N__18759;
    wire N__18756;
    wire N__18753;
    wire N__18750;
    wire N__18747;
    wire N__18744;
    wire N__18741;
    wire N__18738;
    wire N__18735;
    wire N__18732;
    wire N__18729;
    wire N__18726;
    wire N__18723;
    wire N__18720;
    wire N__18717;
    wire N__18714;
    wire N__18711;
    wire N__18708;
    wire N__18705;
    wire N__18702;
    wire N__18699;
    wire N__18696;
    wire N__18693;
    wire N__18690;
    wire N__18687;
    wire N__18684;
    wire N__18681;
    wire N__18678;
    wire N__18675;
    wire N__18672;
    wire N__18669;
    wire N__18664;
    wire N__18661;
    wire N__18658;
    wire N__18655;
    wire N__18652;
    wire N__18651;
    wire N__18646;
    wire N__18645;
    wire N__18642;
    wire N__18639;
    wire N__18636;
    wire N__18633;
    wire N__18628;
    wire N__18625;
    wire N__18622;
    wire N__18619;
    wire N__18616;
    wire N__18613;
    wire N__18610;
    wire N__18607;
    wire N__18604;
    wire N__18601;
    wire N__18598;
    wire N__18595;
    wire N__18594;
    wire N__18593;
    wire N__18590;
    wire N__18585;
    wire N__18580;
    wire N__18577;
    wire N__18574;
    wire N__18571;
    wire N__18568;
    wire N__18567;
    wire N__18564;
    wire N__18561;
    wire N__18556;
    wire N__18553;
    wire N__18550;
    wire N__18549;
    wire N__18546;
    wire N__18543;
    wire N__18538;
    wire N__18535;
    wire N__18534;
    wire N__18531;
    wire N__18528;
    wire N__18525;
    wire N__18522;
    wire N__18519;
    wire N__18516;
    wire N__18513;
    wire N__18510;
    wire N__18507;
    wire N__18504;
    wire N__18501;
    wire N__18498;
    wire N__18495;
    wire N__18492;
    wire N__18489;
    wire N__18486;
    wire N__18483;
    wire N__18480;
    wire N__18477;
    wire N__18474;
    wire N__18471;
    wire N__18468;
    wire N__18465;
    wire N__18462;
    wire N__18459;
    wire N__18456;
    wire N__18453;
    wire N__18450;
    wire N__18447;
    wire N__18444;
    wire N__18441;
    wire N__18438;
    wire N__18435;
    wire N__18432;
    wire N__18429;
    wire N__18426;
    wire N__18423;
    wire N__18420;
    wire N__18417;
    wire N__18414;
    wire N__18411;
    wire N__18408;
    wire N__18405;
    wire N__18402;
    wire N__18399;
    wire N__18396;
    wire N__18393;
    wire N__18390;
    wire N__18387;
    wire N__18384;
    wire N__18381;
    wire N__18378;
    wire N__18375;
    wire N__18372;
    wire N__18369;
    wire N__18366;
    wire N__18363;
    wire N__18360;
    wire N__18357;
    wire N__18354;
    wire N__18351;
    wire N__18348;
    wire N__18345;
    wire N__18342;
    wire N__18339;
    wire N__18336;
    wire N__18333;
    wire N__18330;
    wire N__18327;
    wire N__18324;
    wire N__18319;
    wire N__18316;
    wire N__18315;
    wire N__18314;
    wire N__18311;
    wire N__18308;
    wire N__18307;
    wire N__18304;
    wire N__18303;
    wire N__18302;
    wire N__18301;
    wire N__18300;
    wire N__18299;
    wire N__18298;
    wire N__18295;
    wire N__18294;
    wire N__18291;
    wire N__18288;
    wire N__18285;
    wire N__18280;
    wire N__18275;
    wire N__18274;
    wire N__18273;
    wire N__18270;
    wire N__18269;
    wire N__18266;
    wire N__18263;
    wire N__18260;
    wire N__18257;
    wire N__18250;
    wire N__18247;
    wire N__18242;
    wire N__18237;
    wire N__18220;
    wire N__18217;
    wire N__18214;
    wire N__18211;
    wire N__18208;
    wire N__18205;
    wire N__18202;
    wire N__18199;
    wire N__18196;
    wire N__18193;
    wire N__18192;
    wire N__18189;
    wire N__18186;
    wire N__18183;
    wire N__18180;
    wire N__18177;
    wire N__18174;
    wire N__18171;
    wire N__18168;
    wire N__18165;
    wire N__18162;
    wire N__18159;
    wire N__18156;
    wire N__18153;
    wire N__18150;
    wire N__18147;
    wire N__18144;
    wire N__18141;
    wire N__18138;
    wire N__18135;
    wire N__18132;
    wire N__18129;
    wire N__18126;
    wire N__18123;
    wire N__18120;
    wire N__18117;
    wire N__18114;
    wire N__18111;
    wire N__18108;
    wire N__18105;
    wire N__18102;
    wire N__18099;
    wire N__18096;
    wire N__18093;
    wire N__18090;
    wire N__18087;
    wire N__18084;
    wire N__18081;
    wire N__18078;
    wire N__18075;
    wire N__18072;
    wire N__18069;
    wire N__18066;
    wire N__18063;
    wire N__18060;
    wire N__18057;
    wire N__18054;
    wire N__18051;
    wire N__18048;
    wire N__18045;
    wire N__18042;
    wire N__18039;
    wire N__18036;
    wire N__18033;
    wire N__18030;
    wire N__18027;
    wire N__18024;
    wire N__18021;
    wire N__18018;
    wire N__18015;
    wire N__18012;
    wire N__18009;
    wire N__18006;
    wire N__18003;
    wire N__18000;
    wire N__17997;
    wire N__17994;
    wire N__17991;
    wire N__17988;
    wire N__17983;
    wire N__17980;
    wire N__17979;
    wire N__17976;
    wire N__17973;
    wire N__17972;
    wire N__17969;
    wire N__17966;
    wire N__17963;
    wire N__17956;
    wire N__17955;
    wire N__17952;
    wire N__17949;
    wire N__17944;
    wire N__17941;
    wire N__17938;
    wire N__17937;
    wire N__17934;
    wire N__17933;
    wire N__17930;
    wire N__17929;
    wire N__17928;
    wire N__17927;
    wire N__17924;
    wire N__17921;
    wire N__17918;
    wire N__17915;
    wire N__17912;
    wire N__17909;
    wire N__17908;
    wire N__17907;
    wire N__17906;
    wire N__17905;
    wire N__17900;
    wire N__17897;
    wire N__17894;
    wire N__17891;
    wire N__17888;
    wire N__17885;
    wire N__17884;
    wire N__17883;
    wire N__17882;
    wire N__17881;
    wire N__17878;
    wire N__17875;
    wire N__17872;
    wire N__17863;
    wire N__17858;
    wire N__17855;
    wire N__17852;
    wire N__17849;
    wire N__17846;
    wire N__17827;
    wire N__17824;
    wire N__17821;
    wire N__17820;
    wire N__17817;
    wire N__17814;
    wire N__17809;
    wire N__17808;
    wire N__17807;
    wire N__17800;
    wire N__17797;
    wire N__17796;
    wire N__17793;
    wire N__17790;
    wire N__17785;
    wire N__17782;
    wire N__17779;
    wire N__17778;
    wire N__17775;
    wire N__17774;
    wire N__17771;
    wire N__17770;
    wire N__17767;
    wire N__17766;
    wire N__17763;
    wire N__17762;
    wire N__17759;
    wire N__17756;
    wire N__17753;
    wire N__17750;
    wire N__17747;
    wire N__17744;
    wire N__17743;
    wire N__17738;
    wire N__17733;
    wire N__17728;
    wire N__17725;
    wire N__17720;
    wire N__17717;
    wire N__17714;
    wire N__17707;
    wire N__17704;
    wire N__17701;
    wire N__17698;
    wire N__17697;
    wire N__17694;
    wire N__17693;
    wire N__17690;
    wire N__17687;
    wire N__17684;
    wire N__17681;
    wire N__17678;
    wire N__17675;
    wire N__17672;
    wire N__17669;
    wire N__17666;
    wire N__17663;
    wire N__17660;
    wire N__17657;
    wire N__17654;
    wire N__17651;
    wire N__17646;
    wire N__17643;
    wire N__17638;
    wire N__17635;
    wire N__17632;
    wire N__17629;
    wire N__17628;
    wire N__17625;
    wire N__17624;
    wire N__17621;
    wire N__17618;
    wire N__17615;
    wire N__17612;
    wire N__17609;
    wire N__17606;
    wire N__17601;
    wire N__17598;
    wire N__17595;
    wire N__17592;
    wire N__17589;
    wire N__17586;
    wire N__17581;
    wire N__17578;
    wire N__17575;
    wire N__17572;
    wire N__17569;
    wire N__17566;
    wire N__17563;
    wire N__17560;
    wire N__17557;
    wire N__17554;
    wire N__17551;
    wire N__17548;
    wire N__17545;
    wire N__17542;
    wire N__17539;
    wire N__17536;
    wire N__17533;
    wire N__17530;
    wire N__17527;
    wire N__17524;
    wire N__17521;
    wire N__17518;
    wire N__17515;
    wire N__17512;
    wire N__17509;
    wire N__17506;
    wire N__17503;
    wire N__17500;
    wire N__17497;
    wire N__17494;
    wire N__17491;
    wire N__17488;
    wire N__17485;
    wire N__17482;
    wire N__17479;
    wire N__17476;
    wire N__17473;
    wire N__17470;
    wire N__17467;
    wire N__17464;
    wire N__17461;
    wire N__17458;
    wire N__17455;
    wire N__17452;
    wire N__17449;
    wire N__17446;
    wire N__17443;
    wire N__17440;
    wire N__17437;
    wire N__17434;
    wire N__17431;
    wire N__17428;
    wire N__17425;
    wire N__17422;
    wire N__17419;
    wire N__17416;
    wire N__17413;
    wire N__17410;
    wire N__17407;
    wire N__17404;
    wire N__17401;
    wire N__17398;
    wire N__17395;
    wire N__17392;
    wire N__17389;
    wire N__17386;
    wire N__17383;
    wire N__17380;
    wire N__17377;
    wire N__17374;
    wire N__17371;
    wire N__17368;
    wire N__17365;
    wire N__17362;
    wire N__17359;
    wire N__17356;
    wire N__17353;
    wire N__17352;
    wire N__17351;
    wire N__17350;
    wire N__17347;
    wire N__17342;
    wire N__17337;
    wire N__17332;
    wire N__17331;
    wire N__17330;
    wire N__17329;
    wire N__17326;
    wire N__17323;
    wire N__17320;
    wire N__17315;
    wire N__17308;
    wire N__17305;
    wire N__17302;
    wire N__17299;
    wire N__17296;
    wire N__17293;
    wire N__17292;
    wire N__17287;
    wire N__17284;
    wire N__17283;
    wire N__17280;
    wire N__17277;
    wire N__17274;
    wire N__17271;
    wire N__17268;
    wire N__17265;
    wire N__17262;
    wire N__17259;
    wire N__17256;
    wire N__17253;
    wire N__17250;
    wire N__17247;
    wire N__17244;
    wire N__17241;
    wire N__17238;
    wire N__17235;
    wire N__17232;
    wire N__17229;
    wire N__17226;
    wire N__17223;
    wire N__17220;
    wire N__17217;
    wire N__17214;
    wire N__17211;
    wire N__17208;
    wire N__17205;
    wire N__17202;
    wire N__17199;
    wire N__17196;
    wire N__17193;
    wire N__17190;
    wire N__17187;
    wire N__17184;
    wire N__17181;
    wire N__17178;
    wire N__17175;
    wire N__17172;
    wire N__17169;
    wire N__17166;
    wire N__17163;
    wire N__17160;
    wire N__17157;
    wire N__17154;
    wire N__17151;
    wire N__17148;
    wire N__17145;
    wire N__17142;
    wire N__17139;
    wire N__17136;
    wire N__17133;
    wire N__17130;
    wire N__17127;
    wire N__17124;
    wire N__17121;
    wire N__17118;
    wire N__17115;
    wire N__17112;
    wire N__17109;
    wire N__17106;
    wire N__17103;
    wire N__17100;
    wire N__17097;
    wire N__17094;
    wire N__17091;
    wire N__17088;
    wire N__17085;
    wire N__17082;
    wire N__17079;
    wire N__17076;
    wire N__17073;
    wire N__17070;
    wire N__17067;
    wire N__17064;
    wire N__17061;
    wire N__17058;
    wire N__17053;
    wire N__17050;
    wire N__17047;
    wire N__17044;
    wire N__17041;
    wire N__17040;
    wire N__17037;
    wire N__17034;
    wire N__17033;
    wire N__17028;
    wire N__17025;
    wire N__17024;
    wire N__17019;
    wire N__17016;
    wire N__17013;
    wire N__17010;
    wire N__17007;
    wire N__17004;
    wire N__17001;
    wire N__16998;
    wire N__16995;
    wire N__16992;
    wire N__16987;
    wire N__16986;
    wire N__16983;
    wire N__16980;
    wire N__16977;
    wire N__16976;
    wire N__16973;
    wire N__16972;
    wire N__16969;
    wire N__16966;
    wire N__16963;
    wire N__16960;
    wire N__16957;
    wire N__16954;
    wire N__16949;
    wire N__16942;
    wire N__16939;
    wire N__16936;
    wire N__16935;
    wire N__16932;
    wire N__16929;
    wire N__16928;
    wire N__16925;
    wire N__16922;
    wire N__16919;
    wire N__16912;
    wire N__16909;
    wire N__16908;
    wire N__16905;
    wire N__16902;
    wire N__16897;
    wire N__16894;
    wire N__16891;
    wire N__16888;
    wire N__16885;
    wire N__16882;
    wire N__16879;
    wire N__16876;
    wire N__16873;
    wire N__16870;
    wire N__16867;
    wire N__16864;
    wire N__16863;
    wire N__16862;
    wire N__16859;
    wire N__16858;
    wire N__16855;
    wire N__16852;
    wire N__16849;
    wire N__16846;
    wire N__16843;
    wire N__16834;
    wire N__16831;
    wire N__16828;
    wire N__16825;
    wire N__16824;
    wire N__16821;
    wire N__16818;
    wire N__16817;
    wire N__16812;
    wire N__16809;
    wire N__16808;
    wire N__16803;
    wire N__16800;
    wire N__16795;
    wire N__16792;
    wire N__16789;
    wire N__16786;
    wire N__16785;
    wire N__16784;
    wire N__16783;
    wire N__16782;
    wire N__16781;
    wire N__16780;
    wire N__16779;
    wire N__16776;
    wire N__16773;
    wire N__16772;
    wire N__16769;
    wire N__16762;
    wire N__16757;
    wire N__16750;
    wire N__16741;
    wire N__16740;
    wire N__16739;
    wire N__16738;
    wire N__16737;
    wire N__16736;
    wire N__16735;
    wire N__16732;
    wire N__16729;
    wire N__16726;
    wire N__16725;
    wire N__16724;
    wire N__16721;
    wire N__16718;
    wire N__16711;
    wire N__16708;
    wire N__16705;
    wire N__16698;
    wire N__16687;
    wire N__16686;
    wire N__16685;
    wire N__16682;
    wire N__16679;
    wire N__16678;
    wire N__16677;
    wire N__16676;
    wire N__16675;
    wire N__16674;
    wire N__16673;
    wire N__16670;
    wire N__16665;
    wire N__16662;
    wire N__16657;
    wire N__16650;
    wire N__16639;
    wire N__16638;
    wire N__16635;
    wire N__16634;
    wire N__16631;
    wire N__16628;
    wire N__16625;
    wire N__16624;
    wire N__16621;
    wire N__16618;
    wire N__16615;
    wire N__16612;
    wire N__16609;
    wire N__16604;
    wire N__16601;
    wire N__16598;
    wire N__16595;
    wire N__16592;
    wire N__16587;
    wire N__16584;
    wire N__16581;
    wire N__16578;
    wire N__16573;
    wire N__16570;
    wire N__16567;
    wire N__16564;
    wire N__16561;
    wire N__16558;
    wire N__16555;
    wire N__16552;
    wire N__16549;
    wire N__16546;
    wire N__16543;
    wire N__16540;
    wire N__16537;
    wire N__16534;
    wire N__16531;
    wire N__16528;
    wire N__16525;
    wire N__16522;
    wire N__16519;
    wire N__16516;
    wire N__16513;
    wire N__16510;
    wire N__16507;
    wire N__16504;
    wire N__16501;
    wire N__16498;
    wire N__16495;
    wire N__16492;
    wire N__16491;
    wire N__16490;
    wire N__16487;
    wire N__16484;
    wire N__16483;
    wire N__16480;
    wire N__16475;
    wire N__16472;
    wire N__16469;
    wire N__16464;
    wire N__16461;
    wire N__16458;
    wire N__16455;
    wire N__16452;
    wire N__16447;
    wire N__16446;
    wire N__16443;
    wire N__16440;
    wire N__16439;
    wire N__16438;
    wire N__16433;
    wire N__16430;
    wire N__16427;
    wire N__16420;
    wire N__16417;
    wire N__16414;
    wire N__16411;
    wire N__16408;
    wire N__16405;
    wire N__16404;
    wire N__16401;
    wire N__16398;
    wire N__16397;
    wire N__16396;
    wire N__16391;
    wire N__16388;
    wire N__16385;
    wire N__16380;
    wire N__16377;
    wire N__16374;
    wire N__16371;
    wire N__16368;
    wire N__16365;
    wire N__16362;
    wire N__16357;
    wire N__16356;
    wire N__16353;
    wire N__16350;
    wire N__16345;
    wire N__16342;
    wire N__16341;
    wire N__16338;
    wire N__16335;
    wire N__16330;
    wire N__16327;
    wire N__16326;
    wire N__16323;
    wire N__16320;
    wire N__16315;
    wire N__16312;
    wire N__16311;
    wire N__16308;
    wire N__16305;
    wire N__16300;
    wire N__16297;
    wire N__16296;
    wire N__16293;
    wire N__16290;
    wire N__16285;
    wire N__16282;
    wire N__16279;
    wire N__16278;
    wire N__16275;
    wire N__16272;
    wire N__16267;
    wire N__16266;
    wire N__16263;
    wire N__16260;
    wire N__16257;
    wire N__16254;
    wire N__16251;
    wire N__16248;
    wire N__16243;
    wire N__16240;
    wire N__16237;
    wire N__16234;
    wire N__16231;
    wire N__16228;
    wire N__16225;
    wire N__16222;
    wire N__16219;
    wire N__16216;
    wire N__16215;
    wire N__16212;
    wire N__16209;
    wire N__16206;
    wire N__16203;
    wire N__16200;
    wire N__16197;
    wire N__16194;
    wire N__16191;
    wire N__16188;
    wire N__16185;
    wire N__16182;
    wire N__16179;
    wire N__16176;
    wire N__16173;
    wire N__16170;
    wire N__16167;
    wire N__16164;
    wire N__16161;
    wire N__16158;
    wire N__16155;
    wire N__16152;
    wire N__16149;
    wire N__16146;
    wire N__16143;
    wire N__16140;
    wire N__16137;
    wire N__16134;
    wire N__16131;
    wire N__16128;
    wire N__16125;
    wire N__16122;
    wire N__16119;
    wire N__16116;
    wire N__16113;
    wire N__16110;
    wire N__16107;
    wire N__16104;
    wire N__16101;
    wire N__16098;
    wire N__16095;
    wire N__16092;
    wire N__16089;
    wire N__16086;
    wire N__16083;
    wire N__16080;
    wire N__16077;
    wire N__16074;
    wire N__16071;
    wire N__16068;
    wire N__16065;
    wire N__16062;
    wire N__16059;
    wire N__16056;
    wire N__16053;
    wire N__16050;
    wire N__16047;
    wire N__16044;
    wire N__16041;
    wire N__16038;
    wire N__16035;
    wire N__16032;
    wire N__16029;
    wire N__16026;
    wire N__16023;
    wire N__16020;
    wire N__16017;
    wire N__16014;
    wire N__16011;
    wire N__16010;
    wire N__16007;
    wire N__16004;
    wire N__16001;
    wire N__15998;
    wire N__15995;
    wire N__15994;
    wire N__15991;
    wire N__15986;
    wire N__15983;
    wire N__15978;
    wire N__15973;
    wire N__15970;
    wire N__15967;
    wire N__15964;
    wire N__15961;
    wire N__15958;
    wire N__15957;
    wire N__15954;
    wire N__15951;
    wire N__15948;
    wire N__15945;
    wire N__15942;
    wire N__15939;
    wire N__15936;
    wire N__15933;
    wire N__15930;
    wire N__15927;
    wire N__15924;
    wire N__15921;
    wire N__15918;
    wire N__15915;
    wire N__15912;
    wire N__15909;
    wire N__15906;
    wire N__15903;
    wire N__15900;
    wire N__15897;
    wire N__15894;
    wire N__15891;
    wire N__15888;
    wire N__15885;
    wire N__15882;
    wire N__15879;
    wire N__15876;
    wire N__15873;
    wire N__15870;
    wire N__15867;
    wire N__15864;
    wire N__15861;
    wire N__15858;
    wire N__15855;
    wire N__15852;
    wire N__15849;
    wire N__15846;
    wire N__15843;
    wire N__15840;
    wire N__15837;
    wire N__15834;
    wire N__15831;
    wire N__15828;
    wire N__15825;
    wire N__15822;
    wire N__15819;
    wire N__15816;
    wire N__15813;
    wire N__15810;
    wire N__15807;
    wire N__15804;
    wire N__15801;
    wire N__15798;
    wire N__15795;
    wire N__15792;
    wire N__15789;
    wire N__15786;
    wire N__15783;
    wire N__15780;
    wire N__15777;
    wire N__15774;
    wire N__15771;
    wire N__15768;
    wire N__15765;
    wire N__15762;
    wire N__15759;
    wire N__15758;
    wire N__15755;
    wire N__15752;
    wire N__15751;
    wire N__15748;
    wire N__15745;
    wire N__15742;
    wire N__15739;
    wire N__15736;
    wire N__15733;
    wire N__15730;
    wire N__15725;
    wire N__15720;
    wire N__15715;
    wire N__15712;
    wire N__15709;
    wire N__15706;
    wire N__15703;
    wire N__15700;
    wire N__15697;
    wire N__15694;
    wire N__15691;
    wire N__15688;
    wire N__15685;
    wire N__15682;
    wire N__15679;
    wire N__15676;
    wire N__15673;
    wire N__15670;
    wire N__15667;
    wire N__15664;
    wire N__15661;
    wire N__15658;
    wire N__15657;
    wire N__15654;
    wire N__15651;
    wire N__15648;
    wire N__15645;
    wire N__15642;
    wire N__15639;
    wire N__15636;
    wire N__15633;
    wire N__15630;
    wire N__15627;
    wire N__15624;
    wire N__15621;
    wire N__15618;
    wire N__15615;
    wire N__15612;
    wire N__15609;
    wire N__15606;
    wire N__15603;
    wire N__15600;
    wire N__15597;
    wire N__15594;
    wire N__15591;
    wire N__15588;
    wire N__15585;
    wire N__15582;
    wire N__15579;
    wire N__15576;
    wire N__15573;
    wire N__15570;
    wire N__15567;
    wire N__15564;
    wire N__15561;
    wire N__15558;
    wire N__15555;
    wire N__15552;
    wire N__15549;
    wire N__15546;
    wire N__15543;
    wire N__15540;
    wire N__15537;
    wire N__15534;
    wire N__15531;
    wire N__15528;
    wire N__15525;
    wire N__15522;
    wire N__15519;
    wire N__15516;
    wire N__15513;
    wire N__15510;
    wire N__15507;
    wire N__15504;
    wire N__15501;
    wire N__15498;
    wire N__15495;
    wire N__15492;
    wire N__15489;
    wire N__15486;
    wire N__15483;
    wire N__15480;
    wire N__15479;
    wire N__15476;
    wire N__15473;
    wire N__15470;
    wire N__15467;
    wire N__15464;
    wire N__15461;
    wire N__15458;
    wire N__15455;
    wire N__15452;
    wire N__15449;
    wire N__15446;
    wire N__15443;
    wire N__15442;
    wire N__15439;
    wire N__15436;
    wire N__15433;
    wire N__15430;
    wire N__15427;
    wire N__15424;
    wire N__15415;
    wire N__15412;
    wire N__15409;
    wire N__15406;
    wire N__15403;
    wire N__15400;
    wire N__15399;
    wire N__15396;
    wire N__15393;
    wire N__15390;
    wire N__15387;
    wire N__15384;
    wire N__15381;
    wire N__15378;
    wire N__15375;
    wire N__15372;
    wire N__15369;
    wire N__15366;
    wire N__15363;
    wire N__15360;
    wire N__15357;
    wire N__15354;
    wire N__15351;
    wire N__15348;
    wire N__15345;
    wire N__15342;
    wire N__15339;
    wire N__15336;
    wire N__15333;
    wire N__15330;
    wire N__15327;
    wire N__15324;
    wire N__15321;
    wire N__15318;
    wire N__15315;
    wire N__15312;
    wire N__15309;
    wire N__15306;
    wire N__15303;
    wire N__15300;
    wire N__15297;
    wire N__15294;
    wire N__15291;
    wire N__15288;
    wire N__15285;
    wire N__15282;
    wire N__15279;
    wire N__15276;
    wire N__15273;
    wire N__15270;
    wire N__15267;
    wire N__15264;
    wire N__15261;
    wire N__15258;
    wire N__15255;
    wire N__15252;
    wire N__15249;
    wire N__15246;
    wire N__15243;
    wire N__15240;
    wire N__15237;
    wire N__15234;
    wire N__15231;
    wire N__15228;
    wire N__15225;
    wire N__15222;
    wire N__15219;
    wire N__15218;
    wire N__15215;
    wire N__15212;
    wire N__15209;
    wire N__15206;
    wire N__15203;
    wire N__15202;
    wire N__15199;
    wire N__15196;
    wire N__15193;
    wire N__15190;
    wire N__15183;
    wire N__15178;
    wire N__15175;
    wire N__15172;
    wire N__15169;
    wire N__15166;
    wire N__15163;
    wire N__15162;
    wire N__15159;
    wire N__15156;
    wire N__15153;
    wire N__15150;
    wire N__15147;
    wire N__15144;
    wire N__15141;
    wire N__15138;
    wire N__15135;
    wire N__15132;
    wire N__15129;
    wire N__15126;
    wire N__15123;
    wire N__15120;
    wire N__15117;
    wire N__15114;
    wire N__15111;
    wire N__15108;
    wire N__15105;
    wire N__15102;
    wire N__15099;
    wire N__15096;
    wire N__15093;
    wire N__15090;
    wire N__15087;
    wire N__15084;
    wire N__15081;
    wire N__15078;
    wire N__15075;
    wire N__15072;
    wire N__15069;
    wire N__15066;
    wire N__15063;
    wire N__15060;
    wire N__15057;
    wire N__15054;
    wire N__15051;
    wire N__15048;
    wire N__15045;
    wire N__15042;
    wire N__15039;
    wire N__15036;
    wire N__15033;
    wire N__15030;
    wire N__15027;
    wire N__15024;
    wire N__15021;
    wire N__15018;
    wire N__15015;
    wire N__15012;
    wire N__15009;
    wire N__15006;
    wire N__15003;
    wire N__15000;
    wire N__14997;
    wire N__14994;
    wire N__14991;
    wire N__14990;
    wire N__14987;
    wire N__14984;
    wire N__14981;
    wire N__14978;
    wire N__14975;
    wire N__14972;
    wire N__14969;
    wire N__14966;
    wire N__14963;
    wire N__14960;
    wire N__14957;
    wire N__14956;
    wire N__14953;
    wire N__14950;
    wire N__14947;
    wire N__14944;
    wire N__14941;
    wire N__14938;
    wire N__14935;
    wire N__14932;
    wire N__14929;
    wire N__14926;
    wire N__14923;
    wire N__14914;
    wire N__14911;
    wire N__14908;
    wire N__14905;
    wire N__14902;
    wire N__14899;
    wire N__14896;
    wire N__14895;
    wire N__14892;
    wire N__14889;
    wire N__14886;
    wire N__14883;
    wire N__14880;
    wire N__14877;
    wire N__14874;
    wire N__14871;
    wire N__14868;
    wire N__14865;
    wire N__14862;
    wire N__14859;
    wire N__14856;
    wire N__14853;
    wire N__14850;
    wire N__14847;
    wire N__14844;
    wire N__14841;
    wire N__14838;
    wire N__14835;
    wire N__14832;
    wire N__14829;
    wire N__14826;
    wire N__14823;
    wire N__14820;
    wire N__14817;
    wire N__14814;
    wire N__14811;
    wire N__14808;
    wire N__14805;
    wire N__14802;
    wire N__14799;
    wire N__14796;
    wire N__14793;
    wire N__14790;
    wire N__14787;
    wire N__14784;
    wire N__14781;
    wire N__14778;
    wire N__14775;
    wire N__14772;
    wire N__14769;
    wire N__14766;
    wire N__14763;
    wire N__14760;
    wire N__14757;
    wire N__14754;
    wire N__14751;
    wire N__14748;
    wire N__14745;
    wire N__14742;
    wire N__14739;
    wire N__14736;
    wire N__14733;
    wire N__14730;
    wire N__14727;
    wire N__14724;
    wire N__14721;
    wire N__14718;
    wire N__14715;
    wire N__14714;
    wire N__14711;
    wire N__14708;
    wire N__14705;
    wire N__14702;
    wire N__14699;
    wire N__14696;
    wire N__14693;
    wire N__14690;
    wire N__14687;
    wire N__14686;
    wire N__14683;
    wire N__14680;
    wire N__14677;
    wire N__14674;
    wire N__14669;
    wire N__14662;
    wire N__14659;
    wire N__14656;
    wire N__14653;
    wire N__14650;
    wire N__14647;
    wire N__14646;
    wire N__14643;
    wire N__14640;
    wire N__14637;
    wire N__14634;
    wire N__14631;
    wire N__14628;
    wire N__14625;
    wire N__14622;
    wire N__14619;
    wire N__14616;
    wire N__14613;
    wire N__14610;
    wire N__14607;
    wire N__14604;
    wire N__14601;
    wire N__14598;
    wire N__14595;
    wire N__14592;
    wire N__14589;
    wire N__14586;
    wire N__14583;
    wire N__14580;
    wire N__14577;
    wire N__14574;
    wire N__14571;
    wire N__14568;
    wire N__14565;
    wire N__14562;
    wire N__14559;
    wire N__14556;
    wire N__14553;
    wire N__14550;
    wire N__14547;
    wire N__14544;
    wire N__14541;
    wire N__14538;
    wire N__14535;
    wire N__14532;
    wire N__14529;
    wire N__14526;
    wire N__14523;
    wire N__14520;
    wire N__14517;
    wire N__14514;
    wire N__14511;
    wire N__14508;
    wire N__14505;
    wire N__14502;
    wire N__14499;
    wire N__14496;
    wire N__14493;
    wire N__14490;
    wire N__14487;
    wire N__14484;
    wire N__14481;
    wire N__14478;
    wire N__14475;
    wire N__14472;
    wire N__14469;
    wire N__14466;
    wire N__14463;
    wire N__14462;
    wire N__14459;
    wire N__14456;
    wire N__14453;
    wire N__14450;
    wire N__14447;
    wire N__14446;
    wire N__14443;
    wire N__14440;
    wire N__14437;
    wire N__14434;
    wire N__14431;
    wire N__14428;
    wire N__14425;
    wire N__14422;
    wire N__14419;
    wire N__14414;
    wire N__14407;
    wire N__14404;
    wire N__14401;
    wire N__14398;
    wire N__14395;
    wire N__14392;
    wire N__14391;
    wire N__14388;
    wire N__14385;
    wire N__14382;
    wire N__14379;
    wire N__14376;
    wire N__14373;
    wire N__14370;
    wire N__14367;
    wire N__14364;
    wire N__14361;
    wire N__14358;
    wire N__14355;
    wire N__14352;
    wire N__14349;
    wire N__14346;
    wire N__14343;
    wire N__14340;
    wire N__14337;
    wire N__14334;
    wire N__14331;
    wire N__14328;
    wire N__14325;
    wire N__14322;
    wire N__14319;
    wire N__14316;
    wire N__14313;
    wire N__14310;
    wire N__14307;
    wire N__14304;
    wire N__14301;
    wire N__14298;
    wire N__14295;
    wire N__14292;
    wire N__14289;
    wire N__14286;
    wire N__14283;
    wire N__14280;
    wire N__14277;
    wire N__14274;
    wire N__14271;
    wire N__14268;
    wire N__14265;
    wire N__14262;
    wire N__14259;
    wire N__14256;
    wire N__14253;
    wire N__14250;
    wire N__14247;
    wire N__14244;
    wire N__14241;
    wire N__14238;
    wire N__14235;
    wire N__14232;
    wire N__14229;
    wire N__14226;
    wire N__14223;
    wire N__14220;
    wire N__14217;
    wire N__14214;
    wire N__14211;
    wire N__14210;
    wire N__14207;
    wire N__14204;
    wire N__14201;
    wire N__14198;
    wire N__14195;
    wire N__14192;
    wire N__14189;
    wire N__14186;
    wire N__14183;
    wire N__14182;
    wire N__14179;
    wire N__14176;
    wire N__14173;
    wire N__14170;
    wire N__14165;
    wire N__14158;
    wire N__14155;
    wire N__14152;
    wire N__14149;
    wire N__14146;
    wire N__14143;
    wire N__14140;
    wire N__14139;
    wire N__14136;
    wire N__14133;
    wire N__14130;
    wire N__14127;
    wire N__14124;
    wire N__14121;
    wire N__14118;
    wire N__14115;
    wire N__14112;
    wire N__14109;
    wire N__14106;
    wire N__14103;
    wire N__14100;
    wire N__14097;
    wire N__14094;
    wire N__14091;
    wire N__14088;
    wire N__14085;
    wire N__14082;
    wire N__14079;
    wire N__14076;
    wire N__14073;
    wire N__14070;
    wire N__14067;
    wire N__14064;
    wire N__14061;
    wire N__14058;
    wire N__14055;
    wire N__14052;
    wire N__14049;
    wire N__14046;
    wire N__14043;
    wire N__14040;
    wire N__14037;
    wire N__14034;
    wire N__14031;
    wire N__14028;
    wire N__14025;
    wire N__14022;
    wire N__14019;
    wire N__14016;
    wire N__14013;
    wire N__14010;
    wire N__14007;
    wire N__14004;
    wire N__14001;
    wire N__13998;
    wire N__13995;
    wire N__13992;
    wire N__13989;
    wire N__13986;
    wire N__13983;
    wire N__13980;
    wire N__13977;
    wire N__13976;
    wire N__13973;
    wire N__13970;
    wire N__13967;
    wire N__13964;
    wire N__13961;
    wire N__13958;
    wire N__13955;
    wire N__13952;
    wire N__13949;
    wire N__13946;
    wire N__13943;
    wire N__13942;
    wire N__13939;
    wire N__13936;
    wire N__13933;
    wire N__13930;
    wire N__13927;
    wire N__13924;
    wire N__13921;
    wire N__13918;
    wire N__13915;
    wire N__13912;
    wire N__13909;
    wire N__13900;
    wire N__13897;
    wire N__13894;
    wire N__13891;
    wire N__13888;
    wire N__13885;
    wire N__13882;
    wire N__13879;
    wire N__13876;
    wire N__13873;
    wire N__13870;
    wire N__13867;
    wire N__13864;
    wire N__13861;
    wire N__13858;
    wire N__13855;
    wire N__13852;
    wire N__13849;
    wire N__13846;
    wire N__13843;
    wire N__13842;
    wire N__13839;
    wire N__13836;
    wire N__13833;
    wire N__13830;
    wire N__13827;
    wire N__13822;
    wire N__13819;
    wire N__13816;
    wire N__13813;
    wire N__13810;
    wire N__13807;
    wire N__13804;
    wire N__13801;
    wire N__13798;
    wire N__13795;
    wire N__13792;
    wire N__13789;
    wire N__13786;
    wire N__13783;
    wire N__13782;
    wire N__13779;
    wire N__13776;
    wire N__13773;
    wire N__13770;
    wire N__13767;
    wire N__13764;
    wire N__13761;
    wire N__13758;
    wire N__13755;
    wire N__13752;
    wire N__13749;
    wire N__13746;
    wire N__13743;
    wire N__13740;
    wire N__13737;
    wire N__13734;
    wire N__13731;
    wire N__13728;
    wire N__13725;
    wire N__13722;
    wire N__13719;
    wire N__13716;
    wire N__13713;
    wire N__13710;
    wire N__13707;
    wire N__13704;
    wire N__13701;
    wire N__13698;
    wire N__13695;
    wire N__13692;
    wire N__13689;
    wire N__13686;
    wire N__13683;
    wire N__13680;
    wire N__13677;
    wire N__13674;
    wire N__13671;
    wire N__13668;
    wire N__13665;
    wire N__13662;
    wire N__13659;
    wire N__13656;
    wire N__13653;
    wire N__13650;
    wire N__13647;
    wire N__13644;
    wire N__13641;
    wire N__13638;
    wire N__13635;
    wire N__13632;
    wire N__13629;
    wire N__13626;
    wire N__13623;
    wire N__13620;
    wire N__13617;
    wire N__13614;
    wire N__13611;
    wire N__13608;
    wire N__13605;
    wire N__13602;
    wire N__13599;
    wire N__13596;
    wire N__13593;
    wire N__13590;
    wire N__13589;
    wire N__13586;
    wire N__13583;
    wire N__13580;
    wire N__13577;
    wire N__13574;
    wire N__13571;
    wire N__13570;
    wire N__13567;
    wire N__13564;
    wire N__13561;
    wire N__13558;
    wire N__13553;
    wire N__13546;
    wire N__13545;
    wire N__13544;
    wire N__13543;
    wire N__13540;
    wire N__13537;
    wire N__13534;
    wire N__13531;
    wire N__13528;
    wire N__13525;
    wire N__13522;
    wire N__13513;
    wire N__13510;
    wire N__13507;
    wire N__13504;
    wire N__13501;
    wire N__13498;
    wire N__13497;
    wire N__13496;
    wire N__13495;
    wire N__13492;
    wire N__13487;
    wire N__13484;
    wire N__13477;
    wire N__13474;
    wire N__13471;
    wire N__13468;
    wire N__13465;
    wire N__13462;
    wire N__13459;
    wire N__13456;
    wire N__13455;
    wire N__13454;
    wire N__13451;
    wire N__13448;
    wire N__13445;
    wire N__13440;
    wire N__13439;
    wire N__13434;
    wire N__13431;
    wire N__13426;
    wire N__13423;
    wire N__13422;
    wire N__13419;
    wire N__13416;
    wire N__13413;
    wire N__13410;
    wire N__13407;
    wire N__13404;
    wire N__13399;
    wire N__13396;
    wire N__13393;
    wire N__13390;
    wire N__13389;
    wire N__13386;
    wire N__13385;
    wire N__13384;
    wire N__13381;
    wire N__13378;
    wire N__13373;
    wire N__13370;
    wire N__13363;
    wire N__13360;
    wire N__13357;
    wire N__13354;
    wire N__13351;
    wire N__13348;
    wire N__13345;
    wire N__13342;
    wire N__13339;
    wire N__13338;
    wire N__13337;
    wire N__13336;
    wire N__13333;
    wire N__13330;
    wire N__13327;
    wire N__13324;
    wire N__13315;
    wire N__13312;
    wire N__13309;
    wire N__13306;
    wire N__13305;
    wire N__13304;
    wire N__13301;
    wire N__13298;
    wire N__13297;
    wire N__13294;
    wire N__13289;
    wire N__13286;
    wire N__13283;
    wire N__13276;
    wire N__13273;
    wire N__13270;
    wire N__13267;
    wire N__13266;
    wire N__13265;
    wire N__13262;
    wire N__13259;
    wire N__13258;
    wire N__13255;
    wire N__13252;
    wire N__13249;
    wire N__13246;
    wire N__13243;
    wire N__13234;
    wire N__13231;
    wire N__13228;
    wire N__13225;
    wire N__13222;
    wire N__13219;
    wire N__13216;
    wire N__13213;
    wire N__13210;
    wire N__13207;
    wire N__13204;
    wire N__13201;
    wire N__13198;
    wire N__13195;
    wire N__13192;
    wire N__13189;
    wire N__13186;
    wire N__13183;
    wire N__13180;
    wire N__13177;
    wire N__13174;
    wire N__13171;
    wire N__13168;
    wire N__13165;
    wire N__13164;
    wire N__13161;
    wire N__13160;
    wire N__13159;
    wire N__13156;
    wire N__13153;
    wire N__13148;
    wire N__13141;
    wire N__13140;
    wire N__13137;
    wire N__13134;
    wire N__13129;
    wire N__13126;
    wire N__13123;
    wire N__13122;
    wire N__13121;
    wire N__13120;
    wire N__13117;
    wire N__13114;
    wire N__13109;
    wire N__13102;
    wire N__13099;
    wire N__13096;
    wire N__13093;
    wire N__13092;
    wire N__13089;
    wire N__13086;
    wire N__13083;
    wire N__13080;
    wire N__13075;
    wire N__13072;
    wire N__13069;
    wire N__13066;
    wire N__13063;
    wire N__13060;
    wire N__13057;
    wire N__13054;
    wire N__13053;
    wire N__13050;
    wire N__13047;
    wire N__13044;
    wire N__13041;
    wire N__13038;
    wire N__13033;
    wire N__13030;
    wire N__13027;
    wire N__13024;
    wire N__13021;
    wire N__13018;
    wire N__13015;
    wire N__13014;
    wire N__13011;
    wire N__13008;
    wire N__13005;
    wire N__13002;
    wire N__12999;
    wire N__12996;
    wire N__12993;
    wire N__12990;
    wire N__12987;
    wire N__12984;
    wire N__12981;
    wire N__12978;
    wire N__12975;
    wire N__12972;
    wire N__12969;
    wire N__12966;
    wire N__12963;
    wire N__12960;
    wire N__12957;
    wire N__12954;
    wire N__12951;
    wire N__12948;
    wire N__12945;
    wire N__12942;
    wire N__12939;
    wire N__12936;
    wire N__12933;
    wire N__12930;
    wire N__12927;
    wire N__12924;
    wire N__12921;
    wire N__12918;
    wire N__12915;
    wire N__12912;
    wire N__12909;
    wire N__12906;
    wire N__12903;
    wire N__12900;
    wire N__12897;
    wire N__12894;
    wire N__12891;
    wire N__12888;
    wire N__12885;
    wire N__12882;
    wire N__12879;
    wire N__12876;
    wire N__12873;
    wire N__12870;
    wire N__12867;
    wire N__12864;
    wire N__12861;
    wire N__12858;
    wire N__12855;
    wire N__12852;
    wire N__12849;
    wire N__12846;
    wire N__12843;
    wire N__12840;
    wire N__12837;
    wire N__12834;
    wire N__12831;
    wire N__12828;
    wire N__12825;
    wire N__12822;
    wire N__12819;
    wire N__12816;
    wire N__12813;
    wire N__12810;
    wire N__12805;
    wire N__12802;
    wire N__12801;
    wire N__12798;
    wire N__12795;
    wire N__12792;
    wire N__12789;
    wire N__12786;
    wire N__12781;
    wire N__12778;
    wire N__12777;
    wire N__12774;
    wire N__12771;
    wire N__12768;
    wire N__12763;
    wire N__12762;
    wire N__12759;
    wire N__12756;
    wire N__12753;
    wire N__12750;
    wire N__12747;
    wire N__12744;
    wire N__12741;
    wire N__12738;
    wire N__12735;
    wire N__12732;
    wire N__12729;
    wire N__12726;
    wire N__12723;
    wire N__12720;
    wire N__12717;
    wire N__12714;
    wire N__12711;
    wire N__12708;
    wire N__12705;
    wire N__12702;
    wire N__12699;
    wire N__12696;
    wire N__12693;
    wire N__12690;
    wire N__12687;
    wire N__12684;
    wire N__12681;
    wire N__12678;
    wire N__12675;
    wire N__12672;
    wire N__12669;
    wire N__12666;
    wire N__12663;
    wire N__12660;
    wire N__12657;
    wire N__12654;
    wire N__12651;
    wire N__12648;
    wire N__12645;
    wire N__12642;
    wire N__12639;
    wire N__12636;
    wire N__12633;
    wire N__12630;
    wire N__12627;
    wire N__12624;
    wire N__12621;
    wire N__12618;
    wire N__12615;
    wire N__12612;
    wire N__12609;
    wire N__12606;
    wire N__12603;
    wire N__12600;
    wire N__12597;
    wire N__12594;
    wire N__12591;
    wire N__12588;
    wire N__12585;
    wire N__12582;
    wire N__12579;
    wire N__12576;
    wire N__12573;
    wire N__12570;
    wire N__12567;
    wire N__12564;
    wire N__12561;
    wire N__12558;
    wire N__12553;
    wire N__12550;
    wire N__12547;
    wire N__12544;
    wire N__12543;
    wire N__12540;
    wire N__12537;
    wire N__12532;
    wire N__12529;
    wire N__12526;
    wire N__12523;
    wire N__12520;
    wire N__12517;
    wire N__12514;
    wire N__12513;
    wire N__12508;
    wire N__12505;
    wire N__12502;
    wire N__12499;
    wire N__12496;
    wire N__12495;
    wire N__12492;
    wire N__12489;
    wire N__12486;
    wire N__12481;
    wire N__12478;
    wire N__12475;
    wire N__12472;
    wire N__12469;
    wire N__12468;
    wire N__12465;
    wire N__12462;
    wire N__12459;
    wire N__12456;
    wire N__12453;
    wire N__12450;
    wire N__12447;
    wire N__12444;
    wire N__12441;
    wire N__12438;
    wire N__12435;
    wire N__12432;
    wire N__12429;
    wire N__12426;
    wire N__12423;
    wire N__12420;
    wire N__12417;
    wire N__12414;
    wire N__12411;
    wire N__12408;
    wire N__12405;
    wire N__12402;
    wire N__12399;
    wire N__12396;
    wire N__12393;
    wire N__12390;
    wire N__12387;
    wire N__12384;
    wire N__12381;
    wire N__12378;
    wire N__12375;
    wire N__12372;
    wire N__12369;
    wire N__12366;
    wire N__12363;
    wire N__12360;
    wire N__12357;
    wire N__12354;
    wire N__12351;
    wire N__12348;
    wire N__12345;
    wire N__12342;
    wire N__12339;
    wire N__12336;
    wire N__12333;
    wire N__12330;
    wire N__12327;
    wire N__12324;
    wire N__12321;
    wire N__12318;
    wire N__12315;
    wire N__12312;
    wire N__12309;
    wire N__12306;
    wire N__12303;
    wire N__12300;
    wire N__12297;
    wire N__12294;
    wire N__12291;
    wire N__12288;
    wire N__12285;
    wire N__12282;
    wire N__12279;
    wire N__12276;
    wire N__12273;
    wire N__12270;
    wire N__12267;
    wire N__12264;
    wire N__12261;
    wire N__12258;
    wire N__12255;
    wire N__12252;
    wire N__12247;
    wire N__12244;
    wire N__12241;
    wire N__12238;
    wire N__12235;
    wire N__12232;
    wire N__12229;
    wire N__12226;
    wire N__12223;
    wire N__12220;
    wire N__12219;
    wire N__12216;
    wire N__12215;
    wire N__12212;
    wire N__12209;
    wire N__12206;
    wire N__12203;
    wire N__12200;
    wire N__12197;
    wire N__12194;
    wire N__12191;
    wire N__12188;
    wire N__12185;
    wire N__12180;
    wire N__12177;
    wire N__12172;
    wire N__12169;
    wire N__12168;
    wire N__12167;
    wire N__12164;
    wire N__12161;
    wire N__12158;
    wire N__12155;
    wire N__12152;
    wire N__12149;
    wire N__12146;
    wire N__12143;
    wire N__12140;
    wire N__12137;
    wire N__12134;
    wire N__12131;
    wire N__12126;
    wire N__12121;
    wire N__12118;
    wire N__12115;
    wire N__12112;
    wire N__12109;
    wire N__12106;
    wire N__12103;
    wire N__12100;
    wire N__12097;
    wire N__12094;
    wire N__12091;
    wire N__12088;
    wire N__12085;
    wire N__12082;
    wire N__12079;
    wire N__12078;
    wire N__12075;
    wire N__12072;
    wire N__12069;
    wire N__12066;
    wire N__12063;
    wire N__12060;
    wire N__12057;
    wire N__12052;
    wire N__12051;
    wire N__12048;
    wire N__12045;
    wire N__12042;
    wire N__12039;
    wire N__12036;
    wire N__12031;
    wire N__12028;
    wire N__12027;
    wire N__12024;
    wire N__12021;
    wire N__12018;
    wire N__12015;
    wire N__12012;
    wire N__12009;
    wire N__12006;
    wire N__12003;
    wire N__12000;
    wire N__11997;
    wire N__11994;
    wire N__11991;
    wire N__11988;
    wire N__11985;
    wire N__11982;
    wire N__11979;
    wire N__11976;
    wire N__11973;
    wire N__11970;
    wire N__11967;
    wire N__11964;
    wire N__11961;
    wire N__11958;
    wire N__11955;
    wire N__11952;
    wire N__11949;
    wire N__11946;
    wire N__11943;
    wire N__11940;
    wire N__11937;
    wire N__11934;
    wire N__11931;
    wire N__11928;
    wire N__11925;
    wire N__11922;
    wire N__11919;
    wire N__11916;
    wire N__11913;
    wire N__11910;
    wire N__11907;
    wire N__11904;
    wire N__11901;
    wire N__11898;
    wire N__11895;
    wire N__11892;
    wire N__11889;
    wire N__11886;
    wire N__11883;
    wire N__11880;
    wire N__11877;
    wire N__11874;
    wire N__11871;
    wire N__11868;
    wire N__11865;
    wire N__11862;
    wire N__11859;
    wire N__11856;
    wire N__11853;
    wire N__11850;
    wire N__11847;
    wire N__11844;
    wire N__11841;
    wire N__11838;
    wire N__11835;
    wire N__11832;
    wire N__11829;
    wire N__11826;
    wire N__11823;
    wire N__11820;
    wire N__11817;
    wire N__11812;
    wire N__11809;
    wire N__11806;
    wire N__11803;
    wire N__11802;
    wire N__11799;
    wire N__11796;
    wire N__11793;
    wire N__11788;
    wire N__11785;
    wire N__11784;
    wire N__11781;
    wire N__11778;
    wire N__11775;
    wire N__11772;
    wire N__11769;
    wire N__11766;
    wire N__11763;
    wire N__11760;
    wire N__11757;
    wire N__11754;
    wire N__11751;
    wire N__11748;
    wire N__11745;
    wire N__11742;
    wire N__11739;
    wire N__11736;
    wire N__11733;
    wire N__11730;
    wire N__11727;
    wire N__11724;
    wire N__11721;
    wire N__11718;
    wire N__11715;
    wire N__11712;
    wire N__11709;
    wire N__11706;
    wire N__11703;
    wire N__11700;
    wire N__11697;
    wire N__11694;
    wire N__11691;
    wire N__11688;
    wire N__11685;
    wire N__11682;
    wire N__11679;
    wire N__11676;
    wire N__11673;
    wire N__11670;
    wire N__11667;
    wire N__11664;
    wire N__11661;
    wire N__11658;
    wire N__11655;
    wire N__11652;
    wire N__11649;
    wire N__11646;
    wire N__11643;
    wire N__11640;
    wire N__11637;
    wire N__11634;
    wire N__11631;
    wire N__11628;
    wire N__11625;
    wire N__11622;
    wire N__11619;
    wire N__11616;
    wire N__11613;
    wire N__11610;
    wire N__11607;
    wire N__11604;
    wire N__11601;
    wire N__11598;
    wire N__11595;
    wire N__11592;
    wire N__11589;
    wire N__11586;
    wire N__11583;
    wire N__11580;
    wire N__11577;
    wire N__11574;
    wire N__11571;
    wire N__11568;
    wire N__11565;
    wire N__11562;
    wire N__11557;
    wire N__11554;
    wire N__11551;
    wire N__11548;
    wire N__11545;
    wire N__11542;
    wire N__11539;
    wire N__11536;
    wire N__11533;
    wire N__11530;
    wire N__11527;
    wire N__11524;
    wire N__11521;
    wire N__11518;
    wire N__11515;
    wire N__11512;
    wire N__11509;
    wire N__11506;
    wire N__11503;
    wire N__11500;
    wire N__11497;
    wire N__11494;
    wire N__11491;
    wire N__11488;
    wire N__11485;
    wire N__11482;
    wire N__11479;
    wire N__11476;
    wire N__11473;
    wire N__11470;
    wire N__11467;
    wire N__11464;
    wire N__11461;
    wire N__11458;
    wire N__11455;
    wire N__11452;
    wire N__11449;
    wire N__11446;
    wire N__11443;
    wire N__11440;
    wire N__11437;
    wire N__11434;
    wire N__11431;
    wire N__11428;
    wire N__11425;
    wire N__11422;
    wire N__11419;
    wire N__11416;
    wire N__11415;
    wire N__11414;
    wire N__11411;
    wire N__11408;
    wire N__11405;
    wire N__11398;
    wire N__11395;
    wire N__11392;
    wire N__11391;
    wire N__11388;
    wire N__11385;
    wire N__11380;
    wire N__11379;
    wire N__11378;
    wire N__11377;
    wire N__11374;
    wire N__11369;
    wire N__11366;
    wire N__11361;
    wire N__11356;
    wire N__11353;
    wire N__11352;
    wire N__11349;
    wire N__11348;
    wire N__11345;
    wire N__11344;
    wire N__11341;
    wire N__11338;
    wire N__11333;
    wire N__11326;
    wire N__11323;
    wire N__11320;
    wire N__11317;
    wire N__11314;
    wire N__11311;
    wire N__11308;
    wire N__11305;
    wire N__11302;
    wire N__11299;
    wire N__11296;
    wire N__11295;
    wire N__11292;
    wire N__11289;
    wire N__11284;
    wire N__11283;
    wire N__11282;
    wire N__11281;
    wire N__11278;
    wire N__11271;
    wire N__11266;
    wire N__11265;
    wire N__11264;
    wire N__11263;
    wire N__11260;
    wire N__11253;
    wire N__11248;
    wire N__11247;
    wire N__11246;
    wire N__11245;
    wire N__11242;
    wire N__11239;
    wire N__11232;
    wire N__11227;
    wire N__11226;
    wire N__11225;
    wire N__11222;
    wire N__11217;
    wire N__11212;
    wire N__11211;
    wire N__11210;
    wire N__11207;
    wire N__11204;
    wire N__11201;
    wire N__11194;
    wire N__11191;
    wire N__11188;
    wire N__11185;
    wire N__11182;
    wire N__11179;
    wire N__11178;
    wire N__11177;
    wire N__11176;
    wire N__11173;
    wire N__11170;
    wire N__11165;
    wire N__11158;
    wire N__11155;
    wire N__11152;
    wire N__11149;
    wire N__11146;
    wire N__11143;
    wire N__11140;
    wire N__11137;
    wire N__11134;
    wire N__11131;
    wire N__11128;
    wire N__11127;
    wire N__11124;
    wire N__11123;
    wire N__11122;
    wire N__11119;
    wire N__11116;
    wire N__11113;
    wire N__11110;
    wire N__11107;
    wire N__11106;
    wire N__11103;
    wire N__11100;
    wire N__11097;
    wire N__11094;
    wire N__11091;
    wire N__11086;
    wire N__11079;
    wire N__11074;
    wire N__11073;
    wire N__11070;
    wire N__11069;
    wire N__11066;
    wire N__11065;
    wire N__11064;
    wire N__11061;
    wire N__11058;
    wire N__11055;
    wire N__11052;
    wire N__11049;
    wire N__11044;
    wire N__11041;
    wire N__11038;
    wire N__11035;
    wire N__11032;
    wire N__11027;
    wire N__11024;
    wire N__11017;
    wire N__11016;
    wire N__11013;
    wire N__11012;
    wire N__11011;
    wire N__11008;
    wire N__11005;
    wire N__11000;
    wire N__10993;
    wire N__10992;
    wire N__10989;
    wire N__10988;
    wire N__10985;
    wire N__10982;
    wire N__10981;
    wire N__10978;
    wire N__10973;
    wire N__10970;
    wire N__10963;
    wire N__10960;
    wire N__10957;
    wire N__10954;
    wire N__10951;
    wire N__10948;
    wire N__10945;
    wire N__10942;
    wire N__10939;
    wire N__10936;
    wire N__10933;
    wire N__10930;
    wire N__10927;
    wire N__10924;
    wire N__10921;
    wire N__10918;
    wire N__10915;
    wire N__10912;
    wire N__10909;
    wire N__10906;
    wire N__10903;
    wire N__10900;
    wire N__10897;
    wire N__10894;
    wire N__10891;
    wire N__10888;
    wire N__10885;
    wire N__10882;
    wire N__10879;
    wire N__10876;
    wire N__10873;
    wire N__10870;
    wire N__10867;
    wire N__10864;
    wire N__10861;
    wire N__10858;
    wire N__10855;
    wire N__10852;
    wire N__10849;
    wire N__10846;
    wire N__10843;
    wire N__10840;
    wire N__10837;
    wire N__10834;
    wire N__10831;
    wire N__10828;
    wire N__10827;
    wire N__10824;
    wire N__10821;
    wire N__10818;
    wire N__10815;
    wire N__10812;
    wire N__10809;
    wire N__10806;
    wire N__10803;
    wire N__10800;
    wire N__10797;
    wire N__10794;
    wire N__10791;
    wire N__10788;
    wire N__10785;
    wire N__10782;
    wire N__10779;
    wire N__10776;
    wire N__10773;
    wire N__10770;
    wire N__10767;
    wire N__10764;
    wire N__10761;
    wire N__10758;
    wire N__10755;
    wire N__10752;
    wire N__10749;
    wire N__10746;
    wire N__10743;
    wire N__10740;
    wire N__10737;
    wire N__10734;
    wire N__10731;
    wire N__10728;
    wire N__10725;
    wire N__10722;
    wire N__10719;
    wire N__10716;
    wire N__10713;
    wire N__10710;
    wire N__10707;
    wire N__10704;
    wire N__10701;
    wire N__10698;
    wire N__10695;
    wire N__10692;
    wire N__10689;
    wire N__10686;
    wire N__10683;
    wire N__10680;
    wire N__10677;
    wire N__10674;
    wire N__10671;
    wire N__10668;
    wire N__10665;
    wire N__10662;
    wire N__10659;
    wire N__10656;
    wire N__10653;
    wire N__10650;
    wire N__10647;
    wire N__10644;
    wire N__10641;
    wire N__10638;
    wire N__10635;
    wire N__10632;
    wire N__10629;
    wire N__10626;
    wire N__10623;
    wire N__10618;
    wire N__10615;
    wire N__10614;
    wire N__10613;
    wire N__10610;
    wire N__10609;
    wire N__10604;
    wire N__10599;
    wire N__10594;
    wire N__10591;
    wire N__10590;
    wire N__10585;
    wire N__10584;
    wire N__10583;
    wire N__10580;
    wire N__10575;
    wire N__10570;
    wire N__10567;
    wire N__10564;
    wire N__10561;
    wire N__10558;
    wire N__10557;
    wire N__10556;
    wire N__10553;
    wire N__10548;
    wire N__10547;
    wire N__10546;
    wire N__10545;
    wire N__10542;
    wire N__10539;
    wire N__10532;
    wire N__10525;
    wire N__10522;
    wire N__10521;
    wire N__10518;
    wire N__10515;
    wire N__10510;
    wire N__10507;
    wire N__10504;
    wire N__10501;
    wire N__10498;
    wire N__10495;
    wire N__10492;
    wire N__10491;
    wire N__10490;
    wire N__10489;
    wire N__10486;
    wire N__10485;
    wire N__10480;
    wire N__10477;
    wire N__10474;
    wire N__10471;
    wire N__10468;
    wire N__10459;
    wire N__10456;
    wire N__10455;
    wire N__10452;
    wire N__10449;
    wire N__10444;
    wire N__10441;
    wire N__10438;
    wire N__10435;
    wire N__10432;
    wire N__10431;
    wire N__10428;
    wire N__10425;
    wire N__10422;
    wire N__10419;
    wire N__10416;
    wire N__10413;
    wire N__10410;
    wire N__10407;
    wire N__10404;
    wire N__10401;
    wire N__10398;
    wire N__10395;
    wire N__10392;
    wire N__10389;
    wire N__10386;
    wire N__10383;
    wire N__10380;
    wire N__10377;
    wire N__10374;
    wire N__10371;
    wire N__10368;
    wire N__10365;
    wire N__10362;
    wire N__10359;
    wire N__10356;
    wire N__10353;
    wire N__10350;
    wire N__10347;
    wire N__10344;
    wire N__10341;
    wire N__10338;
    wire N__10335;
    wire N__10332;
    wire N__10329;
    wire N__10326;
    wire N__10323;
    wire N__10320;
    wire N__10317;
    wire N__10314;
    wire N__10311;
    wire N__10308;
    wire N__10305;
    wire N__10302;
    wire N__10299;
    wire N__10296;
    wire N__10293;
    wire N__10290;
    wire N__10287;
    wire N__10284;
    wire N__10281;
    wire N__10278;
    wire N__10275;
    wire N__10272;
    wire N__10269;
    wire N__10266;
    wire N__10263;
    wire N__10260;
    wire N__10257;
    wire N__10254;
    wire N__10251;
    wire N__10248;
    wire N__10245;
    wire N__10242;
    wire N__10239;
    wire N__10236;
    wire N__10233;
    wire N__10230;
    wire N__10227;
    wire N__10224;
    wire N__10221;
    wire N__10216;
    wire N__10213;
    wire N__10210;
    wire N__10207;
    wire N__10204;
    wire N__10201;
    wire N__10198;
    wire N__10195;
    wire N__10192;
    wire N__10189;
    wire N__10188;
    wire N__10183;
    wire N__10180;
    wire N__10179;
    wire N__10178;
    wire N__10177;
    wire N__10172;
    wire N__10169;
    wire N__10166;
    wire N__10163;
    wire N__10156;
    wire N__10155;
    wire N__10154;
    wire N__10153;
    wire N__10150;
    wire N__10147;
    wire N__10142;
    wire N__10135;
    wire N__10134;
    wire N__10133;
    wire N__10130;
    wire N__10125;
    wire N__10120;
    wire N__10119;
    wire N__10118;
    wire N__10117;
    wire N__10114;
    wire N__10111;
    wire N__10106;
    wire N__10099;
    wire N__10096;
    wire N__10095;
    wire N__10094;
    wire N__10093;
    wire N__10090;
    wire N__10087;
    wire N__10082;
    wire N__10075;
    wire N__10074;
    wire N__10073;
    wire N__10072;
    wire N__10069;
    wire N__10066;
    wire N__10061;
    wire N__10054;
    wire N__10053;
    wire N__10052;
    wire N__10051;
    wire N__10050;
    wire N__10049;
    wire N__10046;
    wire N__10043;
    wire N__10040;
    wire N__10039;
    wire N__10036;
    wire N__10035;
    wire N__10032;
    wire N__10029;
    wire N__10028;
    wire N__10025;
    wire N__10024;
    wire N__10021;
    wire N__10018;
    wire N__10015;
    wire N__10012;
    wire N__10009;
    wire N__10006;
    wire N__10003;
    wire N__10000;
    wire N__9997;
    wire N__9994;
    wire N__9989;
    wire N__9986;
    wire N__9981;
    wire N__9976;
    wire N__9973;
    wire N__9968;
    wire N__9965;
    wire N__9962;
    wire N__9959;
    wire N__9954;
    wire N__9951;
    wire N__9940;
    wire N__9937;
    wire N__9934;
    wire N__9931;
    wire N__9928;
    wire N__9925;
    wire N__9922;
    wire N__9919;
    wire N__9916;
    wire N__9913;
    wire N__9910;
    wire N__9907;
    wire N__9904;
    wire N__9901;
    wire N__9898;
    wire N__9895;
    wire N__9892;
    wire N__9889;
    wire N__9886;
    wire N__9883;
    wire N__9880;
    wire N__9877;
    wire N__9874;
    wire N__9871;
    wire N__9868;
    wire N__9865;
    wire N__9862;
    wire N__9859;
    wire N__9856;
    wire N__9853;
    wire N__9850;
    wire N__9849;
    wire N__9846;
    wire N__9843;
    wire N__9838;
    wire N__9835;
    wire N__9832;
    wire N__9829;
    wire N__9826;
    wire N__9823;
    wire N__9820;
    wire N__9817;
    wire N__9814;
    wire N__9811;
    wire N__9808;
    wire N__9805;
    wire N__9802;
    wire N__9799;
    wire N__9796;
    wire N__9793;
    wire N__9790;
    wire N__9787;
    wire N__9786;
    wire N__9783;
    wire N__9782;
    wire N__9779;
    wire N__9778;
    wire N__9775;
    wire N__9772;
    wire N__9769;
    wire N__9766;
    wire N__9759;
    wire N__9754;
    wire N__9751;
    wire N__9748;
    wire N__9745;
    wire N__9742;
    wire N__9739;
    wire N__9736;
    wire N__9733;
    wire N__9730;
    wire N__9727;
    wire N__9724;
    wire N__9721;
    wire N__9718;
    wire N__9715;
    wire N__9712;
    wire N__9709;
    wire N__9706;
    wire N__9703;
    wire N__9700;
    wire N__9697;
    wire N__9694;
    wire N__9691;
    wire N__9690;
    wire N__9689;
    wire N__9688;
    wire N__9683;
    wire N__9680;
    wire N__9677;
    wire N__9674;
    wire N__9667;
    wire N__9664;
    wire N__9663;
    wire N__9662;
    wire N__9661;
    wire N__9658;
    wire N__9655;
    wire N__9652;
    wire N__9649;
    wire N__9640;
    wire N__9639;
    wire N__9636;
    wire N__9635;
    wire N__9630;
    wire N__9629;
    wire N__9626;
    wire N__9623;
    wire N__9620;
    wire N__9613;
    wire N__9612;
    wire N__9607;
    wire N__9606;
    wire N__9603;
    wire N__9602;
    wire N__9599;
    wire N__9596;
    wire N__9593;
    wire N__9586;
    wire N__9583;
    wire N__9580;
    wire N__9577;
    wire N__9576;
    wire N__9575;
    wire N__9574;
    wire N__9569;
    wire N__9566;
    wire N__9563;
    wire N__9556;
    wire N__9553;
    wire N__9552;
    wire N__9551;
    wire N__9550;
    wire N__9545;
    wire N__9542;
    wire N__9539;
    wire N__9532;
    wire N__9529;
    wire N__9526;
    wire N__9523;
    wire N__9520;
    wire N__9517;
    wire N__9514;
    wire N__9511;
    wire N__9508;
    wire N__9505;
    wire N__9502;
    wire N__9499;
    wire N__9496;
    wire N__9493;
    wire N__9490;
    wire N__9487;
    wire N__9484;
    wire N__9481;
    wire N__9478;
    wire N__9475;
    wire N__9472;
    wire N__9469;
    wire N__9466;
    wire N__9463;
    wire N__9460;
    wire N__9457;
    wire N__9454;
    wire N__9451;
    wire N__9448;
    wire N__9445;
    wire N__9442;
    wire N__9439;
    wire N__9436;
    wire N__9433;
    wire N__9432;
    wire N__9427;
    wire N__9424;
    wire N__9421;
    wire N__9420;
    wire N__9419;
    wire N__9416;
    wire N__9415;
    wire N__9412;
    wire N__9409;
    wire N__9406;
    wire N__9403;
    wire N__9394;
    wire N__9393;
    wire N__9392;
    wire N__9391;
    wire N__9388;
    wire N__9385;
    wire N__9382;
    wire N__9379;
    wire N__9370;
    wire N__9367;
    wire N__9364;
    wire N__9361;
    wire N__9358;
    wire N__9355;
    wire N__9352;
    wire N__9349;
    wire N__9346;
    wire N__9343;
    wire N__9340;
    wire N__9337;
    wire N__9334;
    wire N__9331;
    wire N__9328;
    wire N__9325;
    wire N__9322;
    wire N__9319;
    wire N__9316;
    wire N__9313;
    wire N__9310;
    wire N__9307;
    wire N__9304;
    wire N__9301;
    wire N__9298;
    wire N__9295;
    wire N__9292;
    wire N__9289;
    wire N__9286;
    wire N__9283;
    wire N__9280;
    wire N__9277;
    wire N__9274;
    wire N__9271;
    wire N__9268;
    wire N__9265;
    wire N__9262;
    wire N__9259;
    wire N__9256;
    wire N__9253;
    wire N__9250;
    wire N__9247;
    wire N__9244;
    wire N__9241;
    wire N__9238;
    wire N__9235;
    wire N__9232;
    wire N__9229;
    wire N__9226;
    wire N__9223;
    wire N__9220;
    wire N__9217;
    wire N__9214;
    wire N__9211;
    wire N__9208;
    wire N__9207;
    wire N__9206;
    wire N__9203;
    wire N__9198;
    wire N__9193;
    wire N__9190;
    wire N__9189;
    wire N__9188;
    wire N__9187;
    wire N__9184;
    wire N__9181;
    wire N__9174;
    wire N__9169;
    wire N__9166;
    wire N__9165;
    wire N__9164;
    wire N__9163;
    wire N__9160;
    wire N__9153;
    wire N__9148;
    wire N__9145;
    wire N__9142;
    wire N__9139;
    wire N__9136;
    wire N__9133;
    wire N__9130;
    wire N__9127;
    wire N__9124;
    wire N__9121;
    wire N__9118;
    wire N__9115;
    wire N__9112;
    wire N__9109;
    wire N__9106;
    wire N__9103;
    wire N__9100;
    wire N__9097;
    wire N__9094;
    wire N__9091;
    wire N__9088;
    wire N__9085;
    wire N__9082;
    wire N__9079;
    wire N__9076;
    wire N__9073;
    wire N__9070;
    wire N__9067;
    wire N__9064;
    wire N__9061;
    wire N__9058;
    wire N__9055;
    wire N__9052;
    wire N__9049;
    wire N__9046;
    wire N__9043;
    wire N__9040;
    wire N__9037;
    wire N__9034;
    wire N__9031;
    wire N__9028;
    wire N__9025;
    wire N__9022;
    wire N__9019;
    wire N__9016;
    wire N__9013;
    wire N__9010;
    wire N__9007;
    wire N__9004;
    wire N__9001;
    wire N__8998;
    wire N__8995;
    wire N__8992;
    wire N__8989;
    wire N__8986;
    wire N__8983;
    wire N__8980;
    wire N__8977;
    wire N__8974;
    wire N__8971;
    wire N__8968;
    wire N__8965;
    wire N__8962;
    wire N__8959;
    wire N__8956;
    wire N__8953;
    wire N__8950;
    wire N__8947;
    wire N__8944;
    wire N__8941;
    wire N__8938;
    wire N__8935;
    wire N__8932;
    wire N__8929;
    wire N__8926;
    wire N__8923;
    wire N__8920;
    wire N__8917;
    wire N__8914;
    wire N__8911;
    wire N__8908;
    wire N__8905;
    wire N__8902;
    wire N__8899;
    wire N__8896;
    wire N__8893;
    wire N__8890;
    wire N__8887;
    wire N__8884;
    wire N__8881;
    wire N__8878;
    wire N__8875;
    wire N__8874;
    wire N__8871;
    wire N__8868;
    wire N__8863;
    wire N__8862;
    wire N__8859;
    wire N__8856;
    wire N__8855;
    wire N__8850;
    wire N__8847;
    wire N__8842;
    wire N__8841;
    wire N__8840;
    wire N__8837;
    wire N__8834;
    wire N__8831;
    wire N__8826;
    wire N__8823;
    wire N__8822;
    wire N__8819;
    wire N__8816;
    wire N__8813;
    wire N__8810;
    wire N__8809;
    wire N__8806;
    wire N__8803;
    wire N__8800;
    wire N__8797;
    wire N__8792;
    wire N__8787;
    wire N__8784;
    wire N__8781;
    wire N__8778;
    wire N__8775;
    wire N__8770;
    wire N__8767;
    wire N__8764;
    wire N__8761;
    wire N__8758;
    wire N__8755;
    wire N__8754;
    wire N__8753;
    wire N__8750;
    wire N__8747;
    wire N__8744;
    wire N__8741;
    wire N__8740;
    wire N__8739;
    wire N__8734;
    wire N__8731;
    wire N__8728;
    wire N__8727;
    wire N__8724;
    wire N__8721;
    wire N__8716;
    wire N__8713;
    wire N__8712;
    wire N__8711;
    wire N__8708;
    wire N__8701;
    wire N__8698;
    wire N__8695;
    wire N__8692;
    wire N__8689;
    wire N__8686;
    wire N__8683;
    wire N__8680;
    wire N__8677;
    wire N__8674;
    wire N__8671;
    wire N__8668;
    wire N__8665;
    wire N__8662;
    wire N__8659;
    wire N__8654;
    wire N__8649;
    wire N__8644;
    wire N__8641;
    wire N__8640;
    wire N__8639;
    wire N__8636;
    wire N__8633;
    wire N__8630;
    wire N__8629;
    wire N__8628;
    wire N__8621;
    wire N__8618;
    wire N__8615;
    wire N__8614;
    wire N__8609;
    wire N__8606;
    wire N__8603;
    wire N__8600;
    wire N__8597;
    wire N__8594;
    wire N__8593;
    wire N__8588;
    wire N__8585;
    wire N__8582;
    wire N__8579;
    wire N__8576;
    wire N__8573;
    wire N__8572;
    wire N__8569;
    wire N__8566;
    wire N__8563;
    wire N__8560;
    wire N__8551;
    wire N__8548;
    wire N__8545;
    wire N__8544;
    wire N__8541;
    wire N__8538;
    wire N__8537;
    wire N__8534;
    wire N__8533;
    wire N__8532;
    wire N__8529;
    wire N__8526;
    wire N__8523;
    wire N__8520;
    wire N__8517;
    wire N__8516;
    wire N__8513;
    wire N__8510;
    wire N__8505;
    wire N__8502;
    wire N__8501;
    wire N__8500;
    wire N__8497;
    wire N__8494;
    wire N__8491;
    wire N__8488;
    wire N__8485;
    wire N__8482;
    wire N__8479;
    wire N__8476;
    wire N__8473;
    wire N__8470;
    wire N__8467;
    wire N__8462;
    wire N__8459;
    wire N__8456;
    wire N__8453;
    wire N__8448;
    wire N__8443;
    wire N__8440;
    wire N__8431;
    wire N__8430;
    wire N__8427;
    wire N__8424;
    wire N__8421;
    wire N__8420;
    wire N__8417;
    wire N__8414;
    wire N__8411;
    wire N__8410;
    wire N__8407;
    wire N__8402;
    wire N__8399;
    wire N__8396;
    wire N__8395;
    wire N__8390;
    wire N__8389;
    wire N__8386;
    wire N__8383;
    wire N__8382;
    wire N__8379;
    wire N__8376;
    wire N__8371;
    wire N__8368;
    wire N__8363;
    wire N__8358;
    wire N__8357;
    wire N__8354;
    wire N__8351;
    wire N__8348;
    wire N__8345;
    wire N__8340;
    wire N__8337;
    wire N__8334;
    wire N__8329;
    wire N__8326;
    wire N__8325;
    wire N__8322;
    wire N__8321;
    wire N__8318;
    wire N__8315;
    wire N__8314;
    wire N__8311;
    wire N__8308;
    wire N__8307;
    wire N__8304;
    wire N__8301;
    wire N__8298;
    wire N__8295;
    wire N__8292;
    wire N__8291;
    wire N__8286;
    wire N__8285;
    wire N__8282;
    wire N__8277;
    wire N__8274;
    wire N__8271;
    wire N__8268;
    wire N__8265;
    wire N__8260;
    wire N__8255;
    wire N__8254;
    wire N__8251;
    wire N__8248;
    wire N__8245;
    wire N__8242;
    wire N__8237;
    wire N__8232;
    wire N__8229;
    wire N__8226;
    wire N__8221;
    wire N__8218;
    wire N__8215;
    wire N__8214;
    wire N__8213;
    wire N__8212;
    wire N__8209;
    wire N__8206;
    wire N__8205;
    wire N__8202;
    wire N__8201;
    wire N__8198;
    wire N__8193;
    wire N__8190;
    wire N__8187;
    wire N__8184;
    wire N__8181;
    wire N__8176;
    wire N__8173;
    wire N__8170;
    wire N__8169;
    wire N__8166;
    wire N__8163;
    wire N__8160;
    wire N__8157;
    wire N__8154;
    wire N__8151;
    wire N__8148;
    wire N__8145;
    wire N__8142;
    wire N__8139;
    wire N__8138;
    wire N__8135;
    wire N__8132;
    wire N__8125;
    wire N__8122;
    wire N__8119;
    wire N__8116;
    wire N__8113;
    wire N__8110;
    wire N__8107;
    wire N__8104;
    wire N__8101;
    wire N__8098;
    wire N__8089;
    wire N__8088;
    wire N__8085;
    wire N__8082;
    wire N__8081;
    wire N__8078;
    wire N__8075;
    wire N__8072;
    wire N__8071;
    wire N__8068;
    wire N__8065;
    wire N__8062;
    wire N__8061;
    wire N__8058;
    wire N__8057;
    wire N__8056;
    wire N__8053;
    wire N__8050;
    wire N__8047;
    wire N__8044;
    wire N__8041;
    wire N__8038;
    wire N__8037;
    wire N__8034;
    wire N__8029;
    wire N__8026;
    wire N__8023;
    wire N__8020;
    wire N__8017;
    wire N__8014;
    wire N__8011;
    wire N__8006;
    wire N__8003;
    wire N__7996;
    wire N__7993;
    wire N__7988;
    wire N__7985;
    wire N__7982;
    wire TVP_VIDEO_c_3;
    wire VCCG0;
    wire TVP_VIDEO_c_5;
    wire TVP_VIDEO_c_4;
    wire TVP_VIDEO_c_7;
    wire TVP_VIDEO_c_6;
    wire TVP_VIDEO_c_8;
    wire TVP_VIDEO_c_9;
    wire TVP_VIDEO_c_2;
    wire GNDG0;
    wire \transmit_module.X_DELTA_PATTERN_3 ;
    wire \transmit_module.X_DELTA_PATTERN_2 ;
    wire \transmit_module.X_DELTA_PATTERN_4 ;
    wire \transmit_module.X_DELTA_PATTERN_9 ;
    wire \transmit_module.Y_DELTA_PATTERN_87 ;
    wire \transmit_module.Y_DELTA_PATTERN_89 ;
    wire \transmit_module.Y_DELTA_PATTERN_88 ;
    wire \transmit_module.Y_DELTA_PATTERN_90 ;
    wire \transmit_module.Y_DELTA_PATTERN_91 ;
    wire \transmit_module.Y_DELTA_PATTERN_77 ;
    wire \transmit_module.Y_DELTA_PATTERN_92 ;
    wire \transmit_module.Y_DELTA_PATTERN_93 ;
    wire \transmit_module.Y_DELTA_PATTERN_95 ;
    wire \transmit_module.Y_DELTA_PATTERN_94 ;
    wire \transmit_module.X_DELTA_PATTERN_8 ;
    wire \transmit_module.X_DELTA_PATTERN_7 ;
    wire \transmit_module.X_DELTA_PATTERN_10 ;
    wire \transmit_module.X_DELTA_PATTERN_6 ;
    wire \transmit_module.X_DELTA_PATTERN_5 ;
    wire \transmit_module.X_DELTA_PATTERN_15 ;
    wire \transmit_module.X_DELTA_PATTERN_12 ;
    wire \transmit_module.X_DELTA_PATTERN_11 ;
    wire \transmit_module.X_DELTA_PATTERN_14 ;
    wire \transmit_module.X_DELTA_PATTERN_13 ;
    wire \transmit_module.Y_DELTA_PATTERN_64 ;
    wire \transmit_module.Y_DELTA_PATTERN_65 ;
    wire \transmit_module.Y_DELTA_PATTERN_41 ;
    wire \transmit_module.Y_DELTA_PATTERN_63 ;
    wire \transmit_module.Y_DELTA_PATTERN_74 ;
    wire \transmit_module.Y_DELTA_PATTERN_76 ;
    wire \transmit_module.Y_DELTA_PATTERN_75 ;
    wire \transmit_module.Y_DELTA_PATTERN_73 ;
    wire \transmit_module.Y_DELTA_PATTERN_48 ;
    wire \transmit_module.Y_DELTA_PATTERN_47 ;
    wire \transmit_module.Y_DELTA_PATTERN_46 ;
    wire \transmit_module.Y_DELTA_PATTERN_42 ;
    wire \transmit_module.Y_DELTA_PATTERN_96 ;
    wire \transmit_module.Y_DELTA_PATTERN_45 ;
    wire \transmit_module.Y_DELTA_PATTERN_44 ;
    wire \transmit_module.Y_DELTA_PATTERN_43 ;
    wire \transmit_module.video_signal_controller.n3788_cascade_ ;
    wire \transmit_module.video_signal_controller.n2876 ;
    wire \transmit_module.video_signal_controller.VGA_X_0 ;
    wire bfn_10_15_0_;
    wire \transmit_module.video_signal_controller.VGA_X_1 ;
    wire \transmit_module.video_signal_controller.n3279 ;
    wire \transmit_module.video_signal_controller.VGA_X_2 ;
    wire \transmit_module.video_signal_controller.n3280 ;
    wire \transmit_module.video_signal_controller.n3281 ;
    wire \transmit_module.video_signal_controller.n3282 ;
    wire \transmit_module.video_signal_controller.n3283 ;
    wire \transmit_module.video_signal_controller.n3284 ;
    wire \transmit_module.video_signal_controller.n3285 ;
    wire \transmit_module.video_signal_controller.n3286 ;
    wire bfn_10_16_0_;
    wire \transmit_module.video_signal_controller.n3287 ;
    wire \transmit_module.video_signal_controller.n3288 ;
    wire \transmit_module.video_signal_controller.n3289 ;
    wire \transmit_module.Y_DELTA_PATTERN_55 ;
    wire \transmit_module.Y_DELTA_PATTERN_54 ;
    wire \transmit_module.Y_DELTA_PATTERN_40 ;
    wire \transmit_module.Y_DELTA_PATTERN_56 ;
    wire \transmit_module.Y_DELTA_PATTERN_97 ;
    wire \transmit_module.Y_DELTA_PATTERN_36 ;
    wire \transmit_module.Y_DELTA_PATTERN_62 ;
    wire \transmit_module.Y_DELTA_PATTERN_66 ;
    wire \transmit_module.Y_DELTA_PATTERN_53 ;
    wire \transmit_module.Y_DELTA_PATTERN_52 ;
    wire \transmit_module.Y_DELTA_PATTERN_51 ;
    wire \transmit_module.Y_DELTA_PATTERN_81 ;
    wire \transmit_module.Y_DELTA_PATTERN_50 ;
    wire \transmit_module.Y_DELTA_PATTERN_49 ;
    wire \transmit_module.Y_DELTA_PATTERN_35 ;
    wire \transmit_module.Y_DELTA_PATTERN_34 ;
    wire \transmit_module.Y_DELTA_PATTERN_72 ;
    wire \transmit_module.Y_DELTA_PATTERN_82 ;
    wire \transmit_module.Y_DELTA_PATTERN_69 ;
    wire \transmit_module.Y_DELTA_PATTERN_78 ;
    wire \transmit_module.Y_DELTA_PATTERN_80 ;
    wire \transmit_module.Y_DELTA_PATTERN_79 ;
    wire \transmit_module.Y_DELTA_PATTERN_71 ;
    wire \transmit_module.Y_DELTA_PATTERN_70 ;
    wire \transmit_module.Y_DELTA_PATTERN_68 ;
    wire \transmit_module.Y_DELTA_PATTERN_67 ;
    wire \transmit_module.video_signal_controller.n2886 ;
    wire \transmit_module.video_signal_controller.n1983_cascade_ ;
    wire \transmit_module.video_signal_controller.n2926 ;
    wire \transmit_module.video_signal_controller.n2010_cascade_ ;
    wire \transmit_module.video_signal_controller.n1983 ;
    wire \transmit_module.video_signal_controller.n3789 ;
    wire \transmit_module.video_signal_controller.n3467 ;
    wire \transmit_module.video_signal_controller.n18_cascade_ ;
    wire \transmit_module.video_signal_controller.VGA_X_3 ;
    wire \transmit_module.video_signal_controller.VGA_X_5 ;
    wire \transmit_module.video_signal_controller.VGA_X_8 ;
    wire \transmit_module.video_signal_controller.n4_adj_617_cascade_ ;
    wire \transmit_module.video_signal_controller.VGA_X_6 ;
    wire \transmit_module.video_signal_controller.VGA_X_9 ;
    wire \transmit_module.video_signal_controller.VGA_X_10 ;
    wire \transmit_module.video_signal_controller.n4 ;
    wire \transmit_module.video_signal_controller.VGA_X_7 ;
    wire \transmit_module.video_signal_controller.n3794_cascade_ ;
    wire \transmit_module.video_signal_controller.VGA_X_4 ;
    wire \transmit_module.video_signal_controller.n3618 ;
    wire \transmit_module.Y_DELTA_PATTERN_61 ;
    wire \transmit_module.Y_DELTA_PATTERN_37 ;
    wire \transmit_module.Y_DELTA_PATTERN_39 ;
    wire \transmit_module.Y_DELTA_PATTERN_38 ;
    wire \transmit_module.Y_DELTA_PATTERN_58 ;
    wire \transmit_module.Y_DELTA_PATTERN_57 ;
    wire \transmit_module.Y_DELTA_PATTERN_60 ;
    wire \transmit_module.Y_DELTA_PATTERN_59 ;
    wire \transmit_module.Y_DELTA_PATTERN_98 ;
    wire \transmit_module.Y_DELTA_PATTERN_86 ;
    wire \transmit_module.Y_DELTA_PATTERN_85 ;
    wire \transmit_module.Y_DELTA_PATTERN_84 ;
    wire \transmit_module.Y_DELTA_PATTERN_83 ;
    wire \transmit_module.Y_DELTA_PATTERN_99 ;
    wire bfn_12_13_0_;
    wire \transmit_module.video_signal_controller.n3290 ;
    wire \transmit_module.video_signal_controller.n3291 ;
    wire \transmit_module.video_signal_controller.n3292 ;
    wire \transmit_module.video_signal_controller.n3293 ;
    wire \transmit_module.video_signal_controller.n3294 ;
    wire \transmit_module.video_signal_controller.n3295 ;
    wire \transmit_module.video_signal_controller.n3296 ;
    wire \transmit_module.video_signal_controller.n3297 ;
    wire bfn_12_14_0_;
    wire \transmit_module.video_signal_controller.n3298 ;
    wire \transmit_module.video_signal_controller.n3299 ;
    wire \transmit_module.video_signal_controller.n3300 ;
    wire \transmit_module.video_signal_controller.n2010 ;
    wire \transmit_module.video_signal_controller.n2361 ;
    wire \transmit_module.n3787_cascade_ ;
    wire \transmit_module.Y_DELTA_PATTERN_7 ;
    wire \transmit_module.Y_DELTA_PATTERN_6 ;
    wire \transmit_module.Y_DELTA_PATTERN_5 ;
    wire \transmit_module.Y_DELTA_PATTERN_4 ;
    wire \transmit_module.Y_DELTA_PATTERN_3 ;
    wire \line_buffer.n578 ;
    wire \line_buffer.n570 ;
    wire \line_buffer.n577 ;
    wire \line_buffer.n569 ;
    wire bfn_13_10_0_;
    wire \receive_module.rx_counter.n3271 ;
    wire \receive_module.rx_counter.n3272 ;
    wire \receive_module.rx_counter.n3273 ;
    wire \receive_module.rx_counter.n3274 ;
    wire \receive_module.rx_counter.n3275 ;
    wire \receive_module.rx_counter.n3276 ;
    wire \receive_module.rx_counter.n3277 ;
    wire \receive_module.rx_counter.n3278 ;
    wire bfn_13_11_0_;
    wire \transmit_module.video_signal_controller.n3786_cascade_ ;
    wire \transmit_module.video_signal_controller.n8 ;
    wire \transmit_module.video_signal_controller.n7_adj_615_cascade_ ;
    wire \transmit_module.video_signal_controller.n2_cascade_ ;
    wire \transmit_module.video_signal_controller.n3785 ;
    wire \transmit_module.video_signal_controller.n3577_cascade_ ;
    wire \transmit_module.video_signal_controller.n3485 ;
    wire \transmit_module.video_signal_controller.VGA_Y_9 ;
    wire \transmit_module.video_signal_controller.VGA_Y_6 ;
    wire \transmit_module.video_signal_controller.VGA_Y_11 ;
    wire \transmit_module.video_signal_controller.VGA_Y_7 ;
    wire \transmit_module.video_signal_controller.VGA_Y_5 ;
    wire \transmit_module.video_signal_controller.VGA_Y_2 ;
    wire \transmit_module.n3798 ;
    wire \transmit_module.n112_cascade_ ;
    wire n24;
    wire \transmit_module.old_VGA_HS ;
    wire \transmit_module.VGA_VISIBLE_Y ;
    wire ADV_HSYNC_c;
    wire \transmit_module.video_signal_controller.n3486 ;
    wire \transmit_module.video_signal_controller.n7 ;
    wire \transmit_module.video_signal_controller.VGA_X_11 ;
    wire \transmit_module.video_signal_controller.VGA_VISIBLE_N_578 ;
    wire \transmit_module.n111_cascade_ ;
    wire n23;
    wire \transmit_module.ADDR_Y_COMPONENT_4 ;
    wire \transmit_module.ADDR_Y_COMPONENT_5 ;
    wire \line_buffer.n571 ;
    wire \line_buffer.n563 ;
    wire \line_buffer.n514 ;
    wire \line_buffer.n506 ;
    wire \line_buffer.n3764 ;
    wire \line_buffer.n513 ;
    wire \line_buffer.n505 ;
    wire \line_buffer.n3646_cascade_ ;
    wire \line_buffer.n3647 ;
    wire \receive_module.rx_counter.Y_3 ;
    wire \receive_module.rx_counter.Y_2 ;
    wire \receive_module.rx_counter.Y_1 ;
    wire \receive_module.rx_counter.Y_5 ;
    wire \receive_module.rx_counter.Y_6 ;
    wire \receive_module.rx_counter.n4_adj_604 ;
    wire \receive_module.rx_counter.n5_cascade_ ;
    wire \receive_module.rx_counter.n3548 ;
    wire \receive_module.rx_counter.Y_0 ;
    wire \receive_module.rx_counter.n14_adj_611 ;
    wire \receive_module.rx_counter.n10_adj_610 ;
    wire \transmit_module.ADDR_Y_COMPONENT_7 ;
    wire \transmit_module.X_DELTA_PATTERN_1 ;
    wire \transmit_module.n2093 ;
    wire \transmit_module.n2147 ;
    wire \transmit_module.video_signal_controller.VGA_Y_4 ;
    wire \transmit_module.video_signal_controller.VGA_Y_8 ;
    wire \transmit_module.video_signal_controller.VGA_Y_0 ;
    wire \transmit_module.video_signal_controller.VGA_Y_3 ;
    wire \transmit_module.video_signal_controller.n3626_cascade_ ;
    wire \transmit_module.video_signal_controller.VGA_Y_1 ;
    wire \transmit_module.n111 ;
    wire \transmit_module.n143 ;
    wire \transmit_module.n143_cascade_ ;
    wire \transmit_module.n112 ;
    wire \transmit_module.n142 ;
    wire \transmit_module.n141_cascade_ ;
    wire \transmit_module.n137_cascade_ ;
    wire \transmit_module.ADDR_Y_COMPONENT_1 ;
    wire \transmit_module.ADDR_Y_COMPONENT_10 ;
    wire \transmit_module.video_signal_controller.n3632 ;
    wire \transmit_module.video_signal_controller.n18_adj_616 ;
    wire \transmit_module.video_signal_controller.n3614 ;
    wire \transmit_module.video_signal_controller.VGA_Y_10 ;
    wire \transmit_module.n146 ;
    wire \transmit_module.n146_cascade_ ;
    wire \transmit_module.n115 ;
    wire n27;
    wire \transmit_module.Y_DELTA_PATTERN_2 ;
    wire \transmit_module.Y_DELTA_PATTERN_1 ;
    wire \transmit_module.Y_DELTA_PATTERN_9 ;
    wire \transmit_module.Y_DELTA_PATTERN_8 ;
    wire \transmit_module.Y_DELTA_PATTERN_10 ;
    wire \line_buffer.n507 ;
    wire \line_buffer.n499 ;
    wire \line_buffer.n3752 ;
    wire \transmit_module.ADDR_Y_COMPONENT_6 ;
    wire \transmit_module.n106 ;
    wire \transmit_module.n137 ;
    wire n18;
    wire \transmit_module.ADDR_Y_COMPONENT_0 ;
    wire \line_buffer.n3722 ;
    wire TX_DATA_6;
    wire n1792;
    wire n1798;
    wire \line_buffer.n448 ;
    wire \line_buffer.n440 ;
    wire \line_buffer.n3679 ;
    wire \transmit_module.n116 ;
    wire \transmit_module.n147 ;
    wire n28;
    wire \transmit_module.n110 ;
    wire \transmit_module.n141 ;
    wire n22;
    wire \transmit_module.n109 ;
    wire \transmit_module.n140 ;
    wire n21;
    wire LED_c;
    wire \receive_module.rx_counter.n3628_cascade_ ;
    wire \receive_module.rx_counter.n7_adj_609 ;
    wire \receive_module.rx_counter.n11 ;
    wire \receive_module.rx_counter.n11_cascade_ ;
    wire \receive_module.rx_counter.old_VS ;
    wire \line_buffer.n543 ;
    wire \line_buffer.n535 ;
    wire \receive_module.rx_counter.Y_7 ;
    wire \receive_module.rx_counter.n3791 ;
    wire \receive_module.rx_counter.Y_4 ;
    wire \receive_module.rx_counter.n3551 ;
    wire \receive_module.rx_counter.n2045 ;
    wire \receive_module.rx_counter.old_HS ;
    wire bfn_15_11_0_;
    wire \receive_module.n3245 ;
    wire \receive_module.n3246 ;
    wire \receive_module.n3247 ;
    wire \receive_module.n3248 ;
    wire \receive_module.n3249 ;
    wire \receive_module.n3250 ;
    wire \receive_module.n3251 ;
    wire \receive_module.n3252 ;
    wire bfn_15_12_0_;
    wire \receive_module.n3253 ;
    wire \receive_module.n3254 ;
    wire \receive_module.n3255 ;
    wire \receive_module.n3256 ;
    wire \receive_module.n3257 ;
    wire \transmit_module.TX_ADDR_0 ;
    wire \transmit_module.X_DELTA_PATTERN_0 ;
    wire \transmit_module.n132 ;
    wire bfn_15_13_0_;
    wire \transmit_module.TX_ADDR_1 ;
    wire \transmit_module.n131 ;
    wire \transmit_module.n3258 ;
    wire \transmit_module.n3259 ;
    wire \transmit_module.n3260 ;
    wire \transmit_module.TX_ADDR_4 ;
    wire \transmit_module.n128 ;
    wire \transmit_module.n3261 ;
    wire \transmit_module.TX_ADDR_5 ;
    wire \transmit_module.n127 ;
    wire \transmit_module.n3262 ;
    wire \transmit_module.TX_ADDR_6 ;
    wire \transmit_module.n126 ;
    wire \transmit_module.n3263 ;
    wire \transmit_module.TX_ADDR_7 ;
    wire \transmit_module.n125 ;
    wire \transmit_module.n3264 ;
    wire \transmit_module.n3265 ;
    wire bfn_15_14_0_;
    wire \transmit_module.n3266 ;
    wire \transmit_module.TX_ADDR_10 ;
    wire \transmit_module.n122 ;
    wire \transmit_module.n3267 ;
    wire \transmit_module.n3268 ;
    wire \transmit_module.n3269 ;
    wire \transmit_module.n3270 ;
    wire \transmit_module.ADDR_Y_COMPONENT_9 ;
    wire \transmit_module.ADDR_Y_COMPONENT_12 ;
    wire \transmit_module.n120 ;
    wire \transmit_module.n119 ;
    wire \transmit_module.ADDR_Y_COMPONENT_11 ;
    wire \transmit_module.n121 ;
    wire \transmit_module.n2039 ;
    wire \transmit_module.n130 ;
    wire \line_buffer.n3755 ;
    wire TX_DATA_0;
    wire \receive_module.n134 ;
    wire RX_ADDR_2;
    wire \line_buffer.n545 ;
    wire \line_buffer.n537 ;
    wire \line_buffer.n3680 ;
    wire \receive_module.n126 ;
    wire RX_ADDR_10;
    wire \receive_module.n132 ;
    wire RX_ADDR_4;
    wire \receive_module.n131 ;
    wire RX_ADDR_5;
    wire \receive_module.n130 ;
    wire RX_ADDR_6;
    wire \receive_module.n129 ;
    wire RX_ADDR_7;
    wire \receive_module.n128 ;
    wire RX_ADDR_8;
    wire \receive_module.n127 ;
    wire RX_ADDR_9;
    wire \receive_module.rx_counter.FRAME_COUNTER_0 ;
    wire bfn_16_5_0_;
    wire \receive_module.rx_counter.FRAME_COUNTER_1 ;
    wire \receive_module.rx_counter.n3310 ;
    wire \receive_module.rx_counter.FRAME_COUNTER_2 ;
    wire \receive_module.rx_counter.n3311 ;
    wire \receive_module.rx_counter.FRAME_COUNTER_3 ;
    wire \receive_module.rx_counter.n3312 ;
    wire \receive_module.rx_counter.FRAME_COUNTER_4 ;
    wire \receive_module.rx_counter.n3313 ;
    wire \receive_module.rx_counter.n3314 ;
    wire \receive_module.rx_counter.FRAME_COUNTER_5 ;
    wire \receive_module.rx_counter.n3792 ;
    wire \receive_module.rx_counter.n2517 ;
    wire \receive_module.n136 ;
    wire RX_ADDR_0;
    wire \receive_module.n135 ;
    wire RX_ADDR_1;
    wire \line_buffer.n511 ;
    wire \line_buffer.n503 ;
    wire \line_buffer.n509 ;
    wire \line_buffer.n501 ;
    wire \receive_module.rx_counter.n4_cascade_ ;
    wire \receive_module.rx_counter.n6_cascade_ ;
    wire \receive_module.rx_counter.n3534 ;
    wire \receive_module.rx_counter.n3581 ;
    wire \line_buffer.n517 ;
    wire \line_buffer.n452 ;
    wire \line_buffer.n548 ;
    wire \receive_module.n3795 ;
    wire \line_buffer.n451 ;
    wire \line_buffer.n549 ;
    wire \line_buffer.n516 ;
    wire \receive_module.rx_counter.n3575 ;
    wire \receive_module.rx_counter.n4_adj_606 ;
    wire \receive_module.rx_counter.Y_8 ;
    wire \receive_module.rx_counter.n55_adj_607 ;
    wire \line_buffer.n581 ;
    wire RX_ADDR_12;
    wire RX_ADDR_13;
    wire RX_ADDR_11;
    wire \line_buffer.n580 ;
    wire RX_TX_SYNC_BUFF;
    wire RX_TX_SYNC;
    wire \sync_buffer.BUFFER_0 ;
    wire \sync_buffer.BUFFER_1 ;
    wire \INVsync_buffer.WIRE_OUT_8C_net ;
    wire \transmit_module.n124 ;
    wire \transmit_module.n139_cascade_ ;
    wire \transmit_module.ADDR_Y_COMPONENT_8 ;
    wire \transmit_module.TX_ADDR_8 ;
    wire \transmit_module.TX_ADDR_9 ;
    wire \transmit_module.n123 ;
    wire \transmit_module.n138 ;
    wire \transmit_module.n138_cascade_ ;
    wire \transmit_module.n107 ;
    wire n19;
    wire \transmit_module.ADDR_Y_COMPONENT_13 ;
    wire \line_buffer.n3634 ;
    wire \line_buffer.n442 ;
    wire \line_buffer.n434 ;
    wire \line_buffer.n3749 ;
    wire \line_buffer.n541 ;
    wire \line_buffer.n533 ;
    wire \line_buffer.n3676 ;
    wire \line_buffer.n3674 ;
    wire \line_buffer.n3716 ;
    wire \line_buffer.n446 ;
    wire \line_buffer.n438 ;
    wire \line_buffer.n3728 ;
    wire \line_buffer.n3640_cascade_ ;
    wire \line_buffer.n3641 ;
    wire \transmit_module.n114 ;
    wire \transmit_module.n145 ;
    wire n26;
    wire \transmit_module.VGA_VISIBLE ;
    wire \transmit_module.n129 ;
    wire \transmit_module.n144 ;
    wire \transmit_module.n144_cascade_ ;
    wire n25;
    wire \transmit_module.TX_ADDR_2 ;
    wire \transmit_module.ADDR_Y_COMPONENT_2 ;
    wire \transmit_module.Y_DELTA_PATTERN_0 ;
    wire \transmit_module.n113 ;
    wire \transmit_module.TX_ADDR_3 ;
    wire \transmit_module.ADDR_Y_COMPONENT_3 ;
    wire \transmit_module.n2061 ;
    wire TX_DATA_4;
    wire n1794;
    wire TX_DATA_2;
    wire n1796;
    wire \line_buffer.n444 ;
    wire \line_buffer.n436 ;
    wire \line_buffer.n3673 ;
    wire \transmit_module.n3787 ;
    wire \transmit_module.n108 ;
    wire \transmit_module.n139 ;
    wire n20;
    wire GB_BUFFER_TVP_CLK_c_THRU_CO;
    wire TVP_HSYNC_c;
    wire \receive_module.rx_counter.n10 ;
    wire bfn_17_10_0_;
    wire \receive_module.rx_counter.n9 ;
    wire \receive_module.rx_counter.n3301 ;
    wire \receive_module.rx_counter.n8 ;
    wire \receive_module.rx_counter.n3302 ;
    wire \receive_module.rx_counter.X_3 ;
    wire \receive_module.rx_counter.n3303 ;
    wire \receive_module.rx_counter.X_4 ;
    wire \receive_module.rx_counter.n3304 ;
    wire \receive_module.rx_counter.X_5 ;
    wire \receive_module.rx_counter.n3305 ;
    wire \receive_module.rx_counter.X_6 ;
    wire \receive_module.rx_counter.n3306 ;
    wire \receive_module.rx_counter.X_7 ;
    wire \receive_module.rx_counter.n3307 ;
    wire \receive_module.rx_counter.n3308 ;
    wire \receive_module.rx_counter.X_8 ;
    wire bfn_17_11_0_;
    wire \receive_module.rx_counter.n3309 ;
    wire \receive_module.rx_counter.X_9 ;
    wire \receive_module.rx_counter.n3790 ;
    wire \line_buffer.n576 ;
    wire \line_buffer.n568 ;
    wire \line_buffer.n504 ;
    wire \line_buffer.n512 ;
    wire \line_buffer.n3734_cascade_ ;
    wire \transmit_module.Y_DELTA_PATTERN_12 ;
    wire \transmit_module.Y_DELTA_PATTERN_11 ;
    wire \transmit_module.Y_DELTA_PATTERN_25 ;
    wire \transmit_module.Y_DELTA_PATTERN_26 ;
    wire \transmit_module.Y_DELTA_PATTERN_13 ;
    wire \line_buffer.n539 ;
    wire \line_buffer.n531 ;
    wire \line_buffer.n3746 ;
    wire \line_buffer.n573 ;
    wire \line_buffer.n565 ;
    wire \line_buffer.n3677 ;
    wire \line_buffer.n567 ;
    wire \line_buffer.n575 ;
    wire \line_buffer.n3635 ;
    wire \line_buffer.n3737 ;
    wire \line_buffer.n447 ;
    wire \line_buffer.n439 ;
    wire \line_buffer.n3701 ;
    wire TX_DATA_5;
    wire n1793;
    wire CONSTANT_ONE_NET;
    wire \transmit_module.Y_DELTA_PATTERN_33 ;
    wire \transmit_module.Y_DELTA_PATTERN_27 ;
    wire \transmit_module.Y_DELTA_PATTERN_28 ;
    wire \transmit_module.Y_DELTA_PATTERN_29 ;
    wire \transmit_module.Y_DELTA_PATTERN_30 ;
    wire \transmit_module.Y_DELTA_PATTERN_32 ;
    wire \transmit_module.Y_DELTA_PATTERN_31 ;
    wire \transmit_module.Y_DELTA_PATTERN_22 ;
    wire \transmit_module.Y_DELTA_PATTERN_24 ;
    wire \transmit_module.Y_DELTA_PATTERN_23 ;
    wire \transmit_module.Y_DELTA_PATTERN_16 ;
    wire \transmit_module.Y_DELTA_PATTERN_17 ;
    wire \transmit_module.Y_DELTA_PATTERN_19 ;
    wire \transmit_module.Y_DELTA_PATTERN_18 ;
    wire \transmit_module.Y_DELTA_PATTERN_15 ;
    wire \transmit_module.Y_DELTA_PATTERN_14 ;
    wire n1797;
    wire \transmit_module.Y_DELTA_PATTERN_21 ;
    wire \transmit_module.Y_DELTA_PATTERN_20 ;
    wire \transmit_module.n3797 ;
    wire ADV_VSYNC_c;
    wire \line_buffer.n544 ;
    wire \line_buffer.n536 ;
    wire \line_buffer.n3698 ;
    wire \line_buffer.n508 ;
    wire \line_buffer.n500 ;
    wire \line_buffer.n3695_cascade_ ;
    wire TX_DATA_1;
    wire \line_buffer.n572 ;
    wire \line_buffer.n564 ;
    wire \line_buffer.n3692 ;
    wire RX_WE;
    wire \receive_module.n133 ;
    wire TVP_VSYNC_c;
    wire RX_ADDR_3;
    wire TVP_CLK_c;
    wire \receive_module.n3793 ;
    wire \line_buffer.n542 ;
    wire \line_buffer.n534 ;
    wire \line_buffer.n445 ;
    wire \line_buffer.n437 ;
    wire \line_buffer.n3710 ;
    wire \line_buffer.n566 ;
    wire \line_buffer.n574 ;
    wire \line_buffer.n502 ;
    wire \line_buffer.n510 ;
    wire \line_buffer.n3758_cascade_ ;
    wire \line_buffer.n540 ;
    wire \line_buffer.n532 ;
    wire \line_buffer.n435 ;
    wire \line_buffer.n443 ;
    wire \line_buffer.n3740_cascade_ ;
    wire \line_buffer.n3743 ;
    wire \line_buffer.n3761 ;
    wire \line_buffer.n3713 ;
    wire TX_ADDR_13;
    wire \line_buffer.n3767 ;
    wire TX_ADDR_11;
    wire \line_buffer.n546 ;
    wire \line_buffer.n538 ;
    wire TX_DATA_3;
    wire n1795;
    wire TX_DATA_7;
    wire ADV_B_c;
    wire ADV_CLK_c;
    wire \transmit_module.n2354 ;
    wire \line_buffer.n449 ;
    wire TX_ADDR_12;
    wire \line_buffer.n441 ;
    wire \line_buffer.n3704 ;
    wire \line_buffer.n3707 ;
    wire _gnd_net_;

    defparam \tx_pll.TX_PLL_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \tx_pll.TX_PLL_inst .TEST_MODE=1'b0;
    defparam \tx_pll.TX_PLL_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \tx_pll.TX_PLL_inst .PLLOUT_SELECT="GENCLK";
    defparam \tx_pll.TX_PLL_inst .FILTER_RANGE=3'b010;
    defparam \tx_pll.TX_PLL_inst .FEEDBACK_PATH="SIMPLE";
    defparam \tx_pll.TX_PLL_inst .FDA_RELATIVE=4'b0000;
    defparam \tx_pll.TX_PLL_inst .FDA_FEEDBACK=4'b0000;
    defparam \tx_pll.TX_PLL_inst .ENABLE_ICEGATE=1'b0;
    defparam \tx_pll.TX_PLL_inst .DIVR=4'b0000;
    defparam \tx_pll.TX_PLL_inst .DIVQ=3'b100;
    defparam \tx_pll.TX_PLL_inst .DIVF=7'b0100110;
    defparam \tx_pll.TX_PLL_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \tx_pll.TX_PLL_inst  (
            .EXTFEEDBACK(),
            .LATCHINPUTVALUE(),
            .SCLK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(ADV_CLK_c),
            .REFERENCECLK(N__18664),
            .RESETB(N__19656),
            .BYPASS(GNDG0),
            .SDI(),
            .DYNAMICDELAY({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7}),
            .PLLOUTGLOBAL());
    defparam \line_buffer.mem2_physical .WRITE_MODE=3;
    defparam \line_buffer.mem2_physical .READ_MODE=3;
    defparam \line_buffer.mem2_physical .INIT_F=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem2_physical .INIT_E=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem2_physical .INIT_D=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem2_physical .INIT_C=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem2_physical .INIT_B=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem2_physical .INIT_A=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem2_physical .INIT_9=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem2_physical .INIT_8=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem2_physical .INIT_7=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem2_physical .INIT_6=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem2_physical .INIT_5=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem2_physical .INIT_4=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem2_physical .INIT_3=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem2_physical .INIT_2=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem2_physical .INIT_1=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem2_physical .INIT_0=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    SB_RAM40_4K \line_buffer.mem2_physical  (
            .RDATA({dangling_wire_8,dangling_wire_9,dangling_wire_10,dangling_wire_11,\line_buffer.n449 ,dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,\line_buffer.n448 ,dangling_wire_19,dangling_wire_20,dangling_wire_21}),
            .RADDR({N__12333,N__17139,N__18750,N__12621,N__12885,N__10308,N__10683,N__18051,N__18399,N__11649,N__11892}),
            .WADDR({N__15513,N__13995,N__14256,N__14505,N__14760,N__15021,N__15258,N__20280,N__13641,N__15816,N__16071}),
            .MASK({dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29,dangling_wire_30,dangling_wire_31,dangling_wire_32,dangling_wire_33,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37}),
            .WDATA({dangling_wire_38,dangling_wire_39,dangling_wire_40,dangling_wire_41,N__8614,dangling_wire_42,dangling_wire_43,dangling_wire_44,dangling_wire_45,dangling_wire_46,dangling_wire_47,dangling_wire_48,N__8739,dangling_wire_49,dangling_wire_50,dangling_wire_51}),
            .RCLKE(),
            .RCLK(N__22913),
            .RE(N__19629),
            .WCLKE(),
            .WCLK(N__20171),
            .WE(N__16447));
    defparam \line_buffer.mem14_physical .WRITE_MODE=3;
    defparam \line_buffer.mem14_physical .READ_MODE=3;
    defparam \line_buffer.mem14_physical .INIT_F=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem14_physical .INIT_E=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem14_physical .INIT_D=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem14_physical .INIT_C=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem14_physical .INIT_B=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem14_physical .INIT_A=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem14_physical .INIT_9=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem14_physical .INIT_8=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem14_physical .INIT_7=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem14_physical .INIT_6=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem14_physical .INIT_5=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem14_physical .INIT_4=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem14_physical .INIT_3=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    defparam \line_buffer.mem14_physical .INIT_2=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    defparam \line_buffer.mem14_physical .INIT_1=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    defparam \line_buffer.mem14_physical .INIT_0=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    SB_RAM40_4K \line_buffer.mem14_physical  (
            .RDATA({dangling_wire_52,dangling_wire_53,dangling_wire_54,dangling_wire_55,\line_buffer.n536 ,dangling_wire_56,dangling_wire_57,dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,\line_buffer.n535 ,dangling_wire_63,dangling_wire_64,dangling_wire_65}),
            .RADDR({N__12405,N__17211,N__18822,N__12693,N__12957,N__10380,N__10755,N__18123,N__18471,N__11721,N__11964}),
            .WADDR({N__15585,N__14067,N__14328,N__14577,N__14832,N__15093,N__15330,N__20352,N__13713,N__15888,N__16143}),
            .MASK({dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73,dangling_wire_74,dangling_wire_75,dangling_wire_76,dangling_wire_77,dangling_wire_78,dangling_wire_79,dangling_wire_80,dangling_wire_81}),
            .WDATA({dangling_wire_82,dangling_wire_83,dangling_wire_84,dangling_wire_85,N__8537,dangling_wire_86,dangling_wire_87,dangling_wire_88,dangling_wire_89,dangling_wire_90,dangling_wire_91,dangling_wire_92,N__8410,dangling_wire_93,dangling_wire_94,dangling_wire_95}),
            .RCLKE(),
            .RCLK(N__23251),
            .RE(N__19791),
            .WCLKE(),
            .WCLK(N__20154),
            .WE(N__16397));
    defparam \line_buffer.mem5_physical .WRITE_MODE=3;
    defparam \line_buffer.mem5_physical .READ_MODE=3;
    defparam \line_buffer.mem5_physical .INIT_F=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem5_physical .INIT_E=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem5_physical .INIT_D=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem5_physical .INIT_C=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem5_physical .INIT_B=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem5_physical .INIT_A=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem5_physical .INIT_9=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem5_physical .INIT_8=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem5_physical .INIT_7=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem5_physical .INIT_6=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem5_physical .INIT_5=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem5_physical .INIT_4=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem5_physical .INIT_3=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    defparam \line_buffer.mem5_physical .INIT_2=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    defparam \line_buffer.mem5_physical .INIT_1=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    defparam \line_buffer.mem5_physical .INIT_0=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    SB_RAM40_4K \line_buffer.mem5_physical  (
            .RDATA({dangling_wire_96,dangling_wire_97,dangling_wire_98,dangling_wire_99,\line_buffer.n546 ,dangling_wire_100,dangling_wire_101,dangling_wire_102,dangling_wire_103,dangling_wire_104,dangling_wire_105,dangling_wire_106,\line_buffer.n545 ,dangling_wire_107,dangling_wire_108,dangling_wire_109}),
            .RADDR({N__12336,N__17154,N__18753,N__12630,N__12882,N__10299,N__10710,N__18060,N__18402,N__11652,N__11895}),
            .WADDR({N__15534,N__14016,N__14259,N__14514,N__14763,N__15030,N__15267,N__20289,N__13650,N__15825,N__16092}),
            .MASK({dangling_wire_110,dangling_wire_111,dangling_wire_112,dangling_wire_113,dangling_wire_114,dangling_wire_115,dangling_wire_116,dangling_wire_117,dangling_wire_118,dangling_wire_119,dangling_wire_120,dangling_wire_121,dangling_wire_122,dangling_wire_123,dangling_wire_124,dangling_wire_125}),
            .WDATA({dangling_wire_126,dangling_wire_127,dangling_wire_128,dangling_wire_129,N__8639,dangling_wire_130,dangling_wire_131,dangling_wire_132,dangling_wire_133,dangling_wire_134,dangling_wire_135,dangling_wire_136,N__8753,dangling_wire_137,dangling_wire_138,dangling_wire_139}),
            .RCLKE(),
            .RCLK(N__22497),
            .RE(N__19705),
            .WCLKE(),
            .WCLK(N__20166),
            .WE(N__16987));
    defparam \line_buffer.mem11_physical .WRITE_MODE=3;
    defparam \line_buffer.mem11_physical .READ_MODE=3;
    defparam \line_buffer.mem11_physical .INIT_F=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem11_physical .INIT_E=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem11_physical .INIT_D=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem11_physical .INIT_C=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem11_physical .INIT_B=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem11_physical .INIT_A=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem11_physical .INIT_9=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem11_physical .INIT_8=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem11_physical .INIT_7=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem11_physical .INIT_6=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem11_physical .INIT_5=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem11_physical .INIT_4=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem11_physical .INIT_3=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem11_physical .INIT_2=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem11_physical .INIT_1=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem11_physical .INIT_0=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    SB_RAM40_4K \line_buffer.mem11_physical  (
            .RDATA({dangling_wire_140,dangling_wire_141,dangling_wire_142,dangling_wire_143,\line_buffer.n504 ,dangling_wire_144,dangling_wire_145,dangling_wire_146,dangling_wire_147,dangling_wire_148,dangling_wire_149,dangling_wire_150,\line_buffer.n503 ,dangling_wire_151,dangling_wire_152,dangling_wire_153}),
            .RADDR({N__12441,N__17247,N__18858,N__12729,N__12993,N__10416,N__10791,N__18159,N__18507,N__11757,N__12000}),
            .WADDR({N__15621,N__14103,N__14364,N__14613,N__14868,N__15129,N__15366,N__20388,N__13749,N__15924,N__16179}),
            .MASK({dangling_wire_154,dangling_wire_155,dangling_wire_156,dangling_wire_157,dangling_wire_158,dangling_wire_159,dangling_wire_160,dangling_wire_161,dangling_wire_162,dangling_wire_163,dangling_wire_164,dangling_wire_165,dangling_wire_166,dangling_wire_167,dangling_wire_168,dangling_wire_169}),
            .WDATA({dangling_wire_170,dangling_wire_171,dangling_wire_172,dangling_wire_173,N__8501,dangling_wire_174,dangling_wire_175,dangling_wire_176,dangling_wire_177,dangling_wire_178,dangling_wire_179,dangling_wire_180,N__8389,dangling_wire_181,dangling_wire_182,dangling_wire_183}),
            .RCLKE(),
            .RCLK(N__23293),
            .RE(N__19819),
            .WCLKE(),
            .WCLK(N__20146),
            .WE(N__16935));
    defparam \line_buffer.mem21_physical .WRITE_MODE=3;
    defparam \line_buffer.mem21_physical .READ_MODE=3;
    defparam \line_buffer.mem21_physical .INIT_F=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem21_physical .INIT_E=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem21_physical .INIT_D=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem21_physical .INIT_C=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem21_physical .INIT_B=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem21_physical .INIT_A=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem21_physical .INIT_9=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem21_physical .INIT_8=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem21_physical .INIT_7=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem21_physical .INIT_6=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem21_physical .INIT_5=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem21_physical .INIT_4=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem21_physical .INIT_3=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem21_physical .INIT_2=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem21_physical .INIT_1=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem21_physical .INIT_0=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    SB_RAM40_4K \line_buffer.mem21_physical  (
            .RDATA({dangling_wire_184,dangling_wire_185,dangling_wire_186,dangling_wire_187,\line_buffer.n566 ,dangling_wire_188,dangling_wire_189,dangling_wire_190,dangling_wire_191,dangling_wire_192,dangling_wire_193,dangling_wire_194,\line_buffer.n565 ,dangling_wire_195,dangling_wire_196,dangling_wire_197}),
            .RADDR({N__12309,N__17115,N__18726,N__12597,N__12861,N__10284,N__10659,N__18027,N__18375,N__11625,N__11868}),
            .WADDR({N__15489,N__13970,N__14232,N__14481,N__14736,N__14997,N__15234,N__20256,N__13617,N__15792,N__16047}),
            .MASK({dangling_wire_198,dangling_wire_199,dangling_wire_200,dangling_wire_201,dangling_wire_202,dangling_wire_203,dangling_wire_204,dangling_wire_205,dangling_wire_206,dangling_wire_207,dangling_wire_208,dangling_wire_209,dangling_wire_210,dangling_wire_211,dangling_wire_212,dangling_wire_213}),
            .WDATA({dangling_wire_214,dangling_wire_215,dangling_wire_216,dangling_wire_217,N__8321,dangling_wire_218,dangling_wire_219,dangling_wire_220,dangling_wire_221,dangling_wire_222,dangling_wire_223,dangling_wire_224,N__8221,dangling_wire_225,dangling_wire_226,dangling_wire_227}),
            .RCLKE(),
            .RCLK(N__22770),
            .RE(N__19700),
            .WCLKE(),
            .WCLK(N__20175),
            .WE(N__16638));
    defparam \line_buffer.mem12_physical .WRITE_MODE=3;
    defparam \line_buffer.mem12_physical .READ_MODE=3;
    defparam \line_buffer.mem12_physical .INIT_F=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem12_physical .INIT_E=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem12_physical .INIT_D=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem12_physical .INIT_C=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem12_physical .INIT_B=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem12_physical .INIT_A=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem12_physical .INIT_9=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem12_physical .INIT_8=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem12_physical .INIT_7=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem12_physical .INIT_6=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem12_physical .INIT_5=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem12_physical .INIT_4=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem12_physical .INIT_3=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem12_physical .INIT_2=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem12_physical .INIT_1=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem12_physical .INIT_0=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    SB_RAM40_4K \line_buffer.mem12_physical  (
            .RDATA({dangling_wire_228,dangling_wire_229,dangling_wire_230,dangling_wire_231,\line_buffer.n502 ,dangling_wire_232,dangling_wire_233,dangling_wire_234,dangling_wire_235,dangling_wire_236,dangling_wire_237,dangling_wire_238,\line_buffer.n501 ,dangling_wire_239,dangling_wire_240,dangling_wire_241}),
            .RADDR({N__12429,N__17235,N__18846,N__12717,N__12981,N__10404,N__10779,N__18147,N__18495,N__11745,N__11988}),
            .WADDR({N__15609,N__14091,N__14352,N__14601,N__14856,N__15117,N__15354,N__20376,N__13737,N__15912,N__16167}),
            .MASK({dangling_wire_242,dangling_wire_243,dangling_wire_244,dangling_wire_245,dangling_wire_246,dangling_wire_247,dangling_wire_248,dangling_wire_249,dangling_wire_250,dangling_wire_251,dangling_wire_252,dangling_wire_253,dangling_wire_254,dangling_wire_255,dangling_wire_256,dangling_wire_257}),
            .WDATA({dangling_wire_258,dangling_wire_259,dangling_wire_260,dangling_wire_261,N__8291,dangling_wire_262,dangling_wire_263,dangling_wire_264,dangling_wire_265,dangling_wire_266,dangling_wire_267,dangling_wire_268,N__8213,dangling_wire_269,dangling_wire_270,dangling_wire_271}),
            .RCLKE(),
            .RCLK(N__23279),
            .RE(N__19818),
            .WCLKE(),
            .WCLK(N__20148),
            .WE(N__16928));
    defparam \line_buffer.mem18_physical .WRITE_MODE=3;
    defparam \line_buffer.mem18_physical .READ_MODE=3;
    defparam \line_buffer.mem18_physical .INIT_F=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem18_physical .INIT_E=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem18_physical .INIT_D=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem18_physical .INIT_C=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem18_physical .INIT_B=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem18_physical .INIT_A=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem18_physical .INIT_9=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem18_physical .INIT_8=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem18_physical .INIT_7=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem18_physical .INIT_6=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem18_physical .INIT_5=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem18_physical .INIT_4=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem18_physical .INIT_3=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem18_physical .INIT_2=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem18_physical .INIT_1=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem18_physical .INIT_0=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    SB_RAM40_4K \line_buffer.mem18_physical  (
            .RDATA({dangling_wire_272,dangling_wire_273,dangling_wire_274,dangling_wire_275,\line_buffer.n445 ,dangling_wire_276,dangling_wire_277,dangling_wire_278,dangling_wire_279,dangling_wire_280,dangling_wire_281,dangling_wire_282,\line_buffer.n444 ,dangling_wire_283,dangling_wire_284,dangling_wire_285}),
            .RADDR({N__12357,N__17163,N__18774,N__12645,N__12909,N__10332,N__10707,N__18075,N__18423,N__11673,N__11916}),
            .WADDR({N__15537,N__14019,N__14280,N__14529,N__14784,N__15045,N__15282,N__20304,N__13665,N__15840,N__16095}),
            .MASK({dangling_wire_286,dangling_wire_287,dangling_wire_288,dangling_wire_289,dangling_wire_290,dangling_wire_291,dangling_wire_292,dangling_wire_293,dangling_wire_294,dangling_wire_295,dangling_wire_296,dangling_wire_297,dangling_wire_298,dangling_wire_299,dangling_wire_300,dangling_wire_301}),
            .WDATA({dangling_wire_302,dangling_wire_303,dangling_wire_304,dangling_wire_305,N__8325,dangling_wire_306,dangling_wire_307,dangling_wire_308,dangling_wire_309,dangling_wire_310,dangling_wire_311,dangling_wire_312,N__8214,dangling_wire_313,dangling_wire_314,dangling_wire_315}),
            .RCLKE(),
            .RCLK(N__23027),
            .RE(N__19723),
            .WCLKE(),
            .WCLK(N__20163),
            .WE(N__16439));
    defparam \line_buffer.mem24_physical .WRITE_MODE=3;
    defparam \line_buffer.mem24_physical .READ_MODE=3;
    defparam \line_buffer.mem24_physical .INIT_F=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem24_physical .INIT_E=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem24_physical .INIT_D=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem24_physical .INIT_C=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem24_physical .INIT_B=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem24_physical .INIT_A=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem24_physical .INIT_9=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem24_physical .INIT_8=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem24_physical .INIT_7=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem24_physical .INIT_6=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem24_physical .INIT_5=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem24_physical .INIT_4=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem24_physical .INIT_3=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem24_physical .INIT_2=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem24_physical .INIT_1=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem24_physical .INIT_0=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    SB_RAM40_4K \line_buffer.mem24_physical  (
            .RDATA({dangling_wire_316,dangling_wire_317,dangling_wire_318,dangling_wire_319,\line_buffer.n510 ,dangling_wire_320,dangling_wire_321,dangling_wire_322,dangling_wire_323,dangling_wire_324,dangling_wire_325,dangling_wire_326,\line_buffer.n509 ,dangling_wire_327,dangling_wire_328,dangling_wire_329}),
            .RADDR({N__12456,N__17274,N__18873,N__12750,N__13002,N__10419,N__10828,N__18180,N__18522,N__11772,N__12015}),
            .WADDR({N__15654,N__14136,N__14379,N__14634,N__14883,N__15150,N__15387,N__20409,N__13770,N__15945,N__16212}),
            .MASK({dangling_wire_330,dangling_wire_331,dangling_wire_332,dangling_wire_333,dangling_wire_334,dangling_wire_335,dangling_wire_336,dangling_wire_337,dangling_wire_338,dangling_wire_339,dangling_wire_340,dangling_wire_341,dangling_wire_342,dangling_wire_343,dangling_wire_344,dangling_wire_345}),
            .WDATA({dangling_wire_346,dangling_wire_347,dangling_wire_348,dangling_wire_349,N__8254,dangling_wire_350,dangling_wire_351,dangling_wire_352,dangling_wire_353,dangling_wire_354,dangling_wire_355,dangling_wire_356,N__8138,dangling_wire_357,dangling_wire_358,dangling_wire_359}),
            .RCLKE(),
            .RCLK(N__23271),
            .RE(N__19855),
            .WCLKE(),
            .WCLK(N__20138),
            .WE(N__16491));
    defparam \line_buffer.mem1_physical .WRITE_MODE=3;
    defparam \line_buffer.mem1_physical .READ_MODE=3;
    defparam \line_buffer.mem1_physical .INIT_F=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem1_physical .INIT_E=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem1_physical .INIT_D=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem1_physical .INIT_C=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem1_physical .INIT_B=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem1_physical .INIT_A=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem1_physical .INIT_9=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem1_physical .INIT_8=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem1_physical .INIT_7=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem1_physical .INIT_6=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem1_physical .INIT_5=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem1_physical .INIT_4=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem1_physical .INIT_3=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    defparam \line_buffer.mem1_physical .INIT_2=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    defparam \line_buffer.mem1_physical .INIT_1=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    defparam \line_buffer.mem1_physical .INIT_0=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    SB_RAM40_4K \line_buffer.mem1_physical  (
            .RDATA({dangling_wire_360,dangling_wire_361,dangling_wire_362,dangling_wire_363,\line_buffer.n538 ,dangling_wire_364,dangling_wire_365,dangling_wire_366,dangling_wire_367,dangling_wire_368,dangling_wire_369,dangling_wire_370,\line_buffer.n537 ,dangling_wire_371,dangling_wire_372,dangling_wire_373}),
            .RADDR({N__12465,N__17271,N__18882,N__12753,N__13015,N__10435,N__10815,N__18183,N__18531,N__11781,N__12024}),
            .WADDR({N__15645,N__14127,N__14388,N__14637,N__14892,N__15153,N__15390,N__20412,N__13773,N__15948,N__16203}),
            .MASK({dangling_wire_374,dangling_wire_375,dangling_wire_376,dangling_wire_377,dangling_wire_378,dangling_wire_379,dangling_wire_380,dangling_wire_381,dangling_wire_382,dangling_wire_383,dangling_wire_384,dangling_wire_385,dangling_wire_386,dangling_wire_387,dangling_wire_388,dangling_wire_389}),
            .WDATA({dangling_wire_390,dangling_wire_391,dangling_wire_392,dangling_wire_393,N__8593,dangling_wire_394,dangling_wire_395,dangling_wire_396,dangling_wire_397,dangling_wire_398,dangling_wire_399,dangling_wire_400,N__8712,dangling_wire_401,dangling_wire_402,dangling_wire_403}),
            .RCLKE(),
            .RCLK(N__23301),
            .RE(N__19839),
            .WCLKE(),
            .WCLK(N__20136),
            .WE(N__16396));
    defparam \line_buffer.mem15_physical .WRITE_MODE=3;
    defparam \line_buffer.mem15_physical .READ_MODE=3;
    defparam \line_buffer.mem15_physical .INIT_F=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem15_physical .INIT_E=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem15_physical .INIT_D=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem15_physical .INIT_C=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem15_physical .INIT_B=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem15_physical .INIT_A=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem15_physical .INIT_9=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem15_physical .INIT_8=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem15_physical .INIT_7=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem15_physical .INIT_6=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem15_physical .INIT_5=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem15_physical .INIT_4=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem15_physical .INIT_3=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    defparam \line_buffer.mem15_physical .INIT_2=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    defparam \line_buffer.mem15_physical .INIT_1=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    defparam \line_buffer.mem15_physical .INIT_0=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    SB_RAM40_4K \line_buffer.mem15_physical  (
            .RDATA({dangling_wire_404,dangling_wire_405,dangling_wire_406,dangling_wire_407,\line_buffer.n534 ,dangling_wire_408,dangling_wire_409,dangling_wire_410,dangling_wire_411,dangling_wire_412,dangling_wire_413,dangling_wire_414,\line_buffer.n533 ,dangling_wire_415,dangling_wire_416,dangling_wire_417}),
            .RADDR({N__12393,N__17199,N__18810,N__12681,N__12945,N__10368,N__10743,N__18111,N__18459,N__11709,N__11952}),
            .WADDR({N__15573,N__14055,N__14316,N__14565,N__14820,N__15081,N__15318,N__20340,N__13701,N__15876,N__16131}),
            .MASK({dangling_wire_418,dangling_wire_419,dangling_wire_420,dangling_wire_421,dangling_wire_422,dangling_wire_423,dangling_wire_424,dangling_wire_425,dangling_wire_426,dangling_wire_427,dangling_wire_428,dangling_wire_429,dangling_wire_430,dangling_wire_431,dangling_wire_432,dangling_wire_433}),
            .WDATA({dangling_wire_434,dangling_wire_435,dangling_wire_436,dangling_wire_437,N__8307,dangling_wire_438,dangling_wire_439,dangling_wire_440,dangling_wire_441,dangling_wire_442,dangling_wire_443,dangling_wire_444,N__8205,dangling_wire_445,dangling_wire_446,dangling_wire_447}),
            .RCLKE(),
            .RCLK(N__23200),
            .RE(N__19759),
            .WCLKE(),
            .WCLK(N__20156),
            .WE(N__16404));
    defparam \line_buffer.mem27_physical .WRITE_MODE=3;
    defparam \line_buffer.mem27_physical .READ_MODE=3;
    defparam \line_buffer.mem27_physical .INIT_F=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem27_physical .INIT_E=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem27_physical .INIT_D=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem27_physical .INIT_C=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem27_physical .INIT_B=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem27_physical .INIT_A=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem27_physical .INIT_9=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem27_physical .INIT_8=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem27_physical .INIT_7=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem27_physical .INIT_6=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem27_physical .INIT_5=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem27_physical .INIT_4=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem27_physical .INIT_3=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    defparam \line_buffer.mem27_physical .INIT_2=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    defparam \line_buffer.mem27_physical .INIT_1=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    defparam \line_buffer.mem27_physical .INIT_0=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    SB_RAM40_4K \line_buffer.mem27_physical  (
            .RDATA({dangling_wire_448,dangling_wire_449,dangling_wire_450,dangling_wire_451,\line_buffer.n542 ,dangling_wire_452,dangling_wire_453,dangling_wire_454,dangling_wire_455,dangling_wire_456,dangling_wire_457,dangling_wire_458,\line_buffer.n541 ,dangling_wire_459,dangling_wire_460,dangling_wire_461}),
            .RADDR({N__12420,N__17238,N__18837,N__12714,N__12966,N__10383,N__10794,N__18144,N__18486,N__11736,N__11979}),
            .WADDR({N__15618,N__14100,N__14343,N__14598,N__14847,N__15114,N__15351,N__20373,N__13734,N__15909,N__16176}),
            .MASK({dangling_wire_462,dangling_wire_463,dangling_wire_464,dangling_wire_465,dangling_wire_466,dangling_wire_467,dangling_wire_468,dangling_wire_469,dangling_wire_470,dangling_wire_471,dangling_wire_472,dangling_wire_473,dangling_wire_474,dangling_wire_475,dangling_wire_476,dangling_wire_477}),
            .WDATA({dangling_wire_478,dangling_wire_479,dangling_wire_480,dangling_wire_481,N__8285,dangling_wire_482,dangling_wire_483,dangling_wire_484,dangling_wire_485,dangling_wire_486,dangling_wire_487,dangling_wire_488,N__8169,dangling_wire_489,dangling_wire_490,dangling_wire_491}),
            .RCLKE(),
            .RCLK(N__23270),
            .RE(N__19829),
            .WCLKE(),
            .WCLK(N__20149),
            .WE(N__16976));
    defparam \line_buffer.mem4_physical .WRITE_MODE=3;
    defparam \line_buffer.mem4_physical .READ_MODE=3;
    defparam \line_buffer.mem4_physical .INIT_F=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem4_physical .INIT_E=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem4_physical .INIT_D=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem4_physical .INIT_C=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem4_physical .INIT_B=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem4_physical .INIT_A=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem4_physical .INIT_9=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem4_physical .INIT_8=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem4_physical .INIT_7=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem4_physical .INIT_6=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem4_physical .INIT_5=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem4_physical .INIT_4=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem4_physical .INIT_3=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem4_physical .INIT_2=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem4_physical .INIT_1=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem4_physical .INIT_0=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    SB_RAM40_4K \line_buffer.mem4_physical  (
            .RDATA({dangling_wire_492,dangling_wire_493,dangling_wire_494,dangling_wire_495,\line_buffer.n514 ,dangling_wire_496,dangling_wire_497,dangling_wire_498,dangling_wire_499,dangling_wire_500,dangling_wire_501,dangling_wire_502,\line_buffer.n513 ,dangling_wire_503,dangling_wire_504,dangling_wire_505}),
            .RADDR({N__12348,N__17166,N__18765,N__12642,N__12894,N__10311,N__10722,N__18072,N__18414,N__11664,N__11907}),
            .WADDR({N__15546,N__14028,N__14271,N__14526,N__14775,N__15042,N__15279,N__20301,N__13662,N__15837,N__16104}),
            .MASK({dangling_wire_506,dangling_wire_507,dangling_wire_508,dangling_wire_509,dangling_wire_510,dangling_wire_511,dangling_wire_512,dangling_wire_513,dangling_wire_514,dangling_wire_515,dangling_wire_516,dangling_wire_517,dangling_wire_518,dangling_wire_519,dangling_wire_520,dangling_wire_521}),
            .WDATA({dangling_wire_522,dangling_wire_523,dangling_wire_524,dangling_wire_525,N__8629,dangling_wire_526,dangling_wire_527,dangling_wire_528,dangling_wire_529,dangling_wire_530,dangling_wire_531,dangling_wire_532,N__8740,dangling_wire_533,dangling_wire_534,dangling_wire_535}),
            .RCLKE(),
            .RCLK(N__22882),
            .RE(N__19743),
            .WCLKE(),
            .WCLK(N__20164),
            .WE(N__16490));
    defparam \line_buffer.mem16_physical .WRITE_MODE=3;
    defparam \line_buffer.mem16_physical .READ_MODE=3;
    defparam \line_buffer.mem16_physical .INIT_F=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem16_physical .INIT_E=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem16_physical .INIT_D=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem16_physical .INIT_C=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem16_physical .INIT_B=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem16_physical .INIT_A=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem16_physical .INIT_9=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem16_physical .INIT_8=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem16_physical .INIT_7=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem16_physical .INIT_6=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem16_physical .INIT_5=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem16_physical .INIT_4=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem16_physical .INIT_3=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    defparam \line_buffer.mem16_physical .INIT_2=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    defparam \line_buffer.mem16_physical .INIT_1=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    defparam \line_buffer.mem16_physical .INIT_0=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    SB_RAM40_4K \line_buffer.mem16_physical  (
            .RDATA({dangling_wire_536,dangling_wire_537,dangling_wire_538,dangling_wire_539,\line_buffer.n532 ,dangling_wire_540,dangling_wire_541,dangling_wire_542,dangling_wire_543,dangling_wire_544,dangling_wire_545,dangling_wire_546,\line_buffer.n531 ,dangling_wire_547,dangling_wire_548,dangling_wire_549}),
            .RADDR({N__12381,N__17187,N__18798,N__12669,N__12933,N__10356,N__10731,N__18099,N__18447,N__11697,N__11940}),
            .WADDR({N__15561,N__14043,N__14304,N__14553,N__14808,N__15069,N__15306,N__20328,N__13689,N__15864,N__16119}),
            .MASK({dangling_wire_550,dangling_wire_551,dangling_wire_552,dangling_wire_553,dangling_wire_554,dangling_wire_555,dangling_wire_556,dangling_wire_557,dangling_wire_558,dangling_wire_559,dangling_wire_560,dangling_wire_561,dangling_wire_562,dangling_wire_563,dangling_wire_564,dangling_wire_565}),
            .WDATA({dangling_wire_566,dangling_wire_567,dangling_wire_568,dangling_wire_569,N__8088,dangling_wire_570,dangling_wire_571,dangling_wire_572,dangling_wire_573,dangling_wire_574,dangling_wire_575,dangling_wire_576,N__8862,dangling_wire_577,dangling_wire_578,dangling_wire_579}),
            .RCLKE(),
            .RCLK(N__23159),
            .RE(N__19758),
            .WCLKE(),
            .WCLK(N__20159),
            .WE(N__16405));
    defparam \line_buffer.mem30_physical .WRITE_MODE=3;
    defparam \line_buffer.mem30_physical .READ_MODE=3;
    defparam \line_buffer.mem30_physical .INIT_F=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem30_physical .INIT_E=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem30_physical .INIT_D=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem30_physical .INIT_C=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem30_physical .INIT_B=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem30_physical .INIT_A=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem30_physical .INIT_9=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem30_physical .INIT_8=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem30_physical .INIT_7=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem30_physical .INIT_6=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem30_physical .INIT_5=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem30_physical .INIT_4=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem30_physical .INIT_3=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    defparam \line_buffer.mem30_physical .INIT_2=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    defparam \line_buffer.mem30_physical .INIT_1=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    defparam \line_buffer.mem30_physical .INIT_0=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    SB_RAM40_4K \line_buffer.mem30_physical  (
            .RDATA({dangling_wire_580,dangling_wire_581,dangling_wire_582,dangling_wire_583,\line_buffer.n574 ,dangling_wire_584,dangling_wire_585,dangling_wire_586,dangling_wire_587,dangling_wire_588,dangling_wire_589,dangling_wire_590,\line_buffer.n573 ,dangling_wire_591,dangling_wire_592,dangling_wire_593}),
            .RADDR({N__12372,N__17190,N__18789,N__12666,N__12918,N__10335,N__10746,N__18096,N__18438,N__11688,N__11931}),
            .WADDR({N__15570,N__14052,N__14295,N__14550,N__14799,N__15066,N__15303,N__20325,N__13686,N__15861,N__16128}),
            .MASK({dangling_wire_594,dangling_wire_595,dangling_wire_596,dangling_wire_597,dangling_wire_598,dangling_wire_599,dangling_wire_600,dangling_wire_601,dangling_wire_602,dangling_wire_603,dangling_wire_604,dangling_wire_605,dangling_wire_606,dangling_wire_607,dangling_wire_608,dangling_wire_609}),
            .WDATA({dangling_wire_610,dangling_wire_611,dangling_wire_612,dangling_wire_613,N__8314,dangling_wire_614,dangling_wire_615,dangling_wire_616,dangling_wire_617,dangling_wire_618,dangling_wire_619,dangling_wire_620,N__8201,dangling_wire_621,dangling_wire_622,dangling_wire_623}),
            .RCLKE(),
            .RCLK(N__23152),
            .RE(N__19807),
            .WCLKE(),
            .WCLK(N__20160),
            .WE(N__16817));
    defparam \line_buffer.mem7_physical .WRITE_MODE=3;
    defparam \line_buffer.mem7_physical .READ_MODE=3;
    defparam \line_buffer.mem7_physical .INIT_F=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem7_physical .INIT_E=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem7_physical .INIT_D=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem7_physical .INIT_C=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem7_physical .INIT_B=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem7_physical .INIT_A=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem7_physical .INIT_9=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem7_physical .INIT_8=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem7_physical .INIT_7=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem7_physical .INIT_6=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem7_physical .INIT_5=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem7_physical .INIT_4=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem7_physical .INIT_3=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem7_physical .INIT_2=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem7_physical .INIT_1=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem7_physical .INIT_0=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    SB_RAM40_4K \line_buffer.mem7_physical  (
            .RDATA({dangling_wire_624,dangling_wire_625,dangling_wire_626,dangling_wire_627,\line_buffer.n441 ,dangling_wire_628,dangling_wire_629,dangling_wire_630,dangling_wire_631,dangling_wire_632,dangling_wire_633,dangling_wire_634,\line_buffer.n440 ,dangling_wire_635,dangling_wire_636,dangling_wire_637}),
            .RADDR({N__12312,N__17130,N__18729,N__12606,N__12858,N__10275,N__10686,N__18036,N__18378,N__11628,N__11871}),
            .WADDR({N__15510,N__13992,N__14235,N__14490,N__14739,N__15006,N__15243,N__20265,N__13626,N__15801,N__16068}),
            .MASK({dangling_wire_638,dangling_wire_639,dangling_wire_640,dangling_wire_641,dangling_wire_642,dangling_wire_643,dangling_wire_644,dangling_wire_645,dangling_wire_646,dangling_wire_647,dangling_wire_648,dangling_wire_649,dangling_wire_650,dangling_wire_651,dangling_wire_652,dangling_wire_653}),
            .WDATA({dangling_wire_654,dangling_wire_655,dangling_wire_656,dangling_wire_657,N__8644,dangling_wire_658,dangling_wire_659,dangling_wire_660,dangling_wire_661,dangling_wire_662,dangling_wire_663,dangling_wire_664,N__8755,dangling_wire_665,dangling_wire_666,dangling_wire_667}),
            .RCLKE(),
            .RCLK(N__22530),
            .RE(N__19718),
            .WCLKE(),
            .WCLK(N__20174),
            .WE(N__17033));
    defparam \line_buffer.mem20_physical .WRITE_MODE=3;
    defparam \line_buffer.mem20_physical .READ_MODE=3;
    defparam \line_buffer.mem20_physical .INIT_F=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem20_physical .INIT_E=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem20_physical .INIT_D=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem20_physical .INIT_C=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem20_physical .INIT_B=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem20_physical .INIT_A=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem20_physical .INIT_9=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem20_physical .INIT_8=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem20_physical .INIT_7=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem20_physical .INIT_6=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem20_physical .INIT_5=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem20_physical .INIT_4=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem20_physical .INIT_3=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem20_physical .INIT_2=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem20_physical .INIT_1=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem20_physical .INIT_0=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    SB_RAM40_4K \line_buffer.mem20_physical  (
            .RDATA({dangling_wire_668,dangling_wire_669,dangling_wire_670,dangling_wire_671,\line_buffer.n568 ,dangling_wire_672,dangling_wire_673,dangling_wire_674,dangling_wire_675,dangling_wire_676,dangling_wire_677,dangling_wire_678,\line_buffer.n567 ,dangling_wire_679,dangling_wire_680,dangling_wire_681}),
            .RADDR({N__12321,N__17127,N__18738,N__12609,N__12873,N__10296,N__10671,N__18039,N__18387,N__11637,N__11880}),
            .WADDR({N__15501,N__13983,N__14244,N__14493,N__14748,N__15009,N__15246,N__20268,N__13629,N__15804,N__16059}),
            .MASK({dangling_wire_682,dangling_wire_683,dangling_wire_684,dangling_wire_685,dangling_wire_686,dangling_wire_687,dangling_wire_688,dangling_wire_689,dangling_wire_690,dangling_wire_691,dangling_wire_692,dangling_wire_693,dangling_wire_694,dangling_wire_695,dangling_wire_696,dangling_wire_697}),
            .WDATA({dangling_wire_698,dangling_wire_699,dangling_wire_700,dangling_wire_701,N__8544,dangling_wire_702,dangling_wire_703,dangling_wire_704,dangling_wire_705,dangling_wire_706,dangling_wire_707,dangling_wire_708,N__8431,dangling_wire_709,dangling_wire_710,dangling_wire_711}),
            .RCLKE(),
            .RCLK(N__22912),
            .RE(N__19699),
            .WCLKE(),
            .WCLK(N__20173),
            .WE(N__16634));
    defparam \line_buffer.mem13_physical .WRITE_MODE=3;
    defparam \line_buffer.mem13_physical .READ_MODE=3;
    defparam \line_buffer.mem13_physical .INIT_F=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem13_physical .INIT_E=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem13_physical .INIT_D=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem13_physical .INIT_C=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem13_physical .INIT_B=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem13_physical .INIT_A=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem13_physical .INIT_9=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem13_physical .INIT_8=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem13_physical .INIT_7=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem13_physical .INIT_6=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem13_physical .INIT_5=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem13_physical .INIT_4=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem13_physical .INIT_3=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem13_physical .INIT_2=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem13_physical .INIT_1=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem13_physical .INIT_0=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    SB_RAM40_4K \line_buffer.mem13_physical  (
            .RDATA({dangling_wire_712,dangling_wire_713,dangling_wire_714,dangling_wire_715,\line_buffer.n500 ,dangling_wire_716,dangling_wire_717,dangling_wire_718,dangling_wire_719,dangling_wire_720,dangling_wire_721,dangling_wire_722,\line_buffer.n499 ,dangling_wire_723,dangling_wire_724,dangling_wire_725}),
            .RADDR({N__12417,N__17223,N__18834,N__12705,N__12969,N__10392,N__10767,N__18135,N__18483,N__11733,N__11976}),
            .WADDR({N__15597,N__14079,N__14340,N__14589,N__14844,N__15105,N__15342,N__20364,N__13725,N__15900,N__16155}),
            .MASK({dangling_wire_726,dangling_wire_727,dangling_wire_728,dangling_wire_729,dangling_wire_730,dangling_wire_731,dangling_wire_732,dangling_wire_733,dangling_wire_734,dangling_wire_735,dangling_wire_736,dangling_wire_737,dangling_wire_738,dangling_wire_739,dangling_wire_740,dangling_wire_741}),
            .WDATA({dangling_wire_742,dangling_wire_743,dangling_wire_744,dangling_wire_745,N__8057,dangling_wire_746,dangling_wire_747,dangling_wire_748,dangling_wire_749,dangling_wire_750,dangling_wire_751,dangling_wire_752,N__8855,dangling_wire_753,dangling_wire_754,dangling_wire_755}),
            .RCLKE(),
            .RCLK(N__23278),
            .RE(N__19792),
            .WCLKE(),
            .WCLK(N__20150),
            .WE(N__16908));
    defparam \line_buffer.mem19_physical .WRITE_MODE=3;
    defparam \line_buffer.mem19_physical .READ_MODE=3;
    defparam \line_buffer.mem19_physical .INIT_F=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem19_physical .INIT_E=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem19_physical .INIT_D=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem19_physical .INIT_C=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem19_physical .INIT_B=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem19_physical .INIT_A=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem19_physical .INIT_9=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem19_physical .INIT_8=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem19_physical .INIT_7=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem19_physical .INIT_6=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem19_physical .INIT_5=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem19_physical .INIT_4=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem19_physical .INIT_3=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem19_physical .INIT_2=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem19_physical .INIT_1=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem19_physical .INIT_0=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    SB_RAM40_4K \line_buffer.mem19_physical  (
            .RDATA({dangling_wire_756,dangling_wire_757,dangling_wire_758,dangling_wire_759,\line_buffer.n443 ,dangling_wire_760,dangling_wire_761,dangling_wire_762,dangling_wire_763,dangling_wire_764,dangling_wire_765,dangling_wire_766,\line_buffer.n442 ,dangling_wire_767,dangling_wire_768,dangling_wire_769}),
            .RADDR({N__12345,N__17151,N__18762,N__12633,N__12897,N__10320,N__10695,N__18063,N__18411,N__11661,N__11904}),
            .WADDR({N__15525,N__14007,N__14268,N__14517,N__14772,N__15033,N__15270,N__20292,N__13653,N__15828,N__16083}),
            .MASK({dangling_wire_770,dangling_wire_771,dangling_wire_772,dangling_wire_773,dangling_wire_774,dangling_wire_775,dangling_wire_776,dangling_wire_777,dangling_wire_778,dangling_wire_779,dangling_wire_780,dangling_wire_781,dangling_wire_782,dangling_wire_783,dangling_wire_784,dangling_wire_785}),
            .WDATA({dangling_wire_786,dangling_wire_787,dangling_wire_788,dangling_wire_789,N__8071,dangling_wire_790,dangling_wire_791,dangling_wire_792,dangling_wire_793,dangling_wire_794,dangling_wire_795,dangling_wire_796,N__8874,dangling_wire_797,dangling_wire_798,dangling_wire_799}),
            .RCLKE(),
            .RCLK(N__23026),
            .RE(N__19680),
            .WCLKE(),
            .WCLK(N__20165),
            .WE(N__16446));
    defparam \line_buffer.mem23_physical .WRITE_MODE=3;
    defparam \line_buffer.mem23_physical .READ_MODE=3;
    defparam \line_buffer.mem23_physical .INIT_F=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem23_physical .INIT_E=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem23_physical .INIT_D=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem23_physical .INIT_C=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem23_physical .INIT_B=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem23_physical .INIT_A=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem23_physical .INIT_9=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem23_physical .INIT_8=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem23_physical .INIT_7=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem23_physical .INIT_6=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem23_physical .INIT_5=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem23_physical .INIT_4=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem23_physical .INIT_3=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem23_physical .INIT_2=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem23_physical .INIT_1=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem23_physical .INIT_0=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    SB_RAM40_4K \line_buffer.mem23_physical  (
            .RDATA({dangling_wire_800,dangling_wire_801,dangling_wire_802,dangling_wire_803,\line_buffer.n512 ,dangling_wire_804,dangling_wire_805,dangling_wire_806,dangling_wire_807,dangling_wire_808,dangling_wire_809,dangling_wire_810,\line_buffer.n511 ,dangling_wire_811,dangling_wire_812,dangling_wire_813}),
            .RADDR({N__12468,N__17284,N__18885,N__12762,N__13014,N__10431,N__10834,N__18192,N__18534,N__11784,N__12027}),
            .WADDR({N__15661,N__14143,N__14391,N__14646,N__14895,N__15162,N__15399,N__20421,N__13782,N__15957,N__16219}),
            .MASK({dangling_wire_814,dangling_wire_815,dangling_wire_816,dangling_wire_817,dangling_wire_818,dangling_wire_819,dangling_wire_820,dangling_wire_821,dangling_wire_822,dangling_wire_823,dangling_wire_824,dangling_wire_825,dangling_wire_826,dangling_wire_827,dangling_wire_828,dangling_wire_829}),
            .WDATA({dangling_wire_830,dangling_wire_831,dangling_wire_832,dangling_wire_833,N__8516,dangling_wire_834,dangling_wire_835,dangling_wire_836,dangling_wire_837,dangling_wire_838,dangling_wire_839,dangling_wire_840,N__8357,dangling_wire_841,dangling_wire_842,dangling_wire_843}),
            .RCLKE(),
            .RCLK(N__23272),
            .RE(N__19704),
            .WCLKE(),
            .WCLK(N__20134),
            .WE(N__16492));
    defparam \line_buffer.mem0_physical .WRITE_MODE=3;
    defparam \line_buffer.mem0_physical .READ_MODE=3;
    defparam \line_buffer.mem0_physical .INIT_F=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem0_physical .INIT_E=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem0_physical .INIT_D=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem0_physical .INIT_C=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem0_physical .INIT_B=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem0_physical .INIT_A=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem0_physical .INIT_9=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem0_physical .INIT_8=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem0_physical .INIT_7=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem0_physical .INIT_6=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem0_physical .INIT_5=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem0_physical .INIT_4=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem0_physical .INIT_3=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem0_physical .INIT_2=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem0_physical .INIT_1=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem0_physical .INIT_0=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    SB_RAM40_4K \line_buffer.mem0_physical  (
            .RDATA({dangling_wire_844,dangling_wire_845,dangling_wire_846,dangling_wire_847,\line_buffer.n506 ,dangling_wire_848,dangling_wire_849,dangling_wire_850,dangling_wire_851,dangling_wire_852,dangling_wire_853,dangling_wire_854,\line_buffer.n505 ,dangling_wire_855,dangling_wire_856,dangling_wire_857}),
            .RADDR({N__12472,N__17283,N__18889,N__12763,N__13021,N__10441,N__10827,N__18193,N__18538,N__11788,N__12031}),
            .WADDR({N__15657,N__14139,N__14395,N__14647,N__14899,N__15163,N__15400,N__20422,N__13783,N__15958,N__16215}),
            .MASK({dangling_wire_858,dangling_wire_859,dangling_wire_860,dangling_wire_861,dangling_wire_862,dangling_wire_863,dangling_wire_864,dangling_wire_865,dangling_wire_866,dangling_wire_867,dangling_wire_868,dangling_wire_869,dangling_wire_870,dangling_wire_871,dangling_wire_872,dangling_wire_873}),
            .WDATA({dangling_wire_874,dangling_wire_875,dangling_wire_876,dangling_wire_877,N__8572,dangling_wire_878,dangling_wire_879,dangling_wire_880,dangling_wire_881,dangling_wire_882,dangling_wire_883,dangling_wire_884,N__8711,dangling_wire_885,dangling_wire_886,dangling_wire_887}),
            .RCLKE(),
            .RCLK(N__23302),
            .RE(N__19850),
            .WCLKE(),
            .WCLK(N__20132),
            .WE(N__16939));
    defparam \line_buffer.mem26_physical .WRITE_MODE=3;
    defparam \line_buffer.mem26_physical .READ_MODE=3;
    defparam \line_buffer.mem26_physical .INIT_F=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem26_physical .INIT_E=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem26_physical .INIT_D=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem26_physical .INIT_C=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem26_physical .INIT_B=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem26_physical .INIT_A=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem26_physical .INIT_9=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem26_physical .INIT_8=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem26_physical .INIT_7=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem26_physical .INIT_6=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem26_physical .INIT_5=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem26_physical .INIT_4=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem26_physical .INIT_3=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    defparam \line_buffer.mem26_physical .INIT_2=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    defparam \line_buffer.mem26_physical .INIT_1=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    defparam \line_buffer.mem26_physical .INIT_0=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    SB_RAM40_4K \line_buffer.mem26_physical  (
            .RDATA({dangling_wire_888,dangling_wire_889,dangling_wire_890,dangling_wire_891,\line_buffer.n544 ,dangling_wire_892,dangling_wire_893,dangling_wire_894,dangling_wire_895,dangling_wire_896,dangling_wire_897,dangling_wire_898,\line_buffer.n543 ,dangling_wire_899,dangling_wire_900,dangling_wire_901}),
            .RADDR({N__12432,N__17250,N__18849,N__12726,N__12978,N__10395,N__10806,N__18156,N__18498,N__11748,N__11991}),
            .WADDR({N__15630,N__14112,N__14355,N__14610,N__14859,N__15126,N__15363,N__20385,N__13746,N__15921,N__16188}),
            .MASK({dangling_wire_902,dangling_wire_903,dangling_wire_904,dangling_wire_905,dangling_wire_906,dangling_wire_907,dangling_wire_908,dangling_wire_909,dangling_wire_910,dangling_wire_911,dangling_wire_912,dangling_wire_913,dangling_wire_914,dangling_wire_915,dangling_wire_916,dangling_wire_917}),
            .WDATA({dangling_wire_918,dangling_wire_919,dangling_wire_920,dangling_wire_921,N__8500,dangling_wire_922,dangling_wire_923,dangling_wire_924,dangling_wire_925,dangling_wire_926,dangling_wire_927,dangling_wire_928,N__8382,dangling_wire_929,dangling_wire_930,dangling_wire_931}),
            .RCLKE(),
            .RCLK(N__22649),
            .RE(N__19843),
            .WCLKE(),
            .WCLK(N__20147),
            .WE(N__16986));
    defparam \line_buffer.mem3_physical .WRITE_MODE=3;
    defparam \line_buffer.mem3_physical .READ_MODE=3;
    defparam \line_buffer.mem3_physical .INIT_F=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem3_physical .INIT_E=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem3_physical .INIT_D=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem3_physical .INIT_C=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem3_physical .INIT_B=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem3_physical .INIT_A=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem3_physical .INIT_9=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem3_physical .INIT_8=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem3_physical .INIT_7=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem3_physical .INIT_6=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem3_physical .INIT_5=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem3_physical .INIT_4=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem3_physical .INIT_3=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem3_physical .INIT_2=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem3_physical .INIT_1=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem3_physical .INIT_0=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    SB_RAM40_4K \line_buffer.mem3_physical  (
            .RDATA({dangling_wire_932,dangling_wire_933,dangling_wire_934,dangling_wire_935,\line_buffer.n570 ,dangling_wire_936,dangling_wire_937,dangling_wire_938,dangling_wire_939,dangling_wire_940,dangling_wire_941,dangling_wire_942,\line_buffer.n569 ,dangling_wire_943,dangling_wire_944,dangling_wire_945}),
            .RADDR({N__12384,N__17202,N__18801,N__12678,N__12930,N__10347,N__10758,N__18108,N__18450,N__11700,N__11943}),
            .WADDR({N__15582,N__14064,N__14307,N__14562,N__14811,N__15078,N__15315,N__20337,N__13698,N__15873,N__16140}),
            .MASK({dangling_wire_946,dangling_wire_947,dangling_wire_948,dangling_wire_949,dangling_wire_950,dangling_wire_951,dangling_wire_952,dangling_wire_953,dangling_wire_954,dangling_wire_955,dangling_wire_956,dangling_wire_957,dangling_wire_958,dangling_wire_959,dangling_wire_960,dangling_wire_961}),
            .WDATA({dangling_wire_962,dangling_wire_963,dangling_wire_964,dangling_wire_965,N__8628,dangling_wire_966,dangling_wire_967,dangling_wire_968,dangling_wire_969,dangling_wire_970,dangling_wire_971,dangling_wire_972,N__8727,dangling_wire_973,dangling_wire_974,dangling_wire_975}),
            .RCLKE(),
            .RCLK(N__23078),
            .RE(N__19808),
            .WCLKE(),
            .WCLK(N__20157),
            .WE(N__16624));
    defparam \line_buffer.mem17_physical .WRITE_MODE=3;
    defparam \line_buffer.mem17_physical .READ_MODE=3;
    defparam \line_buffer.mem17_physical .INIT_F=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem17_physical .INIT_E=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem17_physical .INIT_D=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem17_physical .INIT_C=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem17_physical .INIT_B=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem17_physical .INIT_A=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem17_physical .INIT_9=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem17_physical .INIT_8=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem17_physical .INIT_7=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem17_physical .INIT_6=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem17_physical .INIT_5=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem17_physical .INIT_4=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem17_physical .INIT_3=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem17_physical .INIT_2=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem17_physical .INIT_1=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem17_physical .INIT_0=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    SB_RAM40_4K \line_buffer.mem17_physical  (
            .RDATA({dangling_wire_976,dangling_wire_977,dangling_wire_978,dangling_wire_979,\line_buffer.n447 ,dangling_wire_980,dangling_wire_981,dangling_wire_982,dangling_wire_983,dangling_wire_984,dangling_wire_985,dangling_wire_986,\line_buffer.n446 ,dangling_wire_987,dangling_wire_988,dangling_wire_989}),
            .RADDR({N__12369,N__17175,N__18786,N__12657,N__12921,N__10344,N__10719,N__18087,N__18435,N__11685,N__11928}),
            .WADDR({N__15549,N__14031,N__14292,N__14541,N__14796,N__15057,N__15294,N__20316,N__13677,N__15852,N__16107}),
            .MASK({dangling_wire_990,dangling_wire_991,dangling_wire_992,dangling_wire_993,dangling_wire_994,dangling_wire_995,dangling_wire_996,dangling_wire_997,dangling_wire_998,dangling_wire_999,dangling_wire_1000,dangling_wire_1001,dangling_wire_1002,dangling_wire_1003,dangling_wire_1004,dangling_wire_1005}),
            .WDATA({dangling_wire_1006,dangling_wire_1007,dangling_wire_1008,dangling_wire_1009,N__8532,dangling_wire_1010,dangling_wire_1011,dangling_wire_1012,dangling_wire_1013,dangling_wire_1014,dangling_wire_1015,dangling_wire_1016,N__8420,dangling_wire_1017,dangling_wire_1018,dangling_wire_1019}),
            .RCLKE(),
            .RCLK(N__23106),
            .RE(N__19724),
            .WCLKE(),
            .WCLK(N__20161),
            .WE(N__16438));
    defparam \line_buffer.mem31_physical .WRITE_MODE=3;
    defparam \line_buffer.mem31_physical .READ_MODE=3;
    defparam \line_buffer.mem31_physical .INIT_F=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem31_physical .INIT_E=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem31_physical .INIT_D=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem31_physical .INIT_C=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem31_physical .INIT_B=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem31_physical .INIT_A=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem31_physical .INIT_9=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem31_physical .INIT_8=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem31_physical .INIT_7=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem31_physical .INIT_6=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem31_physical .INIT_5=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem31_physical .INIT_4=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem31_physical .INIT_3=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    defparam \line_buffer.mem31_physical .INIT_2=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    defparam \line_buffer.mem31_physical .INIT_1=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    defparam \line_buffer.mem31_physical .INIT_0=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    SB_RAM40_4K \line_buffer.mem31_physical  (
            .RDATA({dangling_wire_1020,dangling_wire_1021,dangling_wire_1022,dangling_wire_1023,\line_buffer.n572 ,dangling_wire_1024,dangling_wire_1025,dangling_wire_1026,dangling_wire_1027,dangling_wire_1028,dangling_wire_1029,dangling_wire_1030,\line_buffer.n571 ,dangling_wire_1031,dangling_wire_1032,dangling_wire_1033}),
            .RADDR({N__12360,N__17178,N__18777,N__12654,N__12906,N__10323,N__10734,N__18084,N__18426,N__11676,N__11919}),
            .WADDR({N__15558,N__14040,N__14283,N__14538,N__14787,N__15054,N__15291,N__20313,N__13674,N__15849,N__16116}),
            .MASK({dangling_wire_1034,dangling_wire_1035,dangling_wire_1036,dangling_wire_1037,dangling_wire_1038,dangling_wire_1039,dangling_wire_1040,dangling_wire_1041,dangling_wire_1042,dangling_wire_1043,dangling_wire_1044,dangling_wire_1045,dangling_wire_1046,dangling_wire_1047,dangling_wire_1048,dangling_wire_1049}),
            .WDATA({dangling_wire_1050,dangling_wire_1051,dangling_wire_1052,dangling_wire_1053,N__8061,dangling_wire_1054,dangling_wire_1055,dangling_wire_1056,dangling_wire_1057,dangling_wire_1058,dangling_wire_1059,dangling_wire_1060,N__8840,dangling_wire_1061,dangling_wire_1062,dangling_wire_1063}),
            .RCLKE(),
            .RCLK(N__22545),
            .RE(N__19776),
            .WCLKE(),
            .WCLK(N__20162),
            .WE(N__16824));
    defparam \line_buffer.mem9_physical .INIT_0=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem9_physical .WRITE_MODE=3;
    defparam \line_buffer.mem9_physical .READ_MODE=3;
    defparam \line_buffer.mem9_physical .INIT_F=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem9_physical .INIT_E=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem9_physical .INIT_D=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem9_physical .INIT_C=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem9_physical .INIT_B=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem9_physical .INIT_A=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem9_physical .INIT_9=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem9_physical .INIT_8=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem9_physical .INIT_7=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem9_physical .INIT_6=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem9_physical .INIT_5=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem9_physical .INIT_4=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem9_physical .INIT_3=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem9_physical .INIT_2=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem9_physical .INIT_1=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    SB_RAM40_4K \line_buffer.mem9_physical  (
            .RDATA({dangling_wire_1064,dangling_wire_1065,dangling_wire_1066,dangling_wire_1067,\line_buffer.n437 ,dangling_wire_1068,dangling_wire_1069,dangling_wire_1070,dangling_wire_1071,dangling_wire_1072,dangling_wire_1073,dangling_wire_1074,\line_buffer.n436 ,dangling_wire_1075,dangling_wire_1076,dangling_wire_1077}),
            .RADDR({N__12288,N__17106,N__18705,N__12582,N__12834,N__10251,N__10662,N__18012,N__18354,N__11604,N__11847}),
            .WADDR({N__15486,N__13964,N__14211,N__14466,N__14715,N__14978,N__15219,N__20241,N__13602,N__15777,N__16044}),
            .MASK({dangling_wire_1078,dangling_wire_1079,dangling_wire_1080,dangling_wire_1081,dangling_wire_1082,dangling_wire_1083,dangling_wire_1084,dangling_wire_1085,dangling_wire_1086,dangling_wire_1087,dangling_wire_1088,dangling_wire_1089,dangling_wire_1090,dangling_wire_1091,dangling_wire_1092,dangling_wire_1093}),
            .WDATA({dangling_wire_1094,dangling_wire_1095,dangling_wire_1096,dangling_wire_1097,N__8329,dangling_wire_1098,dangling_wire_1099,dangling_wire_1100,dangling_wire_1101,dangling_wire_1102,dangling_wire_1103,dangling_wire_1104,N__8212,dangling_wire_1105,dangling_wire_1106,dangling_wire_1107}),
            .RCLKE(),
            .RCLK(N__22461),
            .RE(N__19757),
            .WCLKE(),
            .WCLK(N__20178),
            .WE(N__17041));
    defparam \line_buffer.mem29_physical .WRITE_MODE=3;
    defparam \line_buffer.mem29_physical .READ_MODE=3;
    defparam \line_buffer.mem29_physical .INIT_F=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem29_physical .INIT_E=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem29_physical .INIT_D=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem29_physical .INIT_C=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem29_physical .INIT_B=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem29_physical .INIT_A=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem29_physical .INIT_9=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem29_physical .INIT_8=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem29_physical .INIT_7=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem29_physical .INIT_6=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem29_physical .INIT_5=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem29_physical .INIT_4=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem29_physical .INIT_3=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    defparam \line_buffer.mem29_physical .INIT_2=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    defparam \line_buffer.mem29_physical .INIT_1=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    defparam \line_buffer.mem29_physical .INIT_0=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    SB_RAM40_4K \line_buffer.mem29_physical  (
            .RDATA({dangling_wire_1108,dangling_wire_1109,dangling_wire_1110,dangling_wire_1111,\line_buffer.n576 ,dangling_wire_1112,dangling_wire_1113,dangling_wire_1114,dangling_wire_1115,dangling_wire_1116,dangling_wire_1117,dangling_wire_1118,\line_buffer.n575 ,dangling_wire_1119,dangling_wire_1120,dangling_wire_1121}),
            .RADDR({N__12396,N__17214,N__18813,N__12690,N__12942,N__10359,N__10770,N__18120,N__18462,N__11712,N__11955}),
            .WADDR({N__15594,N__14076,N__14319,N__14574,N__14823,N__15090,N__15327,N__20349,N__13710,N__15885,N__16152}),
            .MASK({dangling_wire_1122,dangling_wire_1123,dangling_wire_1124,dangling_wire_1125,dangling_wire_1126,dangling_wire_1127,dangling_wire_1128,dangling_wire_1129,dangling_wire_1130,dangling_wire_1131,dangling_wire_1132,dangling_wire_1133,dangling_wire_1134,dangling_wire_1135,dangling_wire_1136,dangling_wire_1137}),
            .WDATA({dangling_wire_1138,dangling_wire_1139,dangling_wire_1140,dangling_wire_1141,N__8533,dangling_wire_1142,dangling_wire_1143,dangling_wire_1144,dangling_wire_1145,dangling_wire_1146,dangling_wire_1147,dangling_wire_1148,N__8395,dangling_wire_1149,dangling_wire_1150,dangling_wire_1151}),
            .RCLKE(),
            .RCLK(N__23202),
            .RE(N__19652),
            .WCLKE(),
            .WCLK(N__20155),
            .WE(N__16808));
    defparam \line_buffer.mem6_physical .WRITE_MODE=3;
    defparam \line_buffer.mem6_physical .READ_MODE=3;
    defparam \line_buffer.mem6_physical .INIT_F=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem6_physical .INIT_E=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem6_physical .INIT_D=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem6_physical .INIT_C=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem6_physical .INIT_B=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem6_physical .INIT_A=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem6_physical .INIT_9=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem6_physical .INIT_8=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem6_physical .INIT_7=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem6_physical .INIT_6=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem6_physical .INIT_5=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem6_physical .INIT_4=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem6_physical .INIT_3=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    defparam \line_buffer.mem6_physical .INIT_2=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    defparam \line_buffer.mem6_physical .INIT_1=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    defparam \line_buffer.mem6_physical .INIT_0=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    SB_RAM40_4K \line_buffer.mem6_physical  (
            .RDATA({dangling_wire_1152,dangling_wire_1153,dangling_wire_1154,dangling_wire_1155,\line_buffer.n578 ,dangling_wire_1156,dangling_wire_1157,dangling_wire_1158,dangling_wire_1159,dangling_wire_1160,dangling_wire_1161,dangling_wire_1162,\line_buffer.n577 ,dangling_wire_1163,dangling_wire_1164,dangling_wire_1165}),
            .RADDR({N__12324,N__17142,N__18741,N__12618,N__12870,N__10287,N__10698,N__18048,N__18390,N__11640,N__11883}),
            .WADDR({N__15522,N__14004,N__14247,N__14502,N__14751,N__15018,N__15255,N__20277,N__13638,N__15813,N__16080}),
            .MASK({dangling_wire_1166,dangling_wire_1167,dangling_wire_1168,dangling_wire_1169,dangling_wire_1170,dangling_wire_1171,dangling_wire_1172,dangling_wire_1173,dangling_wire_1174,dangling_wire_1175,dangling_wire_1176,dangling_wire_1177,dangling_wire_1178,dangling_wire_1179,dangling_wire_1180,dangling_wire_1181}),
            .WDATA({dangling_wire_1182,dangling_wire_1183,dangling_wire_1184,dangling_wire_1185,N__8640,dangling_wire_1186,dangling_wire_1187,dangling_wire_1188,dangling_wire_1189,dangling_wire_1190,dangling_wire_1191,dangling_wire_1192,N__8754,dangling_wire_1193,dangling_wire_1194,dangling_wire_1195}),
            .RCLKE(),
            .RCLK(N__22746),
            .RE(N__19602),
            .WCLKE(),
            .WCLK(N__20172),
            .WE(N__16828));
    defparam \line_buffer.mem10_physical .WRITE_MODE=3;
    defparam \line_buffer.mem10_physical .READ_MODE=3;
    defparam \line_buffer.mem10_physical .INIT_F=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem10_physical .INIT_E=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem10_physical .INIT_D=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem10_physical .INIT_C=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem10_physical .INIT_B=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem10_physical .INIT_A=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem10_physical .INIT_9=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem10_physical .INIT_8=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem10_physical .INIT_7=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem10_physical .INIT_6=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem10_physical .INIT_5=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem10_physical .INIT_4=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem10_physical .INIT_3=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem10_physical .INIT_2=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem10_physical .INIT_1=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem10_physical .INIT_0=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    SB_RAM40_4K \line_buffer.mem10_physical  (
            .RDATA({dangling_wire_1196,dangling_wire_1197,dangling_wire_1198,dangling_wire_1199,\line_buffer.n435 ,dangling_wire_1200,dangling_wire_1201,dangling_wire_1202,dangling_wire_1203,dangling_wire_1204,dangling_wire_1205,dangling_wire_1206,\line_buffer.n434 ,dangling_wire_1207,dangling_wire_1208,dangling_wire_1209}),
            .RADDR({N__12453,N__17259,N__18870,N__12741,N__13005,N__10428,N__10803,N__18171,N__18519,N__11769,N__12012}),
            .WADDR({N__15633,N__14115,N__14376,N__14625,N__14880,N__15141,N__15378,N__20400,N__13761,N__15936,N__16191}),
            .MASK({dangling_wire_1210,dangling_wire_1211,dangling_wire_1212,dangling_wire_1213,dangling_wire_1214,dangling_wire_1215,dangling_wire_1216,dangling_wire_1217,dangling_wire_1218,dangling_wire_1219,dangling_wire_1220,dangling_wire_1221,dangling_wire_1222,dangling_wire_1223,dangling_wire_1224,dangling_wire_1225}),
            .WDATA({dangling_wire_1226,dangling_wire_1227,dangling_wire_1228,dangling_wire_1229,N__8081,dangling_wire_1230,dangling_wire_1231,dangling_wire_1232,dangling_wire_1233,dangling_wire_1234,dangling_wire_1235,dangling_wire_1236,N__8841,dangling_wire_1237,dangling_wire_1238,dangling_wire_1239}),
            .RCLKE(),
            .RCLK(N__23294),
            .RE(N__19838),
            .WCLKE(),
            .WCLK(N__20140),
            .WE(N__17024));
    defparam \line_buffer.mem22_physical .INIT_0=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem22_physical .WRITE_MODE=3;
    defparam \line_buffer.mem22_physical .READ_MODE=3;
    defparam \line_buffer.mem22_physical .INIT_F=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem22_physical .INIT_E=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem22_physical .INIT_D=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem22_physical .INIT_C=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem22_physical .INIT_B=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem22_physical .INIT_A=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem22_physical .INIT_9=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem22_physical .INIT_8=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem22_physical .INIT_7=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem22_physical .INIT_6=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem22_physical .INIT_5=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem22_physical .INIT_4=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem22_physical .INIT_3=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem22_physical .INIT_2=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem22_physical .INIT_1=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    SB_RAM40_4K \line_buffer.mem22_physical  (
            .RDATA({dangling_wire_1240,dangling_wire_1241,dangling_wire_1242,dangling_wire_1243,\line_buffer.n564 ,dangling_wire_1244,dangling_wire_1245,dangling_wire_1246,dangling_wire_1247,dangling_wire_1248,dangling_wire_1249,dangling_wire_1250,\line_buffer.n563 ,dangling_wire_1251,dangling_wire_1252,dangling_wire_1253}),
            .RADDR({N__12297,N__17103,N__18714,N__12585,N__12849,N__10272,N__10647,N__18015,N__18363,N__11613,N__11856}),
            .WADDR({N__15476,N__13952,N__14220,N__14469,N__14724,N__14984,N__15222,N__20244,N__13605,N__15780,N__16035}),
            .MASK({dangling_wire_1254,dangling_wire_1255,dangling_wire_1256,dangling_wire_1257,dangling_wire_1258,dangling_wire_1259,dangling_wire_1260,dangling_wire_1261,dangling_wire_1262,dangling_wire_1263,dangling_wire_1264,dangling_wire_1265,dangling_wire_1266,dangling_wire_1267,dangling_wire_1268,dangling_wire_1269}),
            .WDATA({dangling_wire_1270,dangling_wire_1271,dangling_wire_1272,dangling_wire_1273,N__8089,dangling_wire_1274,dangling_wire_1275,dangling_wire_1276,dangling_wire_1277,dangling_wire_1278,dangling_wire_1279,dangling_wire_1280,N__8881,dangling_wire_1281,dangling_wire_1282,dangling_wire_1283}),
            .RCLKE(),
            .RCLK(N__22531),
            .RE(N__19742),
            .WCLKE(),
            .WCLK(N__20177),
            .WE(N__16639));
    defparam \line_buffer.mem25_physical .WRITE_MODE=3;
    defparam \line_buffer.mem25_physical .READ_MODE=3;
    defparam \line_buffer.mem25_physical .INIT_F=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem25_physical .INIT_E=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem25_physical .INIT_D=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem25_physical .INIT_C=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem25_physical .INIT_B=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem25_physical .INIT_A=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem25_physical .INIT_9=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem25_physical .INIT_8=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem25_physical .INIT_7=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem25_physical .INIT_6=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem25_physical .INIT_5=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem25_physical .INIT_4=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem25_physical .INIT_3=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem25_physical .INIT_2=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem25_physical .INIT_1=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem25_physical .INIT_0=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    SB_RAM40_4K \line_buffer.mem25_physical  (
            .RDATA({dangling_wire_1284,dangling_wire_1285,dangling_wire_1286,dangling_wire_1287,\line_buffer.n508 ,dangling_wire_1288,dangling_wire_1289,dangling_wire_1290,dangling_wire_1291,dangling_wire_1292,dangling_wire_1293,dangling_wire_1294,\line_buffer.n507 ,dangling_wire_1295,dangling_wire_1296,dangling_wire_1297}),
            .RADDR({N__12444,N__17262,N__18861,N__12738,N__12990,N__10407,N__10818,N__18168,N__18510,N__11760,N__12003}),
            .WADDR({N__15642,N__14124,N__14367,N__14622,N__14871,N__15138,N__15375,N__20397,N__13758,N__15933,N__16200}),
            .MASK({dangling_wire_1298,dangling_wire_1299,dangling_wire_1300,dangling_wire_1301,dangling_wire_1302,dangling_wire_1303,dangling_wire_1304,dangling_wire_1305,dangling_wire_1306,dangling_wire_1307,dangling_wire_1308,dangling_wire_1309,dangling_wire_1310,dangling_wire_1311,dangling_wire_1312,dangling_wire_1313}),
            .WDATA({dangling_wire_1314,dangling_wire_1315,dangling_wire_1316,dangling_wire_1317,N__8056,dangling_wire_1318,dangling_wire_1319,dangling_wire_1320,dangling_wire_1321,dangling_wire_1322,dangling_wire_1323,dangling_wire_1324,N__8809,dangling_wire_1325,dangling_wire_1326,dangling_wire_1327}),
            .RCLKE(),
            .RCLK(N__23235),
            .RE(N__19851),
            .WCLKE(),
            .WCLK(N__20144),
            .WE(N__16483));
    defparam \line_buffer.mem8_physical .WRITE_MODE=3;
    defparam \line_buffer.mem8_physical .READ_MODE=3;
    defparam \line_buffer.mem8_physical .INIT_F=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem8_physical .INIT_E=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem8_physical .INIT_D=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem8_physical .INIT_C=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem8_physical .INIT_B=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem8_physical .INIT_A=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem8_physical .INIT_9=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem8_physical .INIT_8=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem8_physical .INIT_7=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem8_physical .INIT_6=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem8_physical .INIT_5=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem8_physical .INIT_4=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem8_physical .INIT_3=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem8_physical .INIT_2=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem8_physical .INIT_1=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem8_physical .INIT_0=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    SB_RAM40_4K \line_buffer.mem8_physical  (
            .RDATA({dangling_wire_1328,dangling_wire_1329,dangling_wire_1330,dangling_wire_1331,\line_buffer.n439 ,dangling_wire_1332,dangling_wire_1333,dangling_wire_1334,dangling_wire_1335,dangling_wire_1336,dangling_wire_1337,dangling_wire_1338,\line_buffer.n438 ,dangling_wire_1339,dangling_wire_1340,dangling_wire_1341}),
            .RADDR({N__12300,N__17118,N__18717,N__12594,N__12846,N__10263,N__10674,N__18024,N__18366,N__11616,N__11859}),
            .WADDR({N__15498,N__13980,N__14223,N__14478,N__14727,N__14994,N__15231,N__20253,N__13614,N__15789,N__16056}),
            .MASK({dangling_wire_1342,dangling_wire_1343,dangling_wire_1344,dangling_wire_1345,dangling_wire_1346,dangling_wire_1347,dangling_wire_1348,dangling_wire_1349,dangling_wire_1350,dangling_wire_1351,dangling_wire_1352,dangling_wire_1353,dangling_wire_1354,dangling_wire_1355,dangling_wire_1356,dangling_wire_1357}),
            .WDATA({dangling_wire_1358,dangling_wire_1359,dangling_wire_1360,dangling_wire_1361,N__8551,dangling_wire_1362,dangling_wire_1363,dangling_wire_1364,dangling_wire_1365,dangling_wire_1366,dangling_wire_1367,dangling_wire_1368,N__8430,dangling_wire_1369,dangling_wire_1370,dangling_wire_1371}),
            .RCLKE(),
            .RCLK(N__22610),
            .RE(N__19719),
            .WCLKE(),
            .WCLK(N__20176),
            .WE(N__17040));
    defparam \line_buffer.mem28_physical .WRITE_MODE=3;
    defparam \line_buffer.mem28_physical .READ_MODE=3;
    defparam \line_buffer.mem28_physical .INIT_F=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem28_physical .INIT_E=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem28_physical .INIT_D=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem28_physical .INIT_C=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem28_physical .INIT_B=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem28_physical .INIT_A=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem28_physical .INIT_9=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem28_physical .INIT_8=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem28_physical .INIT_7=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem28_physical .INIT_6=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem28_physical .INIT_5=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem28_physical .INIT_4=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem28_physical .INIT_3=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    defparam \line_buffer.mem28_physical .INIT_2=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    defparam \line_buffer.mem28_physical .INIT_1=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    defparam \line_buffer.mem28_physical .INIT_0=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    SB_RAM40_4K \line_buffer.mem28_physical  (
            .RDATA({dangling_wire_1372,dangling_wire_1373,dangling_wire_1374,dangling_wire_1375,\line_buffer.n540 ,dangling_wire_1376,dangling_wire_1377,dangling_wire_1378,dangling_wire_1379,dangling_wire_1380,dangling_wire_1381,dangling_wire_1382,\line_buffer.n539 ,dangling_wire_1383,dangling_wire_1384,dangling_wire_1385}),
            .RADDR({N__12408,N__17226,N__18825,N__12702,N__12954,N__10371,N__10782,N__18132,N__18474,N__11724,N__11967}),
            .WADDR({N__15606,N__14088,N__14331,N__14586,N__14835,N__15102,N__15339,N__20361,N__13722,N__15897,N__16164}),
            .MASK({dangling_wire_1386,dangling_wire_1387,dangling_wire_1388,dangling_wire_1389,dangling_wire_1390,dangling_wire_1391,dangling_wire_1392,dangling_wire_1393,dangling_wire_1394,dangling_wire_1395,dangling_wire_1396,dangling_wire_1397,dangling_wire_1398,dangling_wire_1399,dangling_wire_1400,dangling_wire_1401}),
            .WDATA({dangling_wire_1402,dangling_wire_1403,dangling_wire_1404,dangling_wire_1405,N__8037,dangling_wire_1406,dangling_wire_1407,dangling_wire_1408,dangling_wire_1409,dangling_wire_1410,dangling_wire_1411,dangling_wire_1412,N__8822,dangling_wire_1413,dangling_wire_1414,dangling_wire_1415}),
            .RCLKE(),
            .RCLK(N__23269),
            .RE(N__19809),
            .WCLKE(),
            .WCLK(N__20151),
            .WE(N__16972));
    PRE_IO_GBUF TVP_CLK_pad_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__24119),
            .GLOBALBUFFEROUTPUT(TVP_CLK_c));
    defparam TVP_CLK_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_CLK_pad_iopad.PULLUP=1'b1;
    IO_PAD TVP_CLK_pad_iopad (
            .OE(N__24121),
            .DIN(N__24120),
            .DOUT(N__24119),
            .PACKAGEPIN(TVP_CLK));
    defparam TVP_CLK_pad_preio.PIN_TYPE=6'b000001;
    defparam TVP_CLK_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_CLK_pad_preio (
            .PADOEN(N__24121),
            .PADOUT(N__24120),
            .PADIN(N__24119),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_CLK_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_CLK_pad_iopad.PULLUP=1'b0;
    IO_PAD ADV_CLK_pad_iopad (
            .OE(N__24110),
            .DIN(N__24109),
            .DOUT(N__24108),
            .PACKAGEPIN(ADV_CLK));
    defparam ADV_CLK_pad_preio.PIN_TYPE=6'b011001;
    defparam ADV_CLK_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_CLK_pad_preio (
            .PADOEN(N__24110),
            .PADOUT(N__24109),
            .PADIN(N__24108),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__22632),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_3_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_3_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_3_iopad (
            .OE(N__24101),
            .DIN(N__24100),
            .DOUT(N__24099),
            .PACKAGEPIN(DEBUG[3]));
    defparam DEBUG_pad_3_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_3_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_3_preio (
            .PADOEN(N__24101),
            .PADOUT(N__24100),
            .PADIN(N__24099),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_VIDEO_pad_2_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_VIDEO_pad_2_iopad.PULLUP=1'b1;
    IO_PAD TVP_VIDEO_pad_2_iopad (
            .OE(N__24092),
            .DIN(N__24091),
            .DOUT(N__24090),
            .PACKAGEPIN(TVP_VIDEO[2]));
    defparam TVP_VIDEO_pad_2_preio.PIN_TYPE=6'b000001;
    defparam TVP_VIDEO_pad_2_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_VIDEO_pad_2_preio (
            .PADOEN(N__24092),
            .PADOUT(N__24091),
            .PADIN(N__24090),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_VIDEO_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_5_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_5_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_5_iopad (
            .OE(N__24083),
            .DIN(N__24082),
            .DOUT(N__24081),
            .PACKAGEPIN(ADV_G[5]));
    defparam ADV_G_pad_5_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_5_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_5_preio (
            .PADOEN(N__24083),
            .PADOUT(N__24082),
            .PADIN(N__24081),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__19905),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_3_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_3_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_3_iopad (
            .OE(N__24074),
            .DIN(N__24073),
            .DOUT(N__24072),
            .PACKAGEPIN(ADV_R[3]));
    defparam ADV_R_pad_3_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_3_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_3_preio (
            .PADOEN(N__24074),
            .PADOUT(N__24073),
            .PADIN(N__24072),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__23424),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_7_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_7_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_7_iopad (
            .OE(N__24065),
            .DIN(N__24064),
            .DOUT(N__24063),
            .PACKAGEPIN(DEBUG[7]));
    defparam DEBUG_pad_7_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_7_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_7_preio (
            .PADOEN(N__24065),
            .PADOUT(N__24064),
            .PADIN(N__24063),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_VIDEO_pad_6_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_VIDEO_pad_6_iopad.PULLUP=1'b1;
    IO_PAD TVP_VIDEO_pad_6_iopad (
            .OE(N__24056),
            .DIN(N__24055),
            .DOUT(N__24054),
            .PACKAGEPIN(TVP_VIDEO[6]));
    defparam TVP_VIDEO_pad_6_preio.PIN_TYPE=6'b000001;
    defparam TVP_VIDEO_pad_6_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_VIDEO_pad_6_preio (
            .PADOEN(N__24056),
            .PADOUT(N__24055),
            .PADIN(N__24054),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_VIDEO_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_1_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_1_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_1_iopad (
            .OE(N__24047),
            .DIN(N__24046),
            .DOUT(N__24045),
            .PACKAGEPIN(ADV_G[1]));
    defparam ADV_G_pad_1_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_1_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_1_preio (
            .PADOEN(N__24047),
            .PADOUT(N__24046),
            .PADIN(N__24045),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__21559),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_0_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_0_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_0_iopad (
            .OE(N__24038),
            .DIN(N__24037),
            .DOUT(N__24036),
            .PACKAGEPIN(ADV_R[0]));
    defparam ADV_R_pad_0_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_0_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_0_preio (
            .PADOEN(N__24038),
            .PADOUT(N__24037),
            .PADIN(N__24036),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12172),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_2_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_2_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_2_iopad (
            .OE(N__24029),
            .DIN(N__24028),
            .DOUT(N__24027),
            .PACKAGEPIN(DEBUG[2]));
    defparam DEBUG_pad_2_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_2_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_2_preio (
            .PADOEN(N__24029),
            .PADOUT(N__24028),
            .PADIN(N__24027),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_VIDEO_pad_3_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_VIDEO_pad_3_iopad.PULLUP=1'b1;
    IO_PAD TVP_VIDEO_pad_3_iopad (
            .OE(N__24020),
            .DIN(N__24019),
            .DOUT(N__24018),
            .PACKAGEPIN(TVP_VIDEO[3]));
    defparam TVP_VIDEO_pad_3_preio.PIN_TYPE=6'b000001;
    defparam TVP_VIDEO_pad_3_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_VIDEO_pad_3_preio (
            .PADOEN(N__24020),
            .PADOUT(N__24019),
            .PADIN(N__24018),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_VIDEO_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_4_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_4_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_4_iopad (
            .OE(N__24011),
            .DIN(N__24010),
            .DOUT(N__24009),
            .PACKAGEPIN(ADV_G[4]));
    defparam ADV_G_pad_4_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_4_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_4_preio (
            .PADOEN(N__24011),
            .PADOUT(N__24010),
            .PADIN(N__24009),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__17693),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_5_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_5_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_5_iopad (
            .OE(N__24002),
            .DIN(N__24001),
            .DOUT(N__24000),
            .PACKAGEPIN(ADV_R[5]));
    defparam ADV_R_pad_5_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_5_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_5_preio (
            .PADOEN(N__24002),
            .PADOUT(N__24001),
            .PADIN(N__24000),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__19898),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_VIDEO_pad_9_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_VIDEO_pad_9_iopad.PULLUP=1'b1;
    IO_PAD TVP_VIDEO_pad_9_iopad (
            .OE(N__23993),
            .DIN(N__23992),
            .DOUT(N__23991),
            .PACKAGEPIN(TVP_VIDEO[9]));
    defparam TVP_VIDEO_pad_9_preio.PIN_TYPE=6'b000001;
    defparam TVP_VIDEO_pad_9_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_VIDEO_pad_9_preio (
            .PADOEN(N__23993),
            .PADOUT(N__23992),
            .PADIN(N__23991),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_VIDEO_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_1_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_1_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_1_iopad (
            .OE(N__23984),
            .DIN(N__23983),
            .DOUT(N__23982),
            .PACKAGEPIN(DEBUG[1]));
    defparam DEBUG_pad_1_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_1_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_1_preio (
            .PADOEN(N__23984),
            .PADOUT(N__23983),
            .PADIN(N__23982),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_1_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_1_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_1_iopad (
            .OE(N__23975),
            .DIN(N__23974),
            .DOUT(N__23973),
            .PACKAGEPIN(ADV_B[1]));
    defparam ADV_B_pad_1_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_1_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_1_preio (
            .PADOEN(N__23975),
            .PADOUT(N__23974),
            .PADIN(N__23973),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__21545),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_SYNC_N_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_SYNC_N_pad_iopad.PULLUP=1'b1;
    IO_PAD ADV_SYNC_N_pad_iopad (
            .OE(N__23966),
            .DIN(N__23965),
            .DOUT(N__23964),
            .PACKAGEPIN(ADV_SYNC_N));
    defparam ADV_SYNC_N_pad_preio.PIN_TYPE=6'b011001;
    defparam ADV_SYNC_N_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_SYNC_N_pad_preio (
            .PADOEN(N__23966),
            .PADOUT(N__23965),
            .PADIN(N__23964),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_6_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_6_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_6_iopad (
            .OE(N__23957),
            .DIN(N__23956),
            .DOUT(N__23955),
            .PACKAGEPIN(ADV_B[6]));
    defparam ADV_B_pad_6_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_6_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_6_preio (
            .PADOEN(N__23957),
            .PADOUT(N__23956),
            .PADIN(N__23955),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12223),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_6_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_6_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_6_iopad (
            .OE(N__23948),
            .DIN(N__23947),
            .DOUT(N__23946),
            .PACKAGEPIN(DEBUG[6]));
    defparam DEBUG_pad_6_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_6_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_6_preio (
            .PADOEN(N__23948),
            .PADOUT(N__23947),
            .PADIN(N__23946),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_VIDEO_pad_7_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_VIDEO_pad_7_iopad.PULLUP=1'b1;
    IO_PAD TVP_VIDEO_pad_7_iopad (
            .OE(N__23939),
            .DIN(N__23938),
            .DOUT(N__23937),
            .PACKAGEPIN(TVP_VIDEO[7]));
    defparam TVP_VIDEO_pad_7_preio.PIN_TYPE=6'b000001;
    defparam TVP_VIDEO_pad_7_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_VIDEO_pad_7_preio (
            .PADOEN(N__23939),
            .PADOUT(N__23938),
            .PADIN(N__23937),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_VIDEO_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_0_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_0_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_0_iopad (
            .OE(N__23930),
            .DIN(N__23929),
            .DOUT(N__23928),
            .PACKAGEPIN(ADV_G[0]));
    defparam ADV_G_pad_0_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_0_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_0_preio (
            .PADOEN(N__23930),
            .PADOUT(N__23929),
            .PADIN(N__23928),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12167),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_1_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_1_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_1_iopad (
            .OE(N__23921),
            .DIN(N__23920),
            .DOUT(N__23919),
            .PACKAGEPIN(ADV_R[1]));
    defparam ADV_R_pad_1_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_1_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_1_preio (
            .PADOEN(N__23921),
            .PADOUT(N__23920),
            .PADIN(N__23919),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__21558),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_5_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_5_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_5_iopad (
            .OE(N__23912),
            .DIN(N__23911),
            .DOUT(N__23910),
            .PACKAGEPIN(DEBUG[5]));
    defparam DEBUG_pad_5_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_5_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_5_preio (
            .PADOEN(N__23912),
            .PADOUT(N__23911),
            .PADIN(N__23910),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_HSYNC_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_HSYNC_pad_iopad.PULLUP=1'b1;
    IO_PAD TVP_HSYNC_pad_iopad (
            .OE(N__23903),
            .DIN(N__23902),
            .DOUT(N__23901),
            .PACKAGEPIN(TVP_HSYNC));
    defparam TVP_HSYNC_pad_preio.PIN_TYPE=6'b000001;
    defparam TVP_HSYNC_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_HSYNC_pad_preio (
            .PADOEN(N__23903),
            .PADOUT(N__23902),
            .PADIN(N__23901),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_HSYNC_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_7_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_7_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_7_iopad (
            .OE(N__23894),
            .DIN(N__23893),
            .DOUT(N__23892),
            .PACKAGEPIN(ADV_G[7]));
    defparam ADV_G_pad_7_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_7_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_7_preio (
            .PADOEN(N__23894),
            .PADOUT(N__23893),
            .PADIN(N__23892),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__23357),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_6_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_6_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_6_iopad (
            .OE(N__23885),
            .DIN(N__23884),
            .DOUT(N__23883),
            .PACKAGEPIN(ADV_R[6]));
    defparam ADV_R_pad_6_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_6_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_6_preio (
            .PADOEN(N__23885),
            .PADOUT(N__23884),
            .PADIN(N__23883),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12215),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_VSYNC_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_VSYNC_pad_iopad.PULLUP=1'b1;
    IO_PAD TVP_VSYNC_pad_iopad (
            .OE(N__23876),
            .DIN(N__23875),
            .DOUT(N__23874),
            .PACKAGEPIN(TVP_VSYNC));
    defparam TVP_VSYNC_pad_preio.PIN_TYPE=6'b000001;
    defparam TVP_VSYNC_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_VSYNC_pad_preio (
            .PADOEN(N__23876),
            .PADOUT(N__23875),
            .PADIN(N__23874),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_VSYNC_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_BLANK_N_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_BLANK_N_pad_iopad.PULLUP=1'b1;
    IO_PAD ADV_BLANK_N_pad_iopad (
            .OE(N__23867),
            .DIN(N__23866),
            .DOUT(N__23865),
            .PACKAGEPIN(ADV_BLANK_N));
    defparam ADV_BLANK_N_pad_preio.PIN_TYPE=6'b011001;
    defparam ADV_BLANK_N_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_BLANK_N_pad_preio (
            .PADOEN(N__23867),
            .PADOUT(N__23866),
            .PADIN(N__23865),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__19657),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_0_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_0_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_0_iopad (
            .OE(N__23858),
            .DIN(N__23857),
            .DOUT(N__23856),
            .PACKAGEPIN(DEBUG[0]));
    defparam DEBUG_pad_0_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_0_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_0_preio (
            .PADOEN(N__23858),
            .PADOUT(N__23857),
            .PADIN(N__23856),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_2_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_2_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_2_iopad (
            .OE(N__23849),
            .DIN(N__23848),
            .DOUT(N__23847),
            .PACKAGEPIN(ADV_B[2]));
    defparam ADV_B_pad_2_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_2_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_2_preio (
            .PADOEN(N__23849),
            .PADOUT(N__23848),
            .PADIN(N__23847),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__17624),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_7_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_7_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_7_iopad (
            .OE(N__23840),
            .DIN(N__23839),
            .DOUT(N__23838),
            .PACKAGEPIN(ADV_B[7]));
    defparam ADV_B_pad_7_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_7_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_7_preio (
            .PADOEN(N__23840),
            .PADOUT(N__23839),
            .PADIN(N__23838),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__23364),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam LED_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam LED_pad_iopad.PULLUP=1'b1;
    IO_PAD LED_pad_iopad (
            .OE(N__23831),
            .DIN(N__23830),
            .DOUT(N__23829),
            .PACKAGEPIN(LED));
    defparam LED_pad_preio.PIN_TYPE=6'b011001;
    defparam LED_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO LED_pad_preio (
            .PADOEN(N__23831),
            .PADOUT(N__23830),
            .PADIN(N__23829),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12553),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_VIDEO_pad_4_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_VIDEO_pad_4_iopad.PULLUP=1'b1;
    IO_PAD TVP_VIDEO_pad_4_iopad (
            .OE(N__23822),
            .DIN(N__23821),
            .DOUT(N__23820),
            .PACKAGEPIN(TVP_VIDEO[4]));
    defparam TVP_VIDEO_pad_4_preio.PIN_TYPE=6'b000001;
    defparam TVP_VIDEO_pad_4_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_VIDEO_pad_4_preio (
            .PADOEN(N__23822),
            .PADOUT(N__23821),
            .PADIN(N__23820),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_VIDEO_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_3_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_3_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_3_iopad (
            .OE(N__23813),
            .DIN(N__23812),
            .DOUT(N__23811),
            .PACKAGEPIN(ADV_G[3]));
    defparam ADV_G_pad_3_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_3_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_3_preio (
            .PADOEN(N__23813),
            .PADOUT(N__23812),
            .PADIN(N__23811),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__23434),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_HSYNC_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_HSYNC_pad_iopad.PULLUP=1'b0;
    IO_PAD ADV_HSYNC_pad_iopad (
            .OE(N__23804),
            .DIN(N__23803),
            .DOUT(N__23802),
            .PACKAGEPIN(ADV_HSYNC));
    defparam ADV_HSYNC_pad_preio.PIN_TYPE=6'b011001;
    defparam ADV_HSYNC_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_HSYNC_pad_preio (
            .PADOEN(N__23804),
            .PADOUT(N__23803),
            .PADIN(N__23802),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10570),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_2_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_2_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_2_iopad (
            .OE(N__23795),
            .DIN(N__23794),
            .DOUT(N__23793),
            .PACKAGEPIN(ADV_R[2]));
    defparam ADV_R_pad_2_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_2_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_2_preio (
            .PADOEN(N__23795),
            .PADOUT(N__23794),
            .PADIN(N__23793),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__17629),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_4_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_4_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_4_iopad (
            .OE(N__23786),
            .DIN(N__23785),
            .DOUT(N__23784),
            .PACKAGEPIN(ADV_B[4]));
    defparam ADV_B_pad_4_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_4_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_4_preio (
            .PADOEN(N__23786),
            .PADOUT(N__23785),
            .PADIN(N__23784),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__17697),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_4_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_4_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_4_iopad (
            .OE(N__23777),
            .DIN(N__23776),
            .DOUT(N__23775),
            .PACKAGEPIN(DEBUG[4]));
    defparam DEBUG_pad_4_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_4_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_4_preio (
            .PADOEN(N__23777),
            .PADOUT(N__23776),
            .PADIN(N__23775),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_6_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_6_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_6_iopad (
            .OE(N__23768),
            .DIN(N__23767),
            .DOUT(N__23766),
            .PACKAGEPIN(ADV_G[6]));
    defparam ADV_G_pad_6_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_6_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_6_preio (
            .PADOEN(N__23768),
            .PADOUT(N__23767),
            .PADIN(N__23766),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12219),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_7_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_7_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_7_iopad (
            .OE(N__23759),
            .DIN(N__23758),
            .DOUT(N__23757),
            .PACKAGEPIN(ADV_R[7]));
    defparam ADV_R_pad_7_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_7_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_7_preio (
            .PADOEN(N__23759),
            .PADOUT(N__23758),
            .PADIN(N__23757),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__23365),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_3_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_3_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_3_iopad (
            .OE(N__23750),
            .DIN(N__23749),
            .DOUT(N__23748),
            .PACKAGEPIN(ADV_B[3]));
    defparam ADV_B_pad_3_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_3_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_3_preio (
            .PADOEN(N__23750),
            .PADOUT(N__23749),
            .PADIN(N__23748),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__23417),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_4_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_4_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_4_iopad (
            .OE(N__23741),
            .DIN(N__23740),
            .DOUT(N__23739),
            .PACKAGEPIN(ADV_R[4]));
    defparam ADV_R_pad_4_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_4_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_4_preio (
            .PADOEN(N__23741),
            .PADOUT(N__23740),
            .PADIN(N__23739),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__17698),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_VIDEO_pad_8_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_VIDEO_pad_8_iopad.PULLUP=1'b1;
    IO_PAD TVP_VIDEO_pad_8_iopad (
            .OE(N__23732),
            .DIN(N__23731),
            .DOUT(N__23730),
            .PACKAGEPIN(TVP_VIDEO[8]));
    defparam TVP_VIDEO_pad_8_preio.PIN_TYPE=6'b000001;
    defparam TVP_VIDEO_pad_8_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_VIDEO_pad_8_preio (
            .PADOEN(N__23732),
            .PADOUT(N__23731),
            .PADIN(N__23730),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_VIDEO_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_0_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_0_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_0_iopad (
            .OE(N__23723),
            .DIN(N__23722),
            .DOUT(N__23721),
            .PACKAGEPIN(ADV_B[0]));
    defparam ADV_B_pad_0_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_0_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_0_preio (
            .PADOEN(N__23723),
            .PADOUT(N__23722),
            .PADIN(N__23721),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12168),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_VIDEO_pad_5_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_VIDEO_pad_5_iopad.PULLUP=1'b1;
    IO_PAD TVP_VIDEO_pad_5_iopad (
            .OE(N__23714),
            .DIN(N__23713),
            .DOUT(N__23712),
            .PACKAGEPIN(TVP_VIDEO[5]));
    defparam TVP_VIDEO_pad_5_preio.PIN_TYPE=6'b000001;
    defparam TVP_VIDEO_pad_5_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_VIDEO_pad_5_preio (
            .PADOEN(N__23714),
            .PADOUT(N__23713),
            .PADIN(N__23712),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_VIDEO_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_2_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_2_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_2_iopad (
            .OE(N__23705),
            .DIN(N__23704),
            .DOUT(N__23703),
            .PACKAGEPIN(ADV_G[2]));
    defparam ADV_G_pad_2_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_2_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_2_preio (
            .PADOEN(N__23705),
            .PADOUT(N__23704),
            .PADIN(N__23703),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__17628),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_VSYNC_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_VSYNC_pad_iopad.PULLUP=1'b0;
    IO_PAD ADV_VSYNC_pad_iopad (
            .OE(N__23696),
            .DIN(N__23695),
            .DOUT(N__23694),
            .PACKAGEPIN(ADV_VSYNC));
    defparam ADV_VSYNC_pad_preio.PIN_TYPE=6'b011001;
    defparam ADV_VSYNC_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_VSYNC_pad_preio (
            .PADOEN(N__23696),
            .PADOUT(N__23695),
            .PADIN(N__23694),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__21352),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_5_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_5_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_5_iopad (
            .OE(N__23687),
            .DIN(N__23686),
            .DOUT(N__23685),
            .PACKAGEPIN(ADV_B[5]));
    defparam ADV_B_pad_5_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_5_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_5_preio (
            .PADOEN(N__23687),
            .PADOUT(N__23686),
            .PADIN(N__23685),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__19909),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__5727 (
            .O(N__23668),
            .I(N__23660));
    InMux I__5726 (
            .O(N__23667),
            .I(N__23656));
    CascadeMux I__5725 (
            .O(N__23666),
            .I(N__23650));
    InMux I__5724 (
            .O(N__23665),
            .I(N__23644));
    InMux I__5723 (
            .O(N__23664),
            .I(N__23641));
    InMux I__5722 (
            .O(N__23663),
            .I(N__23634));
    LocalMux I__5721 (
            .O(N__23660),
            .I(N__23631));
    InMux I__5720 (
            .O(N__23659),
            .I(N__23626));
    LocalMux I__5719 (
            .O(N__23656),
            .I(N__23623));
    InMux I__5718 (
            .O(N__23655),
            .I(N__23620));
    InMux I__5717 (
            .O(N__23654),
            .I(N__23617));
    InMux I__5716 (
            .O(N__23653),
            .I(N__23614));
    InMux I__5715 (
            .O(N__23650),
            .I(N__23609));
    InMux I__5714 (
            .O(N__23649),
            .I(N__23609));
    InMux I__5713 (
            .O(N__23648),
            .I(N__23606));
    InMux I__5712 (
            .O(N__23647),
            .I(N__23603));
    LocalMux I__5711 (
            .O(N__23644),
            .I(N__23596));
    LocalMux I__5710 (
            .O(N__23641),
            .I(N__23596));
    InMux I__5709 (
            .O(N__23640),
            .I(N__23593));
    InMux I__5708 (
            .O(N__23639),
            .I(N__23590));
    InMux I__5707 (
            .O(N__23638),
            .I(N__23587));
    InMux I__5706 (
            .O(N__23637),
            .I(N__23584));
    LocalMux I__5705 (
            .O(N__23634),
            .I(N__23581));
    Span4Mux_h I__5704 (
            .O(N__23631),
            .I(N__23578));
    InMux I__5703 (
            .O(N__23630),
            .I(N__23575));
    InMux I__5702 (
            .O(N__23629),
            .I(N__23571));
    LocalMux I__5701 (
            .O(N__23626),
            .I(N__23564));
    Span4Mux_h I__5700 (
            .O(N__23623),
            .I(N__23564));
    LocalMux I__5699 (
            .O(N__23620),
            .I(N__23564));
    LocalMux I__5698 (
            .O(N__23617),
            .I(N__23561));
    LocalMux I__5697 (
            .O(N__23614),
            .I(N__23554));
    LocalMux I__5696 (
            .O(N__23609),
            .I(N__23554));
    LocalMux I__5695 (
            .O(N__23606),
            .I(N__23554));
    LocalMux I__5694 (
            .O(N__23603),
            .I(N__23551));
    InMux I__5693 (
            .O(N__23602),
            .I(N__23548));
    InMux I__5692 (
            .O(N__23601),
            .I(N__23545));
    Span4Mux_h I__5691 (
            .O(N__23596),
            .I(N__23536));
    LocalMux I__5690 (
            .O(N__23593),
            .I(N__23536));
    LocalMux I__5689 (
            .O(N__23590),
            .I(N__23536));
    LocalMux I__5688 (
            .O(N__23587),
            .I(N__23529));
    LocalMux I__5687 (
            .O(N__23584),
            .I(N__23529));
    Span4Mux_h I__5686 (
            .O(N__23581),
            .I(N__23529));
    Span4Mux_v I__5685 (
            .O(N__23578),
            .I(N__23524));
    LocalMux I__5684 (
            .O(N__23575),
            .I(N__23524));
    InMux I__5683 (
            .O(N__23574),
            .I(N__23521));
    LocalMux I__5682 (
            .O(N__23571),
            .I(N__23516));
    Span4Mux_v I__5681 (
            .O(N__23564),
            .I(N__23516));
    Span4Mux_v I__5680 (
            .O(N__23561),
            .I(N__23507));
    Span4Mux_v I__5679 (
            .O(N__23554),
            .I(N__23507));
    Span4Mux_v I__5678 (
            .O(N__23551),
            .I(N__23507));
    LocalMux I__5677 (
            .O(N__23548),
            .I(N__23507));
    LocalMux I__5676 (
            .O(N__23545),
            .I(N__23504));
    InMux I__5675 (
            .O(N__23544),
            .I(N__23501));
    InMux I__5674 (
            .O(N__23543),
            .I(N__23498));
    Span4Mux_v I__5673 (
            .O(N__23536),
            .I(N__23489));
    Span4Mux_v I__5672 (
            .O(N__23529),
            .I(N__23489));
    Span4Mux_v I__5671 (
            .O(N__23524),
            .I(N__23489));
    LocalMux I__5670 (
            .O(N__23521),
            .I(N__23489));
    Span4Mux_v I__5669 (
            .O(N__23516),
            .I(N__23484));
    Span4Mux_h I__5668 (
            .O(N__23507),
            .I(N__23484));
    Odrv4 I__5667 (
            .O(N__23504),
            .I(TX_ADDR_11));
    LocalMux I__5666 (
            .O(N__23501),
            .I(TX_ADDR_11));
    LocalMux I__5665 (
            .O(N__23498),
            .I(TX_ADDR_11));
    Odrv4 I__5664 (
            .O(N__23489),
            .I(TX_ADDR_11));
    Odrv4 I__5663 (
            .O(N__23484),
            .I(TX_ADDR_11));
    InMux I__5662 (
            .O(N__23473),
            .I(N__23470));
    LocalMux I__5661 (
            .O(N__23470),
            .I(N__23467));
    Span12Mux_v I__5660 (
            .O(N__23467),
            .I(N__23464));
    Span12Mux_h I__5659 (
            .O(N__23464),
            .I(N__23461));
    Odrv12 I__5658 (
            .O(N__23461),
            .I(\line_buffer.n546 ));
    InMux I__5657 (
            .O(N__23458),
            .I(N__23455));
    LocalMux I__5656 (
            .O(N__23455),
            .I(N__23452));
    Span12Mux_h I__5655 (
            .O(N__23452),
            .I(N__23449));
    Span12Mux_v I__5654 (
            .O(N__23449),
            .I(N__23446));
    Odrv12 I__5653 (
            .O(N__23446),
            .I(\line_buffer.n538 ));
    InMux I__5652 (
            .O(N__23443),
            .I(N__23440));
    LocalMux I__5651 (
            .O(N__23440),
            .I(N__23437));
    Odrv4 I__5650 (
            .O(N__23437),
            .I(TX_DATA_3));
    IoInMux I__5649 (
            .O(N__23434),
            .I(N__23431));
    LocalMux I__5648 (
            .O(N__23431),
            .I(N__23428));
    IoSpan4Mux I__5647 (
            .O(N__23428),
            .I(N__23425));
    IoSpan4Mux I__5646 (
            .O(N__23425),
            .I(N__23421));
    IoInMux I__5645 (
            .O(N__23424),
            .I(N__23418));
    IoSpan4Mux I__5644 (
            .O(N__23421),
            .I(N__23412));
    LocalMux I__5643 (
            .O(N__23418),
            .I(N__23412));
    IoInMux I__5642 (
            .O(N__23417),
            .I(N__23409));
    Span4Mux_s3_h I__5641 (
            .O(N__23412),
            .I(N__23406));
    LocalMux I__5640 (
            .O(N__23409),
            .I(N__23403));
    Span4Mux_h I__5639 (
            .O(N__23406),
            .I(N__23400));
    IoSpan4Mux I__5638 (
            .O(N__23403),
            .I(N__23397));
    Span4Mux_h I__5637 (
            .O(N__23400),
            .I(N__23394));
    IoSpan4Mux I__5636 (
            .O(N__23397),
            .I(N__23391));
    Span4Mux_h I__5635 (
            .O(N__23394),
            .I(N__23388));
    Span4Mux_s2_v I__5634 (
            .O(N__23391),
            .I(N__23385));
    Span4Mux_h I__5633 (
            .O(N__23388),
            .I(N__23382));
    Sp12to4 I__5632 (
            .O(N__23385),
            .I(N__23379));
    Odrv4 I__5631 (
            .O(N__23382),
            .I(n1795));
    Odrv12 I__5630 (
            .O(N__23379),
            .I(n1795));
    InMux I__5629 (
            .O(N__23374),
            .I(N__23371));
    LocalMux I__5628 (
            .O(N__23371),
            .I(N__23368));
    Odrv12 I__5627 (
            .O(N__23368),
            .I(TX_DATA_7));
    IoInMux I__5626 (
            .O(N__23365),
            .I(N__23361));
    IoInMux I__5625 (
            .O(N__23364),
            .I(N__23358));
    LocalMux I__5624 (
            .O(N__23361),
            .I(N__23354));
    LocalMux I__5623 (
            .O(N__23358),
            .I(N__23351));
    IoInMux I__5622 (
            .O(N__23357),
            .I(N__23348));
    Span4Mux_s2_h I__5621 (
            .O(N__23354),
            .I(N__23345));
    Span4Mux_s2_v I__5620 (
            .O(N__23351),
            .I(N__23342));
    LocalMux I__5619 (
            .O(N__23348),
            .I(N__23339));
    Span4Mux_v I__5618 (
            .O(N__23345),
            .I(N__23336));
    Span4Mux_h I__5617 (
            .O(N__23342),
            .I(N__23333));
    IoSpan4Mux I__5616 (
            .O(N__23339),
            .I(N__23330));
    Span4Mux_v I__5615 (
            .O(N__23336),
            .I(N__23327));
    Span4Mux_v I__5614 (
            .O(N__23333),
            .I(N__23324));
    Span4Mux_s3_v I__5613 (
            .O(N__23330),
            .I(N__23321));
    Sp12to4 I__5612 (
            .O(N__23327),
            .I(N__23318));
    Span4Mux_v I__5611 (
            .O(N__23324),
            .I(N__23315));
    Sp12to4 I__5610 (
            .O(N__23321),
            .I(N__23312));
    Span12Mux_h I__5609 (
            .O(N__23318),
            .I(N__23305));
    Sp12to4 I__5608 (
            .O(N__23315),
            .I(N__23305));
    Span12Mux_s10_v I__5607 (
            .O(N__23312),
            .I(N__23305));
    Odrv12 I__5606 (
            .O(N__23305),
            .I(ADV_B_c));
    ClkMux I__5605 (
            .O(N__23302),
            .I(N__23298));
    ClkMux I__5604 (
            .O(N__23301),
            .I(N__23295));
    LocalMux I__5603 (
            .O(N__23298),
            .I(N__23289));
    LocalMux I__5602 (
            .O(N__23295),
            .I(N__23286));
    ClkMux I__5601 (
            .O(N__23294),
            .I(N__23283));
    ClkMux I__5600 (
            .O(N__23293),
            .I(N__23280));
    ClkMux I__5599 (
            .O(N__23292),
            .I(N__23275));
    Span4Mux_s2_v I__5598 (
            .O(N__23289),
            .I(N__23261));
    Span4Mux_h I__5597 (
            .O(N__23286),
            .I(N__23261));
    LocalMux I__5596 (
            .O(N__23283),
            .I(N__23261));
    LocalMux I__5595 (
            .O(N__23280),
            .I(N__23258));
    ClkMux I__5594 (
            .O(N__23279),
            .I(N__23255));
    ClkMux I__5593 (
            .O(N__23278),
            .I(N__23252));
    LocalMux I__5592 (
            .O(N__23275),
            .I(N__23248));
    ClkMux I__5591 (
            .O(N__23274),
            .I(N__23245));
    ClkMux I__5590 (
            .O(N__23273),
            .I(N__23242));
    ClkMux I__5589 (
            .O(N__23272),
            .I(N__23239));
    ClkMux I__5588 (
            .O(N__23271),
            .I(N__23236));
    ClkMux I__5587 (
            .O(N__23270),
            .I(N__23232));
    ClkMux I__5586 (
            .O(N__23269),
            .I(N__23229));
    ClkMux I__5585 (
            .O(N__23268),
            .I(N__23226));
    Span4Mux_v I__5584 (
            .O(N__23261),
            .I(N__23217));
    Span4Mux_h I__5583 (
            .O(N__23258),
            .I(N__23217));
    LocalMux I__5582 (
            .O(N__23255),
            .I(N__23217));
    LocalMux I__5581 (
            .O(N__23252),
            .I(N__23214));
    ClkMux I__5580 (
            .O(N__23251),
            .I(N__23211));
    Span4Mux_h I__5579 (
            .O(N__23248),
            .I(N__23204));
    LocalMux I__5578 (
            .O(N__23245),
            .I(N__23204));
    LocalMux I__5577 (
            .O(N__23242),
            .I(N__23204));
    LocalMux I__5576 (
            .O(N__23239),
            .I(N__23194));
    LocalMux I__5575 (
            .O(N__23236),
            .I(N__23194));
    ClkMux I__5574 (
            .O(N__23235),
            .I(N__23191));
    LocalMux I__5573 (
            .O(N__23232),
            .I(N__23182));
    LocalMux I__5572 (
            .O(N__23229),
            .I(N__23182));
    LocalMux I__5571 (
            .O(N__23226),
            .I(N__23182));
    ClkMux I__5570 (
            .O(N__23225),
            .I(N__23179));
    ClkMux I__5569 (
            .O(N__23224),
            .I(N__23176));
    Span4Mux_v I__5568 (
            .O(N__23217),
            .I(N__23167));
    Span4Mux_h I__5567 (
            .O(N__23214),
            .I(N__23167));
    LocalMux I__5566 (
            .O(N__23211),
            .I(N__23167));
    Span4Mux_v I__5565 (
            .O(N__23204),
            .I(N__23164));
    ClkMux I__5564 (
            .O(N__23203),
            .I(N__23161));
    ClkMux I__5563 (
            .O(N__23202),
            .I(N__23156));
    ClkMux I__5562 (
            .O(N__23201),
            .I(N__23153));
    ClkMux I__5561 (
            .O(N__23200),
            .I(N__23148));
    ClkMux I__5560 (
            .O(N__23199),
            .I(N__23145));
    Span4Mux_s3_v I__5559 (
            .O(N__23194),
            .I(N__23138));
    LocalMux I__5558 (
            .O(N__23191),
            .I(N__23138));
    ClkMux I__5557 (
            .O(N__23190),
            .I(N__23135));
    ClkMux I__5556 (
            .O(N__23189),
            .I(N__23131));
    Span4Mux_v I__5555 (
            .O(N__23182),
            .I(N__23125));
    LocalMux I__5554 (
            .O(N__23179),
            .I(N__23125));
    LocalMux I__5553 (
            .O(N__23176),
            .I(N__23122));
    ClkMux I__5552 (
            .O(N__23175),
            .I(N__23119));
    ClkMux I__5551 (
            .O(N__23174),
            .I(N__23116));
    Span4Mux_v I__5550 (
            .O(N__23167),
            .I(N__23113));
    Span4Mux_v I__5549 (
            .O(N__23164),
            .I(N__23108));
    LocalMux I__5548 (
            .O(N__23161),
            .I(N__23108));
    ClkMux I__5547 (
            .O(N__23160),
            .I(N__23102));
    ClkMux I__5546 (
            .O(N__23159),
            .I(N__23097));
    LocalMux I__5545 (
            .O(N__23156),
            .I(N__23091));
    LocalMux I__5544 (
            .O(N__23153),
            .I(N__23091));
    ClkMux I__5543 (
            .O(N__23152),
            .I(N__23088));
    ClkMux I__5542 (
            .O(N__23151),
            .I(N__23083));
    LocalMux I__5541 (
            .O(N__23148),
            .I(N__23074));
    LocalMux I__5540 (
            .O(N__23145),
            .I(N__23070));
    ClkMux I__5539 (
            .O(N__23144),
            .I(N__23067));
    ClkMux I__5538 (
            .O(N__23143),
            .I(N__23064));
    Span4Mux_v I__5537 (
            .O(N__23138),
            .I(N__23059));
    LocalMux I__5536 (
            .O(N__23135),
            .I(N__23059));
    ClkMux I__5535 (
            .O(N__23134),
            .I(N__23056));
    LocalMux I__5534 (
            .O(N__23131),
            .I(N__23052));
    ClkMux I__5533 (
            .O(N__23130),
            .I(N__23049));
    Span4Mux_v I__5532 (
            .O(N__23125),
            .I(N__23042));
    Span4Mux_h I__5531 (
            .O(N__23122),
            .I(N__23042));
    LocalMux I__5530 (
            .O(N__23119),
            .I(N__23042));
    LocalMux I__5529 (
            .O(N__23116),
            .I(N__23039));
    Span4Mux_h I__5528 (
            .O(N__23113),
            .I(N__23034));
    Span4Mux_h I__5527 (
            .O(N__23108),
            .I(N__23034));
    ClkMux I__5526 (
            .O(N__23107),
            .I(N__23031));
    ClkMux I__5525 (
            .O(N__23106),
            .I(N__23028));
    ClkMux I__5524 (
            .O(N__23105),
            .I(N__23023));
    LocalMux I__5523 (
            .O(N__23102),
            .I(N__23020));
    ClkMux I__5522 (
            .O(N__23101),
            .I(N__23017));
    ClkMux I__5521 (
            .O(N__23100),
            .I(N__23014));
    LocalMux I__5520 (
            .O(N__23097),
            .I(N__23011));
    ClkMux I__5519 (
            .O(N__23096),
            .I(N__23008));
    Span4Mux_h I__5518 (
            .O(N__23091),
            .I(N__23005));
    LocalMux I__5517 (
            .O(N__23088),
            .I(N__23002));
    ClkMux I__5516 (
            .O(N__23087),
            .I(N__22999));
    ClkMux I__5515 (
            .O(N__23086),
            .I(N__22991));
    LocalMux I__5514 (
            .O(N__23083),
            .I(N__22986));
    ClkMux I__5513 (
            .O(N__23082),
            .I(N__22983));
    ClkMux I__5512 (
            .O(N__23081),
            .I(N__22976));
    ClkMux I__5511 (
            .O(N__23080),
            .I(N__22973));
    ClkMux I__5510 (
            .O(N__23079),
            .I(N__22969));
    ClkMux I__5509 (
            .O(N__23078),
            .I(N__22965));
    ClkMux I__5508 (
            .O(N__23077),
            .I(N__22962));
    Span4Mux_h I__5507 (
            .O(N__23074),
            .I(N__22958));
    ClkMux I__5506 (
            .O(N__23073),
            .I(N__22955));
    Span4Mux_v I__5505 (
            .O(N__23070),
            .I(N__22948));
    LocalMux I__5504 (
            .O(N__23067),
            .I(N__22948));
    LocalMux I__5503 (
            .O(N__23064),
            .I(N__22948));
    Span4Mux_v I__5502 (
            .O(N__23059),
            .I(N__22942));
    LocalMux I__5501 (
            .O(N__23056),
            .I(N__22942));
    ClkMux I__5500 (
            .O(N__23055),
            .I(N__22939));
    Span4Mux_h I__5499 (
            .O(N__23052),
            .I(N__22933));
    LocalMux I__5498 (
            .O(N__23049),
            .I(N__22933));
    Span4Mux_h I__5497 (
            .O(N__23042),
            .I(N__22923));
    Span4Mux_h I__5496 (
            .O(N__23039),
            .I(N__22923));
    Span4Mux_h I__5495 (
            .O(N__23034),
            .I(N__22923));
    LocalMux I__5494 (
            .O(N__23031),
            .I(N__22923));
    LocalMux I__5493 (
            .O(N__23028),
            .I(N__22920));
    ClkMux I__5492 (
            .O(N__23027),
            .I(N__22917));
    ClkMux I__5491 (
            .O(N__23026),
            .I(N__22914));
    LocalMux I__5490 (
            .O(N__23023),
            .I(N__22909));
    Span4Mux_h I__5489 (
            .O(N__23020),
            .I(N__22902));
    LocalMux I__5488 (
            .O(N__23017),
            .I(N__22902));
    LocalMux I__5487 (
            .O(N__23014),
            .I(N__22902));
    Span4Mux_h I__5486 (
            .O(N__23011),
            .I(N__22897));
    LocalMux I__5485 (
            .O(N__23008),
            .I(N__22897));
    Span4Mux_v I__5484 (
            .O(N__23005),
            .I(N__22890));
    Span4Mux_h I__5483 (
            .O(N__23002),
            .I(N__22890));
    LocalMux I__5482 (
            .O(N__22999),
            .I(N__22890));
    ClkMux I__5481 (
            .O(N__22998),
            .I(N__22887));
    ClkMux I__5480 (
            .O(N__22997),
            .I(N__22884));
    ClkMux I__5479 (
            .O(N__22996),
            .I(N__22879));
    ClkMux I__5478 (
            .O(N__22995),
            .I(N__22876));
    ClkMux I__5477 (
            .O(N__22994),
            .I(N__22873));
    LocalMux I__5476 (
            .O(N__22991),
            .I(N__22869));
    ClkMux I__5475 (
            .O(N__22990),
            .I(N__22866));
    ClkMux I__5474 (
            .O(N__22989),
            .I(N__22863));
    Span4Mux_h I__5473 (
            .O(N__22986),
            .I(N__22858));
    LocalMux I__5472 (
            .O(N__22983),
            .I(N__22858));
    ClkMux I__5471 (
            .O(N__22982),
            .I(N__22855));
    ClkMux I__5470 (
            .O(N__22981),
            .I(N__22850));
    ClkMux I__5469 (
            .O(N__22980),
            .I(N__22847));
    ClkMux I__5468 (
            .O(N__22979),
            .I(N__22844));
    LocalMux I__5467 (
            .O(N__22976),
            .I(N__22840));
    LocalMux I__5466 (
            .O(N__22973),
            .I(N__22837));
    ClkMux I__5465 (
            .O(N__22972),
            .I(N__22834));
    LocalMux I__5464 (
            .O(N__22969),
            .I(N__22829));
    ClkMux I__5463 (
            .O(N__22968),
            .I(N__22826));
    LocalMux I__5462 (
            .O(N__22965),
            .I(N__22821));
    LocalMux I__5461 (
            .O(N__22962),
            .I(N__22818));
    ClkMux I__5460 (
            .O(N__22961),
            .I(N__22815));
    Span4Mux_h I__5459 (
            .O(N__22958),
            .I(N__22810));
    LocalMux I__5458 (
            .O(N__22955),
            .I(N__22810));
    Span4Mux_h I__5457 (
            .O(N__22948),
            .I(N__22806));
    ClkMux I__5456 (
            .O(N__22947),
            .I(N__22803));
    Span4Mux_h I__5455 (
            .O(N__22942),
            .I(N__22800));
    LocalMux I__5454 (
            .O(N__22939),
            .I(N__22797));
    ClkMux I__5453 (
            .O(N__22938),
            .I(N__22794));
    Span4Mux_h I__5452 (
            .O(N__22933),
            .I(N__22791));
    ClkMux I__5451 (
            .O(N__22932),
            .I(N__22788));
    Span4Mux_h I__5450 (
            .O(N__22923),
            .I(N__22785));
    Span4Mux_h I__5449 (
            .O(N__22920),
            .I(N__22780));
    LocalMux I__5448 (
            .O(N__22917),
            .I(N__22780));
    LocalMux I__5447 (
            .O(N__22914),
            .I(N__22777));
    ClkMux I__5446 (
            .O(N__22913),
            .I(N__22774));
    ClkMux I__5445 (
            .O(N__22912),
            .I(N__22771));
    Span4Mux_h I__5444 (
            .O(N__22909),
            .I(N__22765));
    Span4Mux_h I__5443 (
            .O(N__22902),
            .I(N__22765));
    Span4Mux_h I__5442 (
            .O(N__22897),
            .I(N__22758));
    Span4Mux_h I__5441 (
            .O(N__22890),
            .I(N__22758));
    LocalMux I__5440 (
            .O(N__22887),
            .I(N__22758));
    LocalMux I__5439 (
            .O(N__22884),
            .I(N__22755));
    ClkMux I__5438 (
            .O(N__22883),
            .I(N__22752));
    ClkMux I__5437 (
            .O(N__22882),
            .I(N__22748));
    LocalMux I__5436 (
            .O(N__22879),
            .I(N__22743));
    LocalMux I__5435 (
            .O(N__22876),
            .I(N__22738));
    LocalMux I__5434 (
            .O(N__22873),
            .I(N__22738));
    ClkMux I__5433 (
            .O(N__22872),
            .I(N__22735));
    Span4Mux_v I__5432 (
            .O(N__22869),
            .I(N__22728));
    LocalMux I__5431 (
            .O(N__22866),
            .I(N__22728));
    LocalMux I__5430 (
            .O(N__22863),
            .I(N__22728));
    Span4Mux_h I__5429 (
            .O(N__22858),
            .I(N__22723));
    LocalMux I__5428 (
            .O(N__22855),
            .I(N__22723));
    ClkMux I__5427 (
            .O(N__22854),
            .I(N__22720));
    ClkMux I__5426 (
            .O(N__22853),
            .I(N__22717));
    LocalMux I__5425 (
            .O(N__22850),
            .I(N__22714));
    LocalMux I__5424 (
            .O(N__22847),
            .I(N__22711));
    LocalMux I__5423 (
            .O(N__22844),
            .I(N__22708));
    ClkMux I__5422 (
            .O(N__22843),
            .I(N__22705));
    Span4Mux_v I__5421 (
            .O(N__22840),
            .I(N__22698));
    Span4Mux_h I__5420 (
            .O(N__22837),
            .I(N__22698));
    LocalMux I__5419 (
            .O(N__22834),
            .I(N__22698));
    ClkMux I__5418 (
            .O(N__22833),
            .I(N__22695));
    ClkMux I__5417 (
            .O(N__22832),
            .I(N__22691));
    Span4Mux_v I__5416 (
            .O(N__22829),
            .I(N__22685));
    LocalMux I__5415 (
            .O(N__22826),
            .I(N__22685));
    ClkMux I__5414 (
            .O(N__22825),
            .I(N__22682));
    ClkMux I__5413 (
            .O(N__22824),
            .I(N__22679));
    Span4Mux_h I__5412 (
            .O(N__22821),
            .I(N__22670));
    Span4Mux_v I__5411 (
            .O(N__22818),
            .I(N__22670));
    LocalMux I__5410 (
            .O(N__22815),
            .I(N__22670));
    Span4Mux_h I__5409 (
            .O(N__22810),
            .I(N__22670));
    ClkMux I__5408 (
            .O(N__22809),
            .I(N__22667));
    Span4Mux_v I__5407 (
            .O(N__22806),
            .I(N__22662));
    LocalMux I__5406 (
            .O(N__22803),
            .I(N__22662));
    Span4Mux_v I__5405 (
            .O(N__22800),
            .I(N__22651));
    Span4Mux_h I__5404 (
            .O(N__22797),
            .I(N__22651));
    LocalMux I__5403 (
            .O(N__22794),
            .I(N__22651));
    Span4Mux_h I__5402 (
            .O(N__22791),
            .I(N__22651));
    LocalMux I__5401 (
            .O(N__22788),
            .I(N__22651));
    Span4Mux_v I__5400 (
            .O(N__22785),
            .I(N__22646));
    Span4Mux_v I__5399 (
            .O(N__22780),
            .I(N__22639));
    Span4Mux_h I__5398 (
            .O(N__22777),
            .I(N__22639));
    LocalMux I__5397 (
            .O(N__22774),
            .I(N__22639));
    LocalMux I__5396 (
            .O(N__22771),
            .I(N__22636));
    ClkMux I__5395 (
            .O(N__22770),
            .I(N__22633));
    Span4Mux_v I__5394 (
            .O(N__22765),
            .I(N__22623));
    Span4Mux_h I__5393 (
            .O(N__22758),
            .I(N__22623));
    Span4Mux_v I__5392 (
            .O(N__22755),
            .I(N__22623));
    LocalMux I__5391 (
            .O(N__22752),
            .I(N__22623));
    ClkMux I__5390 (
            .O(N__22751),
            .I(N__22620));
    LocalMux I__5389 (
            .O(N__22748),
            .I(N__22617));
    ClkMux I__5388 (
            .O(N__22747),
            .I(N__22614));
    ClkMux I__5387 (
            .O(N__22746),
            .I(N__22611));
    Span4Mux_h I__5386 (
            .O(N__22743),
            .I(N__22603));
    Span4Mux_h I__5385 (
            .O(N__22738),
            .I(N__22603));
    LocalMux I__5384 (
            .O(N__22735),
            .I(N__22603));
    Span4Mux_h I__5383 (
            .O(N__22728),
            .I(N__22594));
    Span4Mux_v I__5382 (
            .O(N__22723),
            .I(N__22594));
    LocalMux I__5381 (
            .O(N__22720),
            .I(N__22594));
    LocalMux I__5380 (
            .O(N__22717),
            .I(N__22594));
    Span4Mux_h I__5379 (
            .O(N__22714),
            .I(N__22585));
    Span4Mux_v I__5378 (
            .O(N__22711),
            .I(N__22585));
    Span4Mux_h I__5377 (
            .O(N__22708),
            .I(N__22585));
    LocalMux I__5376 (
            .O(N__22705),
            .I(N__22585));
    Span4Mux_v I__5375 (
            .O(N__22698),
            .I(N__22580));
    LocalMux I__5374 (
            .O(N__22695),
            .I(N__22580));
    ClkMux I__5373 (
            .O(N__22694),
            .I(N__22577));
    LocalMux I__5372 (
            .O(N__22691),
            .I(N__22574));
    ClkMux I__5371 (
            .O(N__22690),
            .I(N__22571));
    Span4Mux_h I__5370 (
            .O(N__22685),
            .I(N__22566));
    LocalMux I__5369 (
            .O(N__22682),
            .I(N__22566));
    LocalMux I__5368 (
            .O(N__22679),
            .I(N__22559));
    Span4Mux_h I__5367 (
            .O(N__22670),
            .I(N__22559));
    LocalMux I__5366 (
            .O(N__22667),
            .I(N__22559));
    Span4Mux_h I__5365 (
            .O(N__22662),
            .I(N__22552));
    Span4Mux_h I__5364 (
            .O(N__22651),
            .I(N__22552));
    ClkMux I__5363 (
            .O(N__22650),
            .I(N__22549));
    ClkMux I__5362 (
            .O(N__22649),
            .I(N__22546));
    Span4Mux_v I__5361 (
            .O(N__22646),
            .I(N__22542));
    Span4Mux_v I__5360 (
            .O(N__22639),
            .I(N__22535));
    Span4Mux_h I__5359 (
            .O(N__22636),
            .I(N__22535));
    LocalMux I__5358 (
            .O(N__22633),
            .I(N__22535));
    IoInMux I__5357 (
            .O(N__22632),
            .I(N__22532));
    Span4Mux_v I__5356 (
            .O(N__22623),
            .I(N__22525));
    LocalMux I__5355 (
            .O(N__22620),
            .I(N__22525));
    Span4Mux_h I__5354 (
            .O(N__22617),
            .I(N__22520));
    LocalMux I__5353 (
            .O(N__22614),
            .I(N__22520));
    LocalMux I__5352 (
            .O(N__22611),
            .I(N__22517));
    ClkMux I__5351 (
            .O(N__22610),
            .I(N__22514));
    Span4Mux_v I__5350 (
            .O(N__22603),
            .I(N__22503));
    Span4Mux_v I__5349 (
            .O(N__22594),
            .I(N__22503));
    Span4Mux_h I__5348 (
            .O(N__22585),
            .I(N__22503));
    Span4Mux_h I__5347 (
            .O(N__22580),
            .I(N__22503));
    LocalMux I__5346 (
            .O(N__22577),
            .I(N__22503));
    Span4Mux_h I__5345 (
            .O(N__22574),
            .I(N__22498));
    LocalMux I__5344 (
            .O(N__22571),
            .I(N__22498));
    Span4Mux_v I__5343 (
            .O(N__22566),
            .I(N__22492));
    Span4Mux_h I__5342 (
            .O(N__22559),
            .I(N__22492));
    ClkMux I__5341 (
            .O(N__22558),
            .I(N__22489));
    ClkMux I__5340 (
            .O(N__22557),
            .I(N__22486));
    Span4Mux_v I__5339 (
            .O(N__22552),
            .I(N__22483));
    LocalMux I__5338 (
            .O(N__22549),
            .I(N__22480));
    LocalMux I__5337 (
            .O(N__22546),
            .I(N__22477));
    ClkMux I__5336 (
            .O(N__22545),
            .I(N__22474));
    Span4Mux_v I__5335 (
            .O(N__22542),
            .I(N__22471));
    Span4Mux_v I__5334 (
            .O(N__22535),
            .I(N__22468));
    LocalMux I__5333 (
            .O(N__22532),
            .I(N__22465));
    ClkMux I__5332 (
            .O(N__22531),
            .I(N__22462));
    ClkMux I__5331 (
            .O(N__22530),
            .I(N__22458));
    Span4Mux_h I__5330 (
            .O(N__22525),
            .I(N__22453));
    Span4Mux_h I__5329 (
            .O(N__22520),
            .I(N__22453));
    Span4Mux_h I__5328 (
            .O(N__22517),
            .I(N__22450));
    LocalMux I__5327 (
            .O(N__22514),
            .I(N__22447));
    Span4Mux_v I__5326 (
            .O(N__22503),
            .I(N__22442));
    Span4Mux_h I__5325 (
            .O(N__22498),
            .I(N__22442));
    ClkMux I__5324 (
            .O(N__22497),
            .I(N__22439));
    Span4Mux_v I__5323 (
            .O(N__22492),
            .I(N__22434));
    LocalMux I__5322 (
            .O(N__22489),
            .I(N__22434));
    LocalMux I__5321 (
            .O(N__22486),
            .I(N__22431));
    Span4Mux_v I__5320 (
            .O(N__22483),
            .I(N__22426));
    Span4Mux_h I__5319 (
            .O(N__22480),
            .I(N__22426));
    Span12Mux_h I__5318 (
            .O(N__22477),
            .I(N__22423));
    LocalMux I__5317 (
            .O(N__22474),
            .I(N__22420));
    Span4Mux_v I__5316 (
            .O(N__22471),
            .I(N__22415));
    Span4Mux_h I__5315 (
            .O(N__22468),
            .I(N__22415));
    Span4Mux_s1_v I__5314 (
            .O(N__22465),
            .I(N__22412));
    LocalMux I__5313 (
            .O(N__22462),
            .I(N__22409));
    ClkMux I__5312 (
            .O(N__22461),
            .I(N__22406));
    LocalMux I__5311 (
            .O(N__22458),
            .I(N__22403));
    Span4Mux_v I__5310 (
            .O(N__22453),
            .I(N__22400));
    Span4Mux_v I__5309 (
            .O(N__22450),
            .I(N__22395));
    Span4Mux_h I__5308 (
            .O(N__22447),
            .I(N__22395));
    Span4Mux_v I__5307 (
            .O(N__22442),
            .I(N__22392));
    LocalMux I__5306 (
            .O(N__22439),
            .I(N__22389));
    Span4Mux_v I__5305 (
            .O(N__22434),
            .I(N__22384));
    Span4Mux_h I__5304 (
            .O(N__22431),
            .I(N__22384));
    Span4Mux_v I__5303 (
            .O(N__22426),
            .I(N__22381));
    Span12Mux_v I__5302 (
            .O(N__22423),
            .I(N__22376));
    Span12Mux_h I__5301 (
            .O(N__22420),
            .I(N__22376));
    Sp12to4 I__5300 (
            .O(N__22415),
            .I(N__22369));
    Sp12to4 I__5299 (
            .O(N__22412),
            .I(N__22369));
    Sp12to4 I__5298 (
            .O(N__22409),
            .I(N__22369));
    LocalMux I__5297 (
            .O(N__22406),
            .I(N__22366));
    Span12Mux_h I__5296 (
            .O(N__22403),
            .I(N__22363));
    Span4Mux_v I__5295 (
            .O(N__22400),
            .I(N__22358));
    Span4Mux_h I__5294 (
            .O(N__22395),
            .I(N__22358));
    Span4Mux_v I__5293 (
            .O(N__22392),
            .I(N__22355));
    Span12Mux_h I__5292 (
            .O(N__22389),
            .I(N__22350));
    Sp12to4 I__5291 (
            .O(N__22384),
            .I(N__22350));
    Span4Mux_v I__5290 (
            .O(N__22381),
            .I(N__22347));
    Span12Mux_v I__5289 (
            .O(N__22376),
            .I(N__22340));
    Span12Mux_h I__5288 (
            .O(N__22369),
            .I(N__22340));
    Span12Mux_h I__5287 (
            .O(N__22366),
            .I(N__22340));
    Odrv12 I__5286 (
            .O(N__22363),
            .I(ADV_CLK_c));
    Odrv4 I__5285 (
            .O(N__22358),
            .I(ADV_CLK_c));
    Odrv4 I__5284 (
            .O(N__22355),
            .I(ADV_CLK_c));
    Odrv12 I__5283 (
            .O(N__22350),
            .I(ADV_CLK_c));
    Odrv4 I__5282 (
            .O(N__22347),
            .I(ADV_CLK_c));
    Odrv12 I__5281 (
            .O(N__22340),
            .I(ADV_CLK_c));
    SRMux I__5280 (
            .O(N__22327),
            .I(N__22323));
    SRMux I__5279 (
            .O(N__22326),
            .I(N__22316));
    LocalMux I__5278 (
            .O(N__22323),
            .I(N__22312));
    SRMux I__5277 (
            .O(N__22322),
            .I(N__22309));
    SRMux I__5276 (
            .O(N__22321),
            .I(N__22306));
    SRMux I__5275 (
            .O(N__22320),
            .I(N__22303));
    SRMux I__5274 (
            .O(N__22319),
            .I(N__22300));
    LocalMux I__5273 (
            .O(N__22316),
            .I(N__22297));
    SRMux I__5272 (
            .O(N__22315),
            .I(N__22294));
    Span4Mux_v I__5271 (
            .O(N__22312),
            .I(N__22289));
    LocalMux I__5270 (
            .O(N__22309),
            .I(N__22289));
    LocalMux I__5269 (
            .O(N__22306),
            .I(N__22286));
    LocalMux I__5268 (
            .O(N__22303),
            .I(N__22283));
    LocalMux I__5267 (
            .O(N__22300),
            .I(N__22280));
    Span4Mux_h I__5266 (
            .O(N__22297),
            .I(N__22275));
    LocalMux I__5265 (
            .O(N__22294),
            .I(N__22275));
    Span4Mux_h I__5264 (
            .O(N__22289),
            .I(N__22272));
    Span4Mux_v I__5263 (
            .O(N__22286),
            .I(N__22267));
    Span4Mux_v I__5262 (
            .O(N__22283),
            .I(N__22267));
    Span4Mux_h I__5261 (
            .O(N__22280),
            .I(N__22264));
    Span4Mux_h I__5260 (
            .O(N__22275),
            .I(N__22261));
    Odrv4 I__5259 (
            .O(N__22272),
            .I(\transmit_module.n2354 ));
    Odrv4 I__5258 (
            .O(N__22267),
            .I(\transmit_module.n2354 ));
    Odrv4 I__5257 (
            .O(N__22264),
            .I(\transmit_module.n2354 ));
    Odrv4 I__5256 (
            .O(N__22261),
            .I(\transmit_module.n2354 ));
    InMux I__5255 (
            .O(N__22252),
            .I(N__22249));
    LocalMux I__5254 (
            .O(N__22249),
            .I(N__22246));
    Span4Mux_v I__5253 (
            .O(N__22246),
            .I(N__22243));
    Span4Mux_h I__5252 (
            .O(N__22243),
            .I(N__22240));
    Odrv4 I__5251 (
            .O(N__22240),
            .I(\line_buffer.n449 ));
    CascadeMux I__5250 (
            .O(N__22237),
            .I(N__22228));
    CascadeMux I__5249 (
            .O(N__22236),
            .I(N__22222));
    CascadeMux I__5248 (
            .O(N__22235),
            .I(N__22219));
    InMux I__5247 (
            .O(N__22234),
            .I(N__22212));
    CascadeMux I__5246 (
            .O(N__22233),
            .I(N__22209));
    CascadeMux I__5245 (
            .O(N__22232),
            .I(N__22206));
    InMux I__5244 (
            .O(N__22231),
            .I(N__22203));
    InMux I__5243 (
            .O(N__22228),
            .I(N__22200));
    InMux I__5242 (
            .O(N__22227),
            .I(N__22190));
    InMux I__5241 (
            .O(N__22226),
            .I(N__22190));
    InMux I__5240 (
            .O(N__22225),
            .I(N__22190));
    InMux I__5239 (
            .O(N__22222),
            .I(N__22190));
    InMux I__5238 (
            .O(N__22219),
            .I(N__22187));
    CascadeMux I__5237 (
            .O(N__22218),
            .I(N__22183));
    CascadeMux I__5236 (
            .O(N__22217),
            .I(N__22180));
    CascadeMux I__5235 (
            .O(N__22216),
            .I(N__22175));
    InMux I__5234 (
            .O(N__22215),
            .I(N__22169));
    LocalMux I__5233 (
            .O(N__22212),
            .I(N__22166));
    InMux I__5232 (
            .O(N__22209),
            .I(N__22163));
    InMux I__5231 (
            .O(N__22206),
            .I(N__22160));
    LocalMux I__5230 (
            .O(N__22203),
            .I(N__22155));
    LocalMux I__5229 (
            .O(N__22200),
            .I(N__22155));
    InMux I__5228 (
            .O(N__22199),
            .I(N__22152));
    LocalMux I__5227 (
            .O(N__22190),
            .I(N__22149));
    LocalMux I__5226 (
            .O(N__22187),
            .I(N__22146));
    InMux I__5225 (
            .O(N__22186),
            .I(N__22143));
    InMux I__5224 (
            .O(N__22183),
            .I(N__22140));
    InMux I__5223 (
            .O(N__22180),
            .I(N__22137));
    InMux I__5222 (
            .O(N__22179),
            .I(N__22134));
    InMux I__5221 (
            .O(N__22178),
            .I(N__22129));
    InMux I__5220 (
            .O(N__22175),
            .I(N__22129));
    CascadeMux I__5219 (
            .O(N__22174),
            .I(N__22126));
    InMux I__5218 (
            .O(N__22173),
            .I(N__22119));
    InMux I__5217 (
            .O(N__22172),
            .I(N__22116));
    LocalMux I__5216 (
            .O(N__22169),
            .I(N__22107));
    Span4Mux_v I__5215 (
            .O(N__22166),
            .I(N__22107));
    LocalMux I__5214 (
            .O(N__22163),
            .I(N__22107));
    LocalMux I__5213 (
            .O(N__22160),
            .I(N__22107));
    Span4Mux_v I__5212 (
            .O(N__22155),
            .I(N__22104));
    LocalMux I__5211 (
            .O(N__22152),
            .I(N__22097));
    Span4Mux_v I__5210 (
            .O(N__22149),
            .I(N__22097));
    Span4Mux_v I__5209 (
            .O(N__22146),
            .I(N__22097));
    LocalMux I__5208 (
            .O(N__22143),
            .I(N__22092));
    LocalMux I__5207 (
            .O(N__22140),
            .I(N__22092));
    LocalMux I__5206 (
            .O(N__22137),
            .I(N__22089));
    LocalMux I__5205 (
            .O(N__22134),
            .I(N__22086));
    LocalMux I__5204 (
            .O(N__22129),
            .I(N__22083));
    InMux I__5203 (
            .O(N__22126),
            .I(N__22080));
    InMux I__5202 (
            .O(N__22125),
            .I(N__22077));
    InMux I__5201 (
            .O(N__22124),
            .I(N__22074));
    InMux I__5200 (
            .O(N__22123),
            .I(N__22069));
    InMux I__5199 (
            .O(N__22122),
            .I(N__22069));
    LocalMux I__5198 (
            .O(N__22119),
            .I(N__22066));
    LocalMux I__5197 (
            .O(N__22116),
            .I(N__22057));
    Span4Mux_v I__5196 (
            .O(N__22107),
            .I(N__22057));
    Span4Mux_h I__5195 (
            .O(N__22104),
            .I(N__22057));
    Span4Mux_h I__5194 (
            .O(N__22097),
            .I(N__22057));
    Span4Mux_v I__5193 (
            .O(N__22092),
            .I(N__22052));
    Span4Mux_v I__5192 (
            .O(N__22089),
            .I(N__22052));
    Span4Mux_v I__5191 (
            .O(N__22086),
            .I(N__22045));
    Span4Mux_v I__5190 (
            .O(N__22083),
            .I(N__22045));
    LocalMux I__5189 (
            .O(N__22080),
            .I(N__22045));
    LocalMux I__5188 (
            .O(N__22077),
            .I(TX_ADDR_12));
    LocalMux I__5187 (
            .O(N__22074),
            .I(TX_ADDR_12));
    LocalMux I__5186 (
            .O(N__22069),
            .I(TX_ADDR_12));
    Odrv4 I__5185 (
            .O(N__22066),
            .I(TX_ADDR_12));
    Odrv4 I__5184 (
            .O(N__22057),
            .I(TX_ADDR_12));
    Odrv4 I__5183 (
            .O(N__22052),
            .I(TX_ADDR_12));
    Odrv4 I__5182 (
            .O(N__22045),
            .I(TX_ADDR_12));
    CascadeMux I__5181 (
            .O(N__22030),
            .I(N__22027));
    InMux I__5180 (
            .O(N__22027),
            .I(N__22024));
    LocalMux I__5179 (
            .O(N__22024),
            .I(N__22021));
    Span12Mux_h I__5178 (
            .O(N__22021),
            .I(N__22018));
    Span12Mux_v I__5177 (
            .O(N__22018),
            .I(N__22015));
    Span12Mux_h I__5176 (
            .O(N__22015),
            .I(N__22012));
    Odrv12 I__5175 (
            .O(N__22012),
            .I(\line_buffer.n441 ));
    InMux I__5174 (
            .O(N__22009),
            .I(N__22006));
    LocalMux I__5173 (
            .O(N__22006),
            .I(\line_buffer.n3704 ));
    InMux I__5172 (
            .O(N__22003),
            .I(N__22000));
    LocalMux I__5171 (
            .O(N__22000),
            .I(\line_buffer.n3707 ));
    SRMux I__5170 (
            .O(N__21997),
            .I(N__21994));
    LocalMux I__5169 (
            .O(N__21994),
            .I(N__21991));
    Span4Mux_h I__5168 (
            .O(N__21991),
            .I(N__21986));
    SRMux I__5167 (
            .O(N__21990),
            .I(N__21983));
    SRMux I__5166 (
            .O(N__21989),
            .I(N__21980));
    Span4Mux_v I__5165 (
            .O(N__21986),
            .I(N__21976));
    LocalMux I__5164 (
            .O(N__21983),
            .I(N__21973));
    LocalMux I__5163 (
            .O(N__21980),
            .I(N__21970));
    SRMux I__5162 (
            .O(N__21979),
            .I(N__21967));
    Span4Mux_v I__5161 (
            .O(N__21976),
            .I(N__21962));
    Span4Mux_h I__5160 (
            .O(N__21973),
            .I(N__21962));
    Span4Mux_h I__5159 (
            .O(N__21970),
            .I(N__21957));
    LocalMux I__5158 (
            .O(N__21967),
            .I(N__21957));
    Span4Mux_v I__5157 (
            .O(N__21962),
            .I(N__21951));
    Span4Mux_h I__5156 (
            .O(N__21957),
            .I(N__21951));
    SRMux I__5155 (
            .O(N__21956),
            .I(N__21948));
    Span4Mux_v I__5154 (
            .O(N__21951),
            .I(N__21943));
    LocalMux I__5153 (
            .O(N__21948),
            .I(N__21940));
    SRMux I__5152 (
            .O(N__21947),
            .I(N__21937));
    SRMux I__5151 (
            .O(N__21946),
            .I(N__21934));
    Span4Mux_v I__5150 (
            .O(N__21943),
            .I(N__21926));
    Span4Mux_h I__5149 (
            .O(N__21940),
            .I(N__21926));
    LocalMux I__5148 (
            .O(N__21937),
            .I(N__21926));
    LocalMux I__5147 (
            .O(N__21934),
            .I(N__21923));
    SRMux I__5146 (
            .O(N__21933),
            .I(N__21920));
    Span4Mux_v I__5145 (
            .O(N__21926),
            .I(N__21917));
    Span4Mux_v I__5144 (
            .O(N__21923),
            .I(N__21914));
    LocalMux I__5143 (
            .O(N__21920),
            .I(N__21911));
    Odrv4 I__5142 (
            .O(N__21917),
            .I(\receive_module.n3793 ));
    Odrv4 I__5141 (
            .O(N__21914),
            .I(\receive_module.n3793 ));
    Odrv12 I__5140 (
            .O(N__21911),
            .I(\receive_module.n3793 ));
    InMux I__5139 (
            .O(N__21904),
            .I(N__21901));
    LocalMux I__5138 (
            .O(N__21901),
            .I(N__21898));
    Span12Mux_v I__5137 (
            .O(N__21898),
            .I(N__21895));
    Odrv12 I__5136 (
            .O(N__21895),
            .I(\line_buffer.n542 ));
    InMux I__5135 (
            .O(N__21892),
            .I(N__21889));
    LocalMux I__5134 (
            .O(N__21889),
            .I(N__21886));
    Odrv12 I__5133 (
            .O(N__21886),
            .I(\line_buffer.n534 ));
    InMux I__5132 (
            .O(N__21883),
            .I(N__21880));
    LocalMux I__5131 (
            .O(N__21880),
            .I(N__21877));
    Span4Mux_v I__5130 (
            .O(N__21877),
            .I(N__21874));
    Span4Mux_h I__5129 (
            .O(N__21874),
            .I(N__21871));
    Odrv4 I__5128 (
            .O(N__21871),
            .I(\line_buffer.n445 ));
    CascadeMux I__5127 (
            .O(N__21868),
            .I(N__21865));
    InMux I__5126 (
            .O(N__21865),
            .I(N__21862));
    LocalMux I__5125 (
            .O(N__21862),
            .I(N__21859));
    Span4Mux_v I__5124 (
            .O(N__21859),
            .I(N__21856));
    Span4Mux_v I__5123 (
            .O(N__21856),
            .I(N__21853));
    Sp12to4 I__5122 (
            .O(N__21853),
            .I(N__21850));
    Span12Mux_h I__5121 (
            .O(N__21850),
            .I(N__21847));
    Odrv12 I__5120 (
            .O(N__21847),
            .I(\line_buffer.n437 ));
    InMux I__5119 (
            .O(N__21844),
            .I(N__21841));
    LocalMux I__5118 (
            .O(N__21841),
            .I(\line_buffer.n3710 ));
    InMux I__5117 (
            .O(N__21838),
            .I(N__21835));
    LocalMux I__5116 (
            .O(N__21835),
            .I(N__21832));
    Span4Mux_v I__5115 (
            .O(N__21832),
            .I(N__21829));
    Span4Mux_h I__5114 (
            .O(N__21829),
            .I(N__21826));
    Sp12to4 I__5113 (
            .O(N__21826),
            .I(N__21823));
    Odrv12 I__5112 (
            .O(N__21823),
            .I(\line_buffer.n566 ));
    InMux I__5111 (
            .O(N__21820),
            .I(N__21817));
    LocalMux I__5110 (
            .O(N__21817),
            .I(N__21814));
    Sp12to4 I__5109 (
            .O(N__21814),
            .I(N__21811));
    Odrv12 I__5108 (
            .O(N__21811),
            .I(\line_buffer.n574 ));
    InMux I__5107 (
            .O(N__21808),
            .I(N__21805));
    LocalMux I__5106 (
            .O(N__21805),
            .I(N__21802));
    Span4Mux_h I__5105 (
            .O(N__21802),
            .I(N__21799));
    Span4Mux_v I__5104 (
            .O(N__21799),
            .I(N__21796));
    Span4Mux_v I__5103 (
            .O(N__21796),
            .I(N__21793));
    Odrv4 I__5102 (
            .O(N__21793),
            .I(\line_buffer.n502 ));
    InMux I__5101 (
            .O(N__21790),
            .I(N__21787));
    LocalMux I__5100 (
            .O(N__21787),
            .I(N__21784));
    Span4Mux_v I__5099 (
            .O(N__21784),
            .I(N__21781));
    Sp12to4 I__5098 (
            .O(N__21781),
            .I(N__21778));
    Span12Mux_v I__5097 (
            .O(N__21778),
            .I(N__21775));
    Odrv12 I__5096 (
            .O(N__21775),
            .I(\line_buffer.n510 ));
    CascadeMux I__5095 (
            .O(N__21772),
            .I(\line_buffer.n3758_cascade_ ));
    InMux I__5094 (
            .O(N__21769),
            .I(N__21766));
    LocalMux I__5093 (
            .O(N__21766),
            .I(N__21763));
    Span12Mux_v I__5092 (
            .O(N__21763),
            .I(N__21760));
    Odrv12 I__5091 (
            .O(N__21760),
            .I(\line_buffer.n540 ));
    InMux I__5090 (
            .O(N__21757),
            .I(N__21754));
    LocalMux I__5089 (
            .O(N__21754),
            .I(N__21751));
    Odrv12 I__5088 (
            .O(N__21751),
            .I(\line_buffer.n532 ));
    InMux I__5087 (
            .O(N__21748),
            .I(N__21745));
    LocalMux I__5086 (
            .O(N__21745),
            .I(N__21742));
    Span4Mux_h I__5085 (
            .O(N__21742),
            .I(N__21739));
    Sp12to4 I__5084 (
            .O(N__21739),
            .I(N__21736));
    Span12Mux_v I__5083 (
            .O(N__21736),
            .I(N__21733));
    Odrv12 I__5082 (
            .O(N__21733),
            .I(\line_buffer.n435 ));
    InMux I__5081 (
            .O(N__21730),
            .I(N__21727));
    LocalMux I__5080 (
            .O(N__21727),
            .I(N__21724));
    Span4Mux_v I__5079 (
            .O(N__21724),
            .I(N__21721));
    Span4Mux_h I__5078 (
            .O(N__21721),
            .I(N__21718));
    Odrv4 I__5077 (
            .O(N__21718),
            .I(\line_buffer.n443 ));
    CascadeMux I__5076 (
            .O(N__21715),
            .I(\line_buffer.n3740_cascade_ ));
    InMux I__5075 (
            .O(N__21712),
            .I(N__21709));
    LocalMux I__5074 (
            .O(N__21709),
            .I(\line_buffer.n3743 ));
    InMux I__5073 (
            .O(N__21706),
            .I(N__21703));
    LocalMux I__5072 (
            .O(N__21703),
            .I(\line_buffer.n3761 ));
    InMux I__5071 (
            .O(N__21700),
            .I(N__21697));
    LocalMux I__5070 (
            .O(N__21697),
            .I(\line_buffer.n3713 ));
    CascadeMux I__5069 (
            .O(N__21694),
            .I(N__21688));
    InMux I__5068 (
            .O(N__21693),
            .I(N__21685));
    InMux I__5067 (
            .O(N__21692),
            .I(N__21679));
    InMux I__5066 (
            .O(N__21691),
            .I(N__21676));
    InMux I__5065 (
            .O(N__21688),
            .I(N__21671));
    LocalMux I__5064 (
            .O(N__21685),
            .I(N__21668));
    InMux I__5063 (
            .O(N__21684),
            .I(N__21665));
    InMux I__5062 (
            .O(N__21683),
            .I(N__21662));
    CascadeMux I__5061 (
            .O(N__21682),
            .I(N__21658));
    LocalMux I__5060 (
            .O(N__21679),
            .I(N__21653));
    LocalMux I__5059 (
            .O(N__21676),
            .I(N__21653));
    CascadeMux I__5058 (
            .O(N__21675),
            .I(N__21649));
    CascadeMux I__5057 (
            .O(N__21674),
            .I(N__21646));
    LocalMux I__5056 (
            .O(N__21671),
            .I(N__21641));
    Span4Mux_v I__5055 (
            .O(N__21668),
            .I(N__21636));
    LocalMux I__5054 (
            .O(N__21665),
            .I(N__21636));
    LocalMux I__5053 (
            .O(N__21662),
            .I(N__21633));
    InMux I__5052 (
            .O(N__21661),
            .I(N__21628));
    InMux I__5051 (
            .O(N__21658),
            .I(N__21628));
    Span4Mux_v I__5050 (
            .O(N__21653),
            .I(N__21625));
    InMux I__5049 (
            .O(N__21652),
            .I(N__21622));
    InMux I__5048 (
            .O(N__21649),
            .I(N__21617));
    InMux I__5047 (
            .O(N__21646),
            .I(N__21617));
    InMux I__5046 (
            .O(N__21645),
            .I(N__21614));
    InMux I__5045 (
            .O(N__21644),
            .I(N__21611));
    Span4Mux_v I__5044 (
            .O(N__21641),
            .I(N__21606));
    Span4Mux_h I__5043 (
            .O(N__21636),
            .I(N__21606));
    Span12Mux_h I__5042 (
            .O(N__21633),
            .I(N__21603));
    LocalMux I__5041 (
            .O(N__21628),
            .I(N__21594));
    Span4Mux_h I__5040 (
            .O(N__21625),
            .I(N__21594));
    LocalMux I__5039 (
            .O(N__21622),
            .I(N__21594));
    LocalMux I__5038 (
            .O(N__21617),
            .I(N__21594));
    LocalMux I__5037 (
            .O(N__21614),
            .I(N__21591));
    LocalMux I__5036 (
            .O(N__21611),
            .I(TX_ADDR_13));
    Odrv4 I__5035 (
            .O(N__21606),
            .I(TX_ADDR_13));
    Odrv12 I__5034 (
            .O(N__21603),
            .I(TX_ADDR_13));
    Odrv4 I__5033 (
            .O(N__21594),
            .I(TX_ADDR_13));
    Odrv4 I__5032 (
            .O(N__21591),
            .I(TX_ADDR_13));
    InMux I__5031 (
            .O(N__21580),
            .I(N__21577));
    LocalMux I__5030 (
            .O(N__21577),
            .I(N__21574));
    Odrv12 I__5029 (
            .O(N__21574),
            .I(\line_buffer.n3767 ));
    InMux I__5028 (
            .O(N__21571),
            .I(N__21568));
    LocalMux I__5027 (
            .O(N__21568),
            .I(\transmit_module.Y_DELTA_PATTERN_15 ));
    InMux I__5026 (
            .O(N__21565),
            .I(N__21562));
    LocalMux I__5025 (
            .O(N__21562),
            .I(\transmit_module.Y_DELTA_PATTERN_14 ));
    IoInMux I__5024 (
            .O(N__21559),
            .I(N__21555));
    IoInMux I__5023 (
            .O(N__21558),
            .I(N__21552));
    LocalMux I__5022 (
            .O(N__21555),
            .I(N__21549));
    LocalMux I__5021 (
            .O(N__21552),
            .I(N__21546));
    IoSpan4Mux I__5020 (
            .O(N__21549),
            .I(N__21542));
    Span4Mux_s1_h I__5019 (
            .O(N__21546),
            .I(N__21539));
    IoInMux I__5018 (
            .O(N__21545),
            .I(N__21536));
    Span4Mux_s3_v I__5017 (
            .O(N__21542),
            .I(N__21533));
    Span4Mux_h I__5016 (
            .O(N__21539),
            .I(N__21530));
    LocalMux I__5015 (
            .O(N__21536),
            .I(N__21527));
    Sp12to4 I__5014 (
            .O(N__21533),
            .I(N__21522));
    Sp12to4 I__5013 (
            .O(N__21530),
            .I(N__21522));
    Span4Mux_s0_v I__5012 (
            .O(N__21527),
            .I(N__21519));
    Span12Mux_s11_v I__5011 (
            .O(N__21522),
            .I(N__21516));
    Span4Mux_v I__5010 (
            .O(N__21519),
            .I(N__21513));
    Span12Mux_h I__5009 (
            .O(N__21516),
            .I(N__21510));
    Span4Mux_v I__5008 (
            .O(N__21513),
            .I(N__21507));
    Odrv12 I__5007 (
            .O(N__21510),
            .I(n1797));
    Odrv4 I__5006 (
            .O(N__21507),
            .I(n1797));
    InMux I__5005 (
            .O(N__21502),
            .I(N__21499));
    LocalMux I__5004 (
            .O(N__21499),
            .I(\transmit_module.Y_DELTA_PATTERN_21 ));
    InMux I__5003 (
            .O(N__21496),
            .I(N__21493));
    LocalMux I__5002 (
            .O(N__21493),
            .I(\transmit_module.Y_DELTA_PATTERN_20 ));
    CEMux I__5001 (
            .O(N__21490),
            .I(N__21485));
    CEMux I__5000 (
            .O(N__21489),
            .I(N__21479));
    SRMux I__4999 (
            .O(N__21488),
            .I(N__21475));
    LocalMux I__4998 (
            .O(N__21485),
            .I(N__21471));
    CEMux I__4997 (
            .O(N__21484),
            .I(N__21468));
    CEMux I__4996 (
            .O(N__21483),
            .I(N__21465));
    CEMux I__4995 (
            .O(N__21482),
            .I(N__21462));
    LocalMux I__4994 (
            .O(N__21479),
            .I(N__21454));
    CEMux I__4993 (
            .O(N__21478),
            .I(N__21450));
    LocalMux I__4992 (
            .O(N__21475),
            .I(N__21446));
    SRMux I__4991 (
            .O(N__21474),
            .I(N__21443));
    Span4Mux_v I__4990 (
            .O(N__21471),
            .I(N__21438));
    LocalMux I__4989 (
            .O(N__21468),
            .I(N__21438));
    LocalMux I__4988 (
            .O(N__21465),
            .I(N__21433));
    LocalMux I__4987 (
            .O(N__21462),
            .I(N__21433));
    CEMux I__4986 (
            .O(N__21461),
            .I(N__21430));
    CEMux I__4985 (
            .O(N__21460),
            .I(N__21427));
    CEMux I__4984 (
            .O(N__21459),
            .I(N__21424));
    SRMux I__4983 (
            .O(N__21458),
            .I(N__21421));
    SRMux I__4982 (
            .O(N__21457),
            .I(N__21418));
    Span4Mux_v I__4981 (
            .O(N__21454),
            .I(N__21415));
    CEMux I__4980 (
            .O(N__21453),
            .I(N__21412));
    LocalMux I__4979 (
            .O(N__21450),
            .I(N__21409));
    CEMux I__4978 (
            .O(N__21449),
            .I(N__21406));
    Span4Mux_h I__4977 (
            .O(N__21446),
            .I(N__21403));
    LocalMux I__4976 (
            .O(N__21443),
            .I(N__21400));
    Span4Mux_v I__4975 (
            .O(N__21438),
            .I(N__21393));
    Span4Mux_v I__4974 (
            .O(N__21433),
            .I(N__21393));
    LocalMux I__4973 (
            .O(N__21430),
            .I(N__21393));
    LocalMux I__4972 (
            .O(N__21427),
            .I(N__21390));
    LocalMux I__4971 (
            .O(N__21424),
            .I(N__21387));
    LocalMux I__4970 (
            .O(N__21421),
            .I(N__21382));
    LocalMux I__4969 (
            .O(N__21418),
            .I(N__21382));
    Sp12to4 I__4968 (
            .O(N__21415),
            .I(N__21377));
    LocalMux I__4967 (
            .O(N__21412),
            .I(N__21377));
    Span4Mux_h I__4966 (
            .O(N__21409),
            .I(N__21368));
    LocalMux I__4965 (
            .O(N__21406),
            .I(N__21368));
    Span4Mux_h I__4964 (
            .O(N__21403),
            .I(N__21368));
    Span4Mux_h I__4963 (
            .O(N__21400),
            .I(N__21368));
    Span4Mux_h I__4962 (
            .O(N__21393),
            .I(N__21359));
    Span4Mux_v I__4961 (
            .O(N__21390),
            .I(N__21359));
    Span4Mux_v I__4960 (
            .O(N__21387),
            .I(N__21359));
    Span4Mux_h I__4959 (
            .O(N__21382),
            .I(N__21359));
    Odrv12 I__4958 (
            .O(N__21377),
            .I(\transmit_module.n3797 ));
    Odrv4 I__4957 (
            .O(N__21368),
            .I(\transmit_module.n3797 ));
    Odrv4 I__4956 (
            .O(N__21359),
            .I(\transmit_module.n3797 ));
    IoInMux I__4955 (
            .O(N__21352),
            .I(N__21344));
    SRMux I__4954 (
            .O(N__21351),
            .I(N__21341));
    SRMux I__4953 (
            .O(N__21350),
            .I(N__21338));
    SRMux I__4952 (
            .O(N__21349),
            .I(N__21335));
    SRMux I__4951 (
            .O(N__21348),
            .I(N__21332));
    SRMux I__4950 (
            .O(N__21347),
            .I(N__21326));
    LocalMux I__4949 (
            .O(N__21344),
            .I(N__21321));
    LocalMux I__4948 (
            .O(N__21341),
            .I(N__21315));
    LocalMux I__4947 (
            .O(N__21338),
            .I(N__21308));
    LocalMux I__4946 (
            .O(N__21335),
            .I(N__21308));
    LocalMux I__4945 (
            .O(N__21332),
            .I(N__21308));
    SRMux I__4944 (
            .O(N__21331),
            .I(N__21305));
    SRMux I__4943 (
            .O(N__21330),
            .I(N__21297));
    SRMux I__4942 (
            .O(N__21329),
            .I(N__21294));
    LocalMux I__4941 (
            .O(N__21326),
            .I(N__21291));
    SRMux I__4940 (
            .O(N__21325),
            .I(N__21288));
    SRMux I__4939 (
            .O(N__21324),
            .I(N__21285));
    IoSpan4Mux I__4938 (
            .O(N__21321),
            .I(N__21277));
    SRMux I__4937 (
            .O(N__21320),
            .I(N__21272));
    SRMux I__4936 (
            .O(N__21319),
            .I(N__21269));
    CascadeMux I__4935 (
            .O(N__21318),
            .I(N__21262));
    Span4Mux_h I__4934 (
            .O(N__21315),
            .I(N__21251));
    Span4Mux_v I__4933 (
            .O(N__21308),
            .I(N__21251));
    LocalMux I__4932 (
            .O(N__21305),
            .I(N__21251));
    SRMux I__4931 (
            .O(N__21304),
            .I(N__21248));
    SRMux I__4930 (
            .O(N__21303),
            .I(N__21245));
    SRMux I__4929 (
            .O(N__21302),
            .I(N__21242));
    SRMux I__4928 (
            .O(N__21301),
            .I(N__21239));
    SRMux I__4927 (
            .O(N__21300),
            .I(N__21236));
    LocalMux I__4926 (
            .O(N__21297),
            .I(N__21230));
    LocalMux I__4925 (
            .O(N__21294),
            .I(N__21221));
    Span4Mux_v I__4924 (
            .O(N__21291),
            .I(N__21221));
    LocalMux I__4923 (
            .O(N__21288),
            .I(N__21221));
    LocalMux I__4922 (
            .O(N__21285),
            .I(N__21221));
    SRMux I__4921 (
            .O(N__21284),
            .I(N__21218));
    SRMux I__4920 (
            .O(N__21283),
            .I(N__21215));
    CascadeMux I__4919 (
            .O(N__21282),
            .I(N__21212));
    CascadeMux I__4918 (
            .O(N__21281),
            .I(N__21209));
    CascadeMux I__4917 (
            .O(N__21280),
            .I(N__21206));
    Span4Mux_s3_h I__4916 (
            .O(N__21277),
            .I(N__21202));
    SRMux I__4915 (
            .O(N__21276),
            .I(N__21199));
    SRMux I__4914 (
            .O(N__21275),
            .I(N__21196));
    LocalMux I__4913 (
            .O(N__21272),
            .I(N__21192));
    LocalMux I__4912 (
            .O(N__21269),
            .I(N__21189));
    CascadeMux I__4911 (
            .O(N__21268),
            .I(N__21186));
    SRMux I__4910 (
            .O(N__21267),
            .I(N__21182));
    SRMux I__4909 (
            .O(N__21266),
            .I(N__21179));
    CascadeMux I__4908 (
            .O(N__21265),
            .I(N__21175));
    InMux I__4907 (
            .O(N__21262),
            .I(N__21172));
    SRMux I__4906 (
            .O(N__21261),
            .I(N__21168));
    SRMux I__4905 (
            .O(N__21260),
            .I(N__21163));
    CascadeMux I__4904 (
            .O(N__21259),
            .I(N__21160));
    CascadeMux I__4903 (
            .O(N__21258),
            .I(N__21157));
    Span4Mux_h I__4902 (
            .O(N__21251),
            .I(N__21152));
    LocalMux I__4901 (
            .O(N__21248),
            .I(N__21152));
    LocalMux I__4900 (
            .O(N__21245),
            .I(N__21145));
    LocalMux I__4899 (
            .O(N__21242),
            .I(N__21145));
    LocalMux I__4898 (
            .O(N__21239),
            .I(N__21145));
    LocalMux I__4897 (
            .O(N__21236),
            .I(N__21142));
    SRMux I__4896 (
            .O(N__21235),
            .I(N__21139));
    CascadeMux I__4895 (
            .O(N__21234),
            .I(N__21135));
    CascadeMux I__4894 (
            .O(N__21233),
            .I(N__21132));
    Span4Mux_v I__4893 (
            .O(N__21230),
            .I(N__21124));
    Span4Mux_v I__4892 (
            .O(N__21221),
            .I(N__21124));
    LocalMux I__4891 (
            .O(N__21218),
            .I(N__21124));
    LocalMux I__4890 (
            .O(N__21215),
            .I(N__21121));
    InMux I__4889 (
            .O(N__21212),
            .I(N__21114));
    InMux I__4888 (
            .O(N__21209),
            .I(N__21111));
    InMux I__4887 (
            .O(N__21206),
            .I(N__21108));
    CascadeMux I__4886 (
            .O(N__21205),
            .I(N__21105));
    Span4Mux_h I__4885 (
            .O(N__21202),
            .I(N__21102));
    LocalMux I__4884 (
            .O(N__21199),
            .I(N__21097));
    LocalMux I__4883 (
            .O(N__21196),
            .I(N__21097));
    SRMux I__4882 (
            .O(N__21195),
            .I(N__21094));
    Span4Mux_h I__4881 (
            .O(N__21192),
            .I(N__21089));
    Span4Mux_v I__4880 (
            .O(N__21189),
            .I(N__21089));
    InMux I__4879 (
            .O(N__21186),
            .I(N__21086));
    SRMux I__4878 (
            .O(N__21185),
            .I(N__21083));
    LocalMux I__4877 (
            .O(N__21182),
            .I(N__21080));
    LocalMux I__4876 (
            .O(N__21179),
            .I(N__21077));
    InMux I__4875 (
            .O(N__21178),
            .I(N__21072));
    InMux I__4874 (
            .O(N__21175),
            .I(N__21072));
    LocalMux I__4873 (
            .O(N__21172),
            .I(N__21069));
    SRMux I__4872 (
            .O(N__21171),
            .I(N__21066));
    LocalMux I__4871 (
            .O(N__21168),
            .I(N__21063));
    CascadeMux I__4870 (
            .O(N__21167),
            .I(N__21060));
    CascadeMux I__4869 (
            .O(N__21166),
            .I(N__21056));
    LocalMux I__4868 (
            .O(N__21163),
            .I(N__21045));
    InMux I__4867 (
            .O(N__21160),
            .I(N__21040));
    InMux I__4866 (
            .O(N__21157),
            .I(N__21040));
    Span4Mux_v I__4865 (
            .O(N__21152),
            .I(N__21037));
    Span4Mux_v I__4864 (
            .O(N__21145),
            .I(N__21030));
    Span4Mux_h I__4863 (
            .O(N__21142),
            .I(N__21030));
    LocalMux I__4862 (
            .O(N__21139),
            .I(N__21030));
    CascadeMux I__4861 (
            .O(N__21138),
            .I(N__21027));
    InMux I__4860 (
            .O(N__21135),
            .I(N__21020));
    InMux I__4859 (
            .O(N__21132),
            .I(N__21020));
    InMux I__4858 (
            .O(N__21131),
            .I(N__21020));
    Span4Mux_h I__4857 (
            .O(N__21124),
            .I(N__21017));
    Span4Mux_h I__4856 (
            .O(N__21121),
            .I(N__21014));
    InMux I__4855 (
            .O(N__21120),
            .I(N__21009));
    InMux I__4854 (
            .O(N__21119),
            .I(N__21009));
    InMux I__4853 (
            .O(N__21118),
            .I(N__21006));
    SRMux I__4852 (
            .O(N__21117),
            .I(N__20999));
    LocalMux I__4851 (
            .O(N__21114),
            .I(N__20992));
    LocalMux I__4850 (
            .O(N__21111),
            .I(N__20992));
    LocalMux I__4849 (
            .O(N__21108),
            .I(N__20992));
    InMux I__4848 (
            .O(N__21105),
            .I(N__20989));
    Span4Mux_h I__4847 (
            .O(N__21102),
            .I(N__20982));
    Span4Mux_v I__4846 (
            .O(N__21097),
            .I(N__20982));
    LocalMux I__4845 (
            .O(N__21094),
            .I(N__20982));
    Span4Mux_h I__4844 (
            .O(N__21089),
            .I(N__20977));
    LocalMux I__4843 (
            .O(N__21086),
            .I(N__20977));
    LocalMux I__4842 (
            .O(N__21083),
            .I(N__20974));
    Span4Mux_v I__4841 (
            .O(N__21080),
            .I(N__20969));
    Span4Mux_v I__4840 (
            .O(N__21077),
            .I(N__20969));
    LocalMux I__4839 (
            .O(N__21072),
            .I(N__20966));
    Span4Mux_v I__4838 (
            .O(N__21069),
            .I(N__20963));
    LocalMux I__4837 (
            .O(N__21066),
            .I(N__20960));
    Span4Mux_v I__4836 (
            .O(N__21063),
            .I(N__20957));
    InMux I__4835 (
            .O(N__21060),
            .I(N__20952));
    InMux I__4834 (
            .O(N__21059),
            .I(N__20952));
    InMux I__4833 (
            .O(N__21056),
            .I(N__20945));
    InMux I__4832 (
            .O(N__21055),
            .I(N__20945));
    InMux I__4831 (
            .O(N__21054),
            .I(N__20945));
    SRMux I__4830 (
            .O(N__21053),
            .I(N__20942));
    InMux I__4829 (
            .O(N__21052),
            .I(N__20937));
    InMux I__4828 (
            .O(N__21051),
            .I(N__20937));
    SRMux I__4827 (
            .O(N__21050),
            .I(N__20934));
    SRMux I__4826 (
            .O(N__21049),
            .I(N__20931));
    SRMux I__4825 (
            .O(N__21048),
            .I(N__20928));
    Span4Mux_v I__4824 (
            .O(N__21045),
            .I(N__20925));
    LocalMux I__4823 (
            .O(N__21040),
            .I(N__20918));
    Span4Mux_h I__4822 (
            .O(N__21037),
            .I(N__20918));
    Span4Mux_h I__4821 (
            .O(N__21030),
            .I(N__20918));
    InMux I__4820 (
            .O(N__21027),
            .I(N__20915));
    LocalMux I__4819 (
            .O(N__21020),
            .I(N__20908));
    Span4Mux_h I__4818 (
            .O(N__21017),
            .I(N__20908));
    Span4Mux_v I__4817 (
            .O(N__21014),
            .I(N__20908));
    LocalMux I__4816 (
            .O(N__21009),
            .I(N__20903));
    LocalMux I__4815 (
            .O(N__21006),
            .I(N__20903));
    InMux I__4814 (
            .O(N__21005),
            .I(N__20898));
    InMux I__4813 (
            .O(N__21004),
            .I(N__20898));
    InMux I__4812 (
            .O(N__21003),
            .I(N__20893));
    InMux I__4811 (
            .O(N__21002),
            .I(N__20893));
    LocalMux I__4810 (
            .O(N__20999),
            .I(N__20886));
    Span12Mux_v I__4809 (
            .O(N__20992),
            .I(N__20886));
    LocalMux I__4808 (
            .O(N__20989),
            .I(N__20886));
    Span4Mux_v I__4807 (
            .O(N__20982),
            .I(N__20873));
    Span4Mux_v I__4806 (
            .O(N__20977),
            .I(N__20873));
    Span4Mux_h I__4805 (
            .O(N__20974),
            .I(N__20873));
    Span4Mux_h I__4804 (
            .O(N__20969),
            .I(N__20873));
    Span4Mux_v I__4803 (
            .O(N__20966),
            .I(N__20873));
    Span4Mux_v I__4802 (
            .O(N__20963),
            .I(N__20873));
    Sp12to4 I__4801 (
            .O(N__20960),
            .I(N__20864));
    Sp12to4 I__4800 (
            .O(N__20957),
            .I(N__20864));
    LocalMux I__4799 (
            .O(N__20952),
            .I(N__20864));
    LocalMux I__4798 (
            .O(N__20945),
            .I(N__20864));
    LocalMux I__4797 (
            .O(N__20942),
            .I(ADV_VSYNC_c));
    LocalMux I__4796 (
            .O(N__20937),
            .I(ADV_VSYNC_c));
    LocalMux I__4795 (
            .O(N__20934),
            .I(ADV_VSYNC_c));
    LocalMux I__4794 (
            .O(N__20931),
            .I(ADV_VSYNC_c));
    LocalMux I__4793 (
            .O(N__20928),
            .I(ADV_VSYNC_c));
    Odrv4 I__4792 (
            .O(N__20925),
            .I(ADV_VSYNC_c));
    Odrv4 I__4791 (
            .O(N__20918),
            .I(ADV_VSYNC_c));
    LocalMux I__4790 (
            .O(N__20915),
            .I(ADV_VSYNC_c));
    Odrv4 I__4789 (
            .O(N__20908),
            .I(ADV_VSYNC_c));
    Odrv12 I__4788 (
            .O(N__20903),
            .I(ADV_VSYNC_c));
    LocalMux I__4787 (
            .O(N__20898),
            .I(ADV_VSYNC_c));
    LocalMux I__4786 (
            .O(N__20893),
            .I(ADV_VSYNC_c));
    Odrv12 I__4785 (
            .O(N__20886),
            .I(ADV_VSYNC_c));
    Odrv4 I__4784 (
            .O(N__20873),
            .I(ADV_VSYNC_c));
    Odrv12 I__4783 (
            .O(N__20864),
            .I(ADV_VSYNC_c));
    InMux I__4782 (
            .O(N__20833),
            .I(N__20830));
    LocalMux I__4781 (
            .O(N__20830),
            .I(N__20827));
    Sp12to4 I__4780 (
            .O(N__20827),
            .I(N__20824));
    Span12Mux_v I__4779 (
            .O(N__20824),
            .I(N__20821));
    Odrv12 I__4778 (
            .O(N__20821),
            .I(\line_buffer.n544 ));
    InMux I__4777 (
            .O(N__20818),
            .I(N__20815));
    LocalMux I__4776 (
            .O(N__20815),
            .I(N__20812));
    Span4Mux_h I__4775 (
            .O(N__20812),
            .I(N__20809));
    Span4Mux_h I__4774 (
            .O(N__20809),
            .I(N__20806));
    Odrv4 I__4773 (
            .O(N__20806),
            .I(\line_buffer.n536 ));
    InMux I__4772 (
            .O(N__20803),
            .I(N__20800));
    LocalMux I__4771 (
            .O(N__20800),
            .I(N__20797));
    Span4Mux_v I__4770 (
            .O(N__20797),
            .I(N__20794));
    Odrv4 I__4769 (
            .O(N__20794),
            .I(\line_buffer.n3698 ));
    InMux I__4768 (
            .O(N__20791),
            .I(N__20788));
    LocalMux I__4767 (
            .O(N__20788),
            .I(N__20785));
    Sp12to4 I__4766 (
            .O(N__20785),
            .I(N__20782));
    Span12Mux_v I__4765 (
            .O(N__20782),
            .I(N__20779));
    Odrv12 I__4764 (
            .O(N__20779),
            .I(\line_buffer.n508 ));
    CascadeMux I__4763 (
            .O(N__20776),
            .I(N__20773));
    InMux I__4762 (
            .O(N__20773),
            .I(N__20770));
    LocalMux I__4761 (
            .O(N__20770),
            .I(N__20767));
    Span4Mux_h I__4760 (
            .O(N__20767),
            .I(N__20764));
    Span4Mux_h I__4759 (
            .O(N__20764),
            .I(N__20761));
    Span4Mux_v I__4758 (
            .O(N__20761),
            .I(N__20758));
    Odrv4 I__4757 (
            .O(N__20758),
            .I(\line_buffer.n500 ));
    CascadeMux I__4756 (
            .O(N__20755),
            .I(\line_buffer.n3695_cascade_ ));
    InMux I__4755 (
            .O(N__20752),
            .I(N__20749));
    LocalMux I__4754 (
            .O(N__20749),
            .I(N__20746));
    Span4Mux_v I__4753 (
            .O(N__20746),
            .I(N__20743));
    Odrv4 I__4752 (
            .O(N__20743),
            .I(TX_DATA_1));
    InMux I__4751 (
            .O(N__20740),
            .I(N__20737));
    LocalMux I__4750 (
            .O(N__20737),
            .I(N__20734));
    Span4Mux_v I__4749 (
            .O(N__20734),
            .I(N__20731));
    Sp12to4 I__4748 (
            .O(N__20731),
            .I(N__20728));
    Odrv12 I__4747 (
            .O(N__20728),
            .I(\line_buffer.n572 ));
    InMux I__4746 (
            .O(N__20725),
            .I(N__20722));
    LocalMux I__4745 (
            .O(N__20722),
            .I(N__20719));
    Span4Mux_v I__4744 (
            .O(N__20719),
            .I(N__20716));
    Sp12to4 I__4743 (
            .O(N__20716),
            .I(N__20713));
    Span12Mux_h I__4742 (
            .O(N__20713),
            .I(N__20710));
    Span12Mux_v I__4741 (
            .O(N__20710),
            .I(N__20707));
    Odrv12 I__4740 (
            .O(N__20707),
            .I(\line_buffer.n564 ));
    InMux I__4739 (
            .O(N__20704),
            .I(N__20701));
    LocalMux I__4738 (
            .O(N__20701),
            .I(\line_buffer.n3692 ));
    InMux I__4737 (
            .O(N__20698),
            .I(N__20680));
    InMux I__4736 (
            .O(N__20697),
            .I(N__20680));
    InMux I__4735 (
            .O(N__20696),
            .I(N__20680));
    InMux I__4734 (
            .O(N__20695),
            .I(N__20680));
    InMux I__4733 (
            .O(N__20694),
            .I(N__20680));
    InMux I__4732 (
            .O(N__20693),
            .I(N__20680));
    LocalMux I__4731 (
            .O(N__20680),
            .I(N__20675));
    InMux I__4730 (
            .O(N__20679),
            .I(N__20669));
    InMux I__4729 (
            .O(N__20678),
            .I(N__20666));
    Span4Mux_v I__4728 (
            .O(N__20675),
            .I(N__20663));
    InMux I__4727 (
            .O(N__20674),
            .I(N__20658));
    InMux I__4726 (
            .O(N__20673),
            .I(N__20658));
    InMux I__4725 (
            .O(N__20672),
            .I(N__20655));
    LocalMux I__4724 (
            .O(N__20669),
            .I(N__20652));
    LocalMux I__4723 (
            .O(N__20666),
            .I(N__20647));
    Span4Mux_v I__4722 (
            .O(N__20663),
            .I(N__20647));
    LocalMux I__4721 (
            .O(N__20658),
            .I(N__20644));
    LocalMux I__4720 (
            .O(N__20655),
            .I(N__20637));
    Span4Mux_h I__4719 (
            .O(N__20652),
            .I(N__20637));
    Span4Mux_v I__4718 (
            .O(N__20647),
            .I(N__20637));
    Span4Mux_v I__4717 (
            .O(N__20644),
            .I(N__20625));
    Span4Mux_v I__4716 (
            .O(N__20637),
            .I(N__20622));
    InMux I__4715 (
            .O(N__20636),
            .I(N__20617));
    InMux I__4714 (
            .O(N__20635),
            .I(N__20617));
    InMux I__4713 (
            .O(N__20634),
            .I(N__20614));
    InMux I__4712 (
            .O(N__20633),
            .I(N__20611));
    InMux I__4711 (
            .O(N__20632),
            .I(N__20608));
    InMux I__4710 (
            .O(N__20631),
            .I(N__20599));
    InMux I__4709 (
            .O(N__20630),
            .I(N__20599));
    InMux I__4708 (
            .O(N__20629),
            .I(N__20599));
    InMux I__4707 (
            .O(N__20628),
            .I(N__20599));
    Odrv4 I__4706 (
            .O(N__20625),
            .I(RX_WE));
    Odrv4 I__4705 (
            .O(N__20622),
            .I(RX_WE));
    LocalMux I__4704 (
            .O(N__20617),
            .I(RX_WE));
    LocalMux I__4703 (
            .O(N__20614),
            .I(RX_WE));
    LocalMux I__4702 (
            .O(N__20611),
            .I(RX_WE));
    LocalMux I__4701 (
            .O(N__20608),
            .I(RX_WE));
    LocalMux I__4700 (
            .O(N__20599),
            .I(RX_WE));
    InMux I__4699 (
            .O(N__20584),
            .I(N__20581));
    LocalMux I__4698 (
            .O(N__20581),
            .I(N__20578));
    Span4Mux_v I__4697 (
            .O(N__20578),
            .I(N__20575));
    Span4Mux_v I__4696 (
            .O(N__20575),
            .I(N__20572));
    Odrv4 I__4695 (
            .O(N__20572),
            .I(\receive_module.n133 ));
    CascadeMux I__4694 (
            .O(N__20569),
            .I(N__20561));
    CascadeMux I__4693 (
            .O(N__20568),
            .I(N__20558));
    CascadeMux I__4692 (
            .O(N__20567),
            .I(N__20554));
    CascadeMux I__4691 (
            .O(N__20566),
            .I(N__20551));
    InMux I__4690 (
            .O(N__20565),
            .I(N__20546));
    InMux I__4689 (
            .O(N__20564),
            .I(N__20546));
    InMux I__4688 (
            .O(N__20561),
            .I(N__20537));
    InMux I__4687 (
            .O(N__20558),
            .I(N__20537));
    InMux I__4686 (
            .O(N__20557),
            .I(N__20537));
    InMux I__4685 (
            .O(N__20554),
            .I(N__20537));
    InMux I__4684 (
            .O(N__20551),
            .I(N__20531));
    LocalMux I__4683 (
            .O(N__20546),
            .I(N__20528));
    LocalMux I__4682 (
            .O(N__20537),
            .I(N__20525));
    CascadeMux I__4681 (
            .O(N__20536),
            .I(N__20522));
    CascadeMux I__4680 (
            .O(N__20535),
            .I(N__20518));
    InMux I__4679 (
            .O(N__20534),
            .I(N__20515));
    LocalMux I__4678 (
            .O(N__20531),
            .I(N__20512));
    Span4Mux_v I__4677 (
            .O(N__20528),
            .I(N__20507));
    Span4Mux_v I__4676 (
            .O(N__20525),
            .I(N__20507));
    InMux I__4675 (
            .O(N__20522),
            .I(N__20504));
    InMux I__4674 (
            .O(N__20521),
            .I(N__20498));
    InMux I__4673 (
            .O(N__20518),
            .I(N__20498));
    LocalMux I__4672 (
            .O(N__20515),
            .I(N__20495));
    Span4Mux_v I__4671 (
            .O(N__20512),
            .I(N__20492));
    Span4Mux_v I__4670 (
            .O(N__20507),
            .I(N__20487));
    LocalMux I__4669 (
            .O(N__20504),
            .I(N__20487));
    CascadeMux I__4668 (
            .O(N__20503),
            .I(N__20484));
    LocalMux I__4667 (
            .O(N__20498),
            .I(N__20480));
    Span4Mux_v I__4666 (
            .O(N__20495),
            .I(N__20477));
    Span4Mux_h I__4665 (
            .O(N__20492),
            .I(N__20472));
    Span4Mux_v I__4664 (
            .O(N__20487),
            .I(N__20472));
    InMux I__4663 (
            .O(N__20484),
            .I(N__20469));
    InMux I__4662 (
            .O(N__20483),
            .I(N__20466));
    Span4Mux_h I__4661 (
            .O(N__20480),
            .I(N__20459));
    Sp12to4 I__4660 (
            .O(N__20477),
            .I(N__20456));
    Sp12to4 I__4659 (
            .O(N__20472),
            .I(N__20449));
    LocalMux I__4658 (
            .O(N__20469),
            .I(N__20449));
    LocalMux I__4657 (
            .O(N__20466),
            .I(N__20449));
    InMux I__4656 (
            .O(N__20465),
            .I(N__20446));
    InMux I__4655 (
            .O(N__20464),
            .I(N__20439));
    InMux I__4654 (
            .O(N__20463),
            .I(N__20439));
    InMux I__4653 (
            .O(N__20462),
            .I(N__20439));
    Span4Mux_v I__4652 (
            .O(N__20459),
            .I(N__20436));
    Span12Mux_h I__4651 (
            .O(N__20456),
            .I(N__20427));
    Span12Mux_v I__4650 (
            .O(N__20449),
            .I(N__20427));
    LocalMux I__4649 (
            .O(N__20446),
            .I(N__20427));
    LocalMux I__4648 (
            .O(N__20439),
            .I(N__20427));
    Odrv4 I__4647 (
            .O(N__20436),
            .I(TVP_VSYNC_c));
    Odrv12 I__4646 (
            .O(N__20427),
            .I(TVP_VSYNC_c));
    CascadeMux I__4645 (
            .O(N__20422),
            .I(N__20418));
    CascadeMux I__4644 (
            .O(N__20421),
            .I(N__20415));
    CascadeBuf I__4643 (
            .O(N__20418),
            .I(N__20412));
    CascadeBuf I__4642 (
            .O(N__20415),
            .I(N__20409));
    CascadeMux I__4641 (
            .O(N__20412),
            .I(N__20406));
    CascadeMux I__4640 (
            .O(N__20409),
            .I(N__20403));
    CascadeBuf I__4639 (
            .O(N__20406),
            .I(N__20400));
    CascadeBuf I__4638 (
            .O(N__20403),
            .I(N__20397));
    CascadeMux I__4637 (
            .O(N__20400),
            .I(N__20394));
    CascadeMux I__4636 (
            .O(N__20397),
            .I(N__20391));
    CascadeBuf I__4635 (
            .O(N__20394),
            .I(N__20388));
    CascadeBuf I__4634 (
            .O(N__20391),
            .I(N__20385));
    CascadeMux I__4633 (
            .O(N__20388),
            .I(N__20382));
    CascadeMux I__4632 (
            .O(N__20385),
            .I(N__20379));
    CascadeBuf I__4631 (
            .O(N__20382),
            .I(N__20376));
    CascadeBuf I__4630 (
            .O(N__20379),
            .I(N__20373));
    CascadeMux I__4629 (
            .O(N__20376),
            .I(N__20370));
    CascadeMux I__4628 (
            .O(N__20373),
            .I(N__20367));
    CascadeBuf I__4627 (
            .O(N__20370),
            .I(N__20364));
    CascadeBuf I__4626 (
            .O(N__20367),
            .I(N__20361));
    CascadeMux I__4625 (
            .O(N__20364),
            .I(N__20358));
    CascadeMux I__4624 (
            .O(N__20361),
            .I(N__20355));
    CascadeBuf I__4623 (
            .O(N__20358),
            .I(N__20352));
    CascadeBuf I__4622 (
            .O(N__20355),
            .I(N__20349));
    CascadeMux I__4621 (
            .O(N__20352),
            .I(N__20346));
    CascadeMux I__4620 (
            .O(N__20349),
            .I(N__20343));
    CascadeBuf I__4619 (
            .O(N__20346),
            .I(N__20340));
    CascadeBuf I__4618 (
            .O(N__20343),
            .I(N__20337));
    CascadeMux I__4617 (
            .O(N__20340),
            .I(N__20334));
    CascadeMux I__4616 (
            .O(N__20337),
            .I(N__20331));
    CascadeBuf I__4615 (
            .O(N__20334),
            .I(N__20328));
    CascadeBuf I__4614 (
            .O(N__20331),
            .I(N__20325));
    CascadeMux I__4613 (
            .O(N__20328),
            .I(N__20322));
    CascadeMux I__4612 (
            .O(N__20325),
            .I(N__20319));
    CascadeBuf I__4611 (
            .O(N__20322),
            .I(N__20316));
    CascadeBuf I__4610 (
            .O(N__20319),
            .I(N__20313));
    CascadeMux I__4609 (
            .O(N__20316),
            .I(N__20310));
    CascadeMux I__4608 (
            .O(N__20313),
            .I(N__20307));
    CascadeBuf I__4607 (
            .O(N__20310),
            .I(N__20304));
    CascadeBuf I__4606 (
            .O(N__20307),
            .I(N__20301));
    CascadeMux I__4605 (
            .O(N__20304),
            .I(N__20298));
    CascadeMux I__4604 (
            .O(N__20301),
            .I(N__20295));
    CascadeBuf I__4603 (
            .O(N__20298),
            .I(N__20292));
    CascadeBuf I__4602 (
            .O(N__20295),
            .I(N__20289));
    CascadeMux I__4601 (
            .O(N__20292),
            .I(N__20286));
    CascadeMux I__4600 (
            .O(N__20289),
            .I(N__20283));
    CascadeBuf I__4599 (
            .O(N__20286),
            .I(N__20280));
    CascadeBuf I__4598 (
            .O(N__20283),
            .I(N__20277));
    CascadeMux I__4597 (
            .O(N__20280),
            .I(N__20274));
    CascadeMux I__4596 (
            .O(N__20277),
            .I(N__20271));
    CascadeBuf I__4595 (
            .O(N__20274),
            .I(N__20268));
    CascadeBuf I__4594 (
            .O(N__20271),
            .I(N__20265));
    CascadeMux I__4593 (
            .O(N__20268),
            .I(N__20262));
    CascadeMux I__4592 (
            .O(N__20265),
            .I(N__20259));
    CascadeBuf I__4591 (
            .O(N__20262),
            .I(N__20256));
    CascadeBuf I__4590 (
            .O(N__20259),
            .I(N__20253));
    CascadeMux I__4589 (
            .O(N__20256),
            .I(N__20250));
    CascadeMux I__4588 (
            .O(N__20253),
            .I(N__20247));
    CascadeBuf I__4587 (
            .O(N__20250),
            .I(N__20244));
    CascadeBuf I__4586 (
            .O(N__20247),
            .I(N__20241));
    CascadeMux I__4585 (
            .O(N__20244),
            .I(N__20237));
    CascadeMux I__4584 (
            .O(N__20241),
            .I(N__20234));
    CascadeMux I__4583 (
            .O(N__20240),
            .I(N__20231));
    InMux I__4582 (
            .O(N__20237),
            .I(N__20228));
    InMux I__4581 (
            .O(N__20234),
            .I(N__20225));
    InMux I__4580 (
            .O(N__20231),
            .I(N__20222));
    LocalMux I__4579 (
            .O(N__20228),
            .I(N__20219));
    LocalMux I__4578 (
            .O(N__20225),
            .I(N__20216));
    LocalMux I__4577 (
            .O(N__20222),
            .I(N__20213));
    Span4Mux_h I__4576 (
            .O(N__20219),
            .I(N__20210));
    Span12Mux_s1_v I__4575 (
            .O(N__20216),
            .I(N__20206));
    Sp12to4 I__4574 (
            .O(N__20213),
            .I(N__20203));
    Sp12to4 I__4573 (
            .O(N__20210),
            .I(N__20200));
    InMux I__4572 (
            .O(N__20209),
            .I(N__20197));
    Span12Mux_v I__4571 (
            .O(N__20206),
            .I(N__20194));
    Span12Mux_v I__4570 (
            .O(N__20203),
            .I(N__20189));
    Span12Mux_v I__4569 (
            .O(N__20200),
            .I(N__20189));
    LocalMux I__4568 (
            .O(N__20197),
            .I(RX_ADDR_3));
    Odrv12 I__4567 (
            .O(N__20194),
            .I(RX_ADDR_3));
    Odrv12 I__4566 (
            .O(N__20189),
            .I(RX_ADDR_3));
    InMux I__4565 (
            .O(N__20182),
            .I(N__20179));
    LocalMux I__4564 (
            .O(N__20179),
            .I(N__20167));
    ClkMux I__4563 (
            .O(N__20178),
            .I(N__20029));
    ClkMux I__4562 (
            .O(N__20177),
            .I(N__20029));
    ClkMux I__4561 (
            .O(N__20176),
            .I(N__20029));
    ClkMux I__4560 (
            .O(N__20175),
            .I(N__20029));
    ClkMux I__4559 (
            .O(N__20174),
            .I(N__20029));
    ClkMux I__4558 (
            .O(N__20173),
            .I(N__20029));
    ClkMux I__4557 (
            .O(N__20172),
            .I(N__20029));
    ClkMux I__4556 (
            .O(N__20171),
            .I(N__20029));
    ClkMux I__4555 (
            .O(N__20170),
            .I(N__20029));
    Glb2LocalMux I__4554 (
            .O(N__20167),
            .I(N__20029));
    ClkMux I__4553 (
            .O(N__20166),
            .I(N__20029));
    ClkMux I__4552 (
            .O(N__20165),
            .I(N__20029));
    ClkMux I__4551 (
            .O(N__20164),
            .I(N__20029));
    ClkMux I__4550 (
            .O(N__20163),
            .I(N__20029));
    ClkMux I__4549 (
            .O(N__20162),
            .I(N__20029));
    ClkMux I__4548 (
            .O(N__20161),
            .I(N__20029));
    ClkMux I__4547 (
            .O(N__20160),
            .I(N__20029));
    ClkMux I__4546 (
            .O(N__20159),
            .I(N__20029));
    ClkMux I__4545 (
            .O(N__20158),
            .I(N__20029));
    ClkMux I__4544 (
            .O(N__20157),
            .I(N__20029));
    ClkMux I__4543 (
            .O(N__20156),
            .I(N__20029));
    ClkMux I__4542 (
            .O(N__20155),
            .I(N__20029));
    ClkMux I__4541 (
            .O(N__20154),
            .I(N__20029));
    ClkMux I__4540 (
            .O(N__20153),
            .I(N__20029));
    ClkMux I__4539 (
            .O(N__20152),
            .I(N__20029));
    ClkMux I__4538 (
            .O(N__20151),
            .I(N__20029));
    ClkMux I__4537 (
            .O(N__20150),
            .I(N__20029));
    ClkMux I__4536 (
            .O(N__20149),
            .I(N__20029));
    ClkMux I__4535 (
            .O(N__20148),
            .I(N__20029));
    ClkMux I__4534 (
            .O(N__20147),
            .I(N__20029));
    ClkMux I__4533 (
            .O(N__20146),
            .I(N__20029));
    ClkMux I__4532 (
            .O(N__20145),
            .I(N__20029));
    ClkMux I__4531 (
            .O(N__20144),
            .I(N__20029));
    ClkMux I__4530 (
            .O(N__20143),
            .I(N__20029));
    ClkMux I__4529 (
            .O(N__20142),
            .I(N__20029));
    ClkMux I__4528 (
            .O(N__20141),
            .I(N__20029));
    ClkMux I__4527 (
            .O(N__20140),
            .I(N__20029));
    ClkMux I__4526 (
            .O(N__20139),
            .I(N__20029));
    ClkMux I__4525 (
            .O(N__20138),
            .I(N__20029));
    ClkMux I__4524 (
            .O(N__20137),
            .I(N__20029));
    ClkMux I__4523 (
            .O(N__20136),
            .I(N__20029));
    ClkMux I__4522 (
            .O(N__20135),
            .I(N__20029));
    ClkMux I__4521 (
            .O(N__20134),
            .I(N__20029));
    ClkMux I__4520 (
            .O(N__20133),
            .I(N__20029));
    ClkMux I__4519 (
            .O(N__20132),
            .I(N__20029));
    ClkMux I__4518 (
            .O(N__20131),
            .I(N__20029));
    ClkMux I__4517 (
            .O(N__20130),
            .I(N__20029));
    ClkMux I__4516 (
            .O(N__20129),
            .I(N__20029));
    ClkMux I__4515 (
            .O(N__20128),
            .I(N__20029));
    GlobalMux I__4514 (
            .O(N__20029),
            .I(N__20026));
    gio2CtrlBuf I__4513 (
            .O(N__20026),
            .I(TVP_CLK_c));
    InMux I__4512 (
            .O(N__20023),
            .I(N__20020));
    LocalMux I__4511 (
            .O(N__20020),
            .I(\transmit_module.Y_DELTA_PATTERN_32 ));
    InMux I__4510 (
            .O(N__20017),
            .I(N__20014));
    LocalMux I__4509 (
            .O(N__20014),
            .I(\transmit_module.Y_DELTA_PATTERN_31 ));
    InMux I__4508 (
            .O(N__20011),
            .I(N__20008));
    LocalMux I__4507 (
            .O(N__20008),
            .I(\transmit_module.Y_DELTA_PATTERN_22 ));
    InMux I__4506 (
            .O(N__20005),
            .I(N__20002));
    LocalMux I__4505 (
            .O(N__20002),
            .I(\transmit_module.Y_DELTA_PATTERN_24 ));
    InMux I__4504 (
            .O(N__19999),
            .I(N__19996));
    LocalMux I__4503 (
            .O(N__19996),
            .I(\transmit_module.Y_DELTA_PATTERN_23 ));
    InMux I__4502 (
            .O(N__19993),
            .I(N__19990));
    LocalMux I__4501 (
            .O(N__19990),
            .I(\transmit_module.Y_DELTA_PATTERN_16 ));
    InMux I__4500 (
            .O(N__19987),
            .I(N__19984));
    LocalMux I__4499 (
            .O(N__19984),
            .I(\transmit_module.Y_DELTA_PATTERN_17 ));
    InMux I__4498 (
            .O(N__19981),
            .I(N__19978));
    LocalMux I__4497 (
            .O(N__19978),
            .I(\transmit_module.Y_DELTA_PATTERN_19 ));
    InMux I__4496 (
            .O(N__19975),
            .I(N__19972));
    LocalMux I__4495 (
            .O(N__19972),
            .I(\transmit_module.Y_DELTA_PATTERN_18 ));
    InMux I__4494 (
            .O(N__19969),
            .I(N__19966));
    LocalMux I__4493 (
            .O(N__19966),
            .I(N__19963));
    Odrv12 I__4492 (
            .O(N__19963),
            .I(\line_buffer.n3737 ));
    InMux I__4491 (
            .O(N__19960),
            .I(N__19957));
    LocalMux I__4490 (
            .O(N__19957),
            .I(N__19954));
    Span4Mux_h I__4489 (
            .O(N__19954),
            .I(N__19951));
    Span4Mux_h I__4488 (
            .O(N__19951),
            .I(N__19948));
    Odrv4 I__4487 (
            .O(N__19948),
            .I(\line_buffer.n447 ));
    CascadeMux I__4486 (
            .O(N__19945),
            .I(N__19942));
    InMux I__4485 (
            .O(N__19942),
            .I(N__19939));
    LocalMux I__4484 (
            .O(N__19939),
            .I(N__19936));
    Span4Mux_v I__4483 (
            .O(N__19936),
            .I(N__19933));
    Sp12to4 I__4482 (
            .O(N__19933),
            .I(N__19930));
    Span12Mux_h I__4481 (
            .O(N__19930),
            .I(N__19927));
    Odrv12 I__4480 (
            .O(N__19927),
            .I(\line_buffer.n439 ));
    InMux I__4479 (
            .O(N__19924),
            .I(N__19921));
    LocalMux I__4478 (
            .O(N__19921),
            .I(\line_buffer.n3701 ));
    InMux I__4477 (
            .O(N__19918),
            .I(N__19915));
    LocalMux I__4476 (
            .O(N__19915),
            .I(N__19912));
    Odrv12 I__4475 (
            .O(N__19912),
            .I(TX_DATA_5));
    IoInMux I__4474 (
            .O(N__19909),
            .I(N__19906));
    LocalMux I__4473 (
            .O(N__19906),
            .I(N__19902));
    IoInMux I__4472 (
            .O(N__19905),
            .I(N__19899));
    IoSpan4Mux I__4471 (
            .O(N__19902),
            .I(N__19895));
    LocalMux I__4470 (
            .O(N__19899),
            .I(N__19892));
    IoInMux I__4469 (
            .O(N__19898),
            .I(N__19889));
    Span4Mux_s3_v I__4468 (
            .O(N__19895),
            .I(N__19886));
    Span4Mux_s3_v I__4467 (
            .O(N__19892),
            .I(N__19883));
    LocalMux I__4466 (
            .O(N__19889),
            .I(N__19880));
    Span4Mux_h I__4465 (
            .O(N__19886),
            .I(N__19877));
    Span4Mux_h I__4464 (
            .O(N__19883),
            .I(N__19874));
    Span12Mux_s4_h I__4463 (
            .O(N__19880),
            .I(N__19871));
    Span4Mux_h I__4462 (
            .O(N__19877),
            .I(N__19866));
    Span4Mux_h I__4461 (
            .O(N__19874),
            .I(N__19866));
    Span12Mux_h I__4460 (
            .O(N__19871),
            .I(N__19863));
    Span4Mux_v I__4459 (
            .O(N__19866),
            .I(N__19860));
    Odrv12 I__4458 (
            .O(N__19863),
            .I(n1793));
    Odrv4 I__4457 (
            .O(N__19860),
            .I(n1793));
    SRMux I__4456 (
            .O(N__19855),
            .I(N__19852));
    LocalMux I__4455 (
            .O(N__19852),
            .I(N__19847));
    SRMux I__4454 (
            .O(N__19851),
            .I(N__19844));
    SRMux I__4453 (
            .O(N__19850),
            .I(N__19840));
    Span4Mux_v I__4452 (
            .O(N__19847),
            .I(N__19833));
    LocalMux I__4451 (
            .O(N__19844),
            .I(N__19833));
    SRMux I__4450 (
            .O(N__19843),
            .I(N__19830));
    LocalMux I__4449 (
            .O(N__19840),
            .I(N__19826));
    SRMux I__4448 (
            .O(N__19839),
            .I(N__19823));
    SRMux I__4447 (
            .O(N__19838),
            .I(N__19820));
    Span4Mux_h I__4446 (
            .O(N__19833),
            .I(N__19813));
    LocalMux I__4445 (
            .O(N__19830),
            .I(N__19813));
    SRMux I__4444 (
            .O(N__19829),
            .I(N__19810));
    Span4Mux_s0_v I__4443 (
            .O(N__19826),
            .I(N__19802));
    LocalMux I__4442 (
            .O(N__19823),
            .I(N__19802));
    LocalMux I__4441 (
            .O(N__19820),
            .I(N__19799));
    SRMux I__4440 (
            .O(N__19819),
            .I(N__19796));
    SRMux I__4439 (
            .O(N__19818),
            .I(N__19793));
    Span4Mux_v I__4438 (
            .O(N__19813),
            .I(N__19786));
    LocalMux I__4437 (
            .O(N__19810),
            .I(N__19786));
    SRMux I__4436 (
            .O(N__19809),
            .I(N__19783));
    SRMux I__4435 (
            .O(N__19808),
            .I(N__19780));
    SRMux I__4434 (
            .O(N__19807),
            .I(N__19777));
    Span4Mux_v I__4433 (
            .O(N__19802),
            .I(N__19769));
    Span4Mux_h I__4432 (
            .O(N__19799),
            .I(N__19769));
    LocalMux I__4431 (
            .O(N__19796),
            .I(N__19769));
    LocalMux I__4430 (
            .O(N__19793),
            .I(N__19766));
    SRMux I__4429 (
            .O(N__19792),
            .I(N__19763));
    SRMux I__4428 (
            .O(N__19791),
            .I(N__19760));
    Span4Mux_h I__4427 (
            .O(N__19786),
            .I(N__19752));
    LocalMux I__4426 (
            .O(N__19783),
            .I(N__19752));
    LocalMux I__4425 (
            .O(N__19780),
            .I(N__19747));
    LocalMux I__4424 (
            .O(N__19777),
            .I(N__19747));
    SRMux I__4423 (
            .O(N__19776),
            .I(N__19744));
    Span4Mux_v I__4422 (
            .O(N__19769),
            .I(N__19739));
    Span4Mux_h I__4421 (
            .O(N__19766),
            .I(N__19734));
    LocalMux I__4420 (
            .O(N__19763),
            .I(N__19734));
    LocalMux I__4419 (
            .O(N__19760),
            .I(N__19731));
    SRMux I__4418 (
            .O(N__19759),
            .I(N__19728));
    SRMux I__4417 (
            .O(N__19758),
            .I(N__19725));
    SRMux I__4416 (
            .O(N__19757),
            .I(N__19720));
    Span4Mux_v I__4415 (
            .O(N__19752),
            .I(N__19715));
    Span4Mux_v I__4414 (
            .O(N__19747),
            .I(N__19712));
    LocalMux I__4413 (
            .O(N__19744),
            .I(N__19709));
    SRMux I__4412 (
            .O(N__19743),
            .I(N__19706));
    SRMux I__4411 (
            .O(N__19742),
            .I(N__19701));
    Span4Mux_v I__4410 (
            .O(N__19739),
            .I(N__19690));
    Span4Mux_v I__4409 (
            .O(N__19734),
            .I(N__19690));
    Span4Mux_h I__4408 (
            .O(N__19731),
            .I(N__19690));
    LocalMux I__4407 (
            .O(N__19728),
            .I(N__19690));
    LocalMux I__4406 (
            .O(N__19725),
            .I(N__19687));
    SRMux I__4405 (
            .O(N__19724),
            .I(N__19684));
    SRMux I__4404 (
            .O(N__19723),
            .I(N__19681));
    LocalMux I__4403 (
            .O(N__19720),
            .I(N__19677));
    SRMux I__4402 (
            .O(N__19719),
            .I(N__19674));
    SRMux I__4401 (
            .O(N__19718),
            .I(N__19671));
    Span4Mux_v I__4400 (
            .O(N__19715),
            .I(N__19668));
    Span4Mux_v I__4399 (
            .O(N__19712),
            .I(N__19661));
    Span4Mux_v I__4398 (
            .O(N__19709),
            .I(N__19661));
    LocalMux I__4397 (
            .O(N__19706),
            .I(N__19661));
    SRMux I__4396 (
            .O(N__19705),
            .I(N__19658));
    SRMux I__4395 (
            .O(N__19704),
            .I(N__19653));
    LocalMux I__4394 (
            .O(N__19701),
            .I(N__19649));
    SRMux I__4393 (
            .O(N__19700),
            .I(N__19646));
    SRMux I__4392 (
            .O(N__19699),
            .I(N__19643));
    Span4Mux_v I__4391 (
            .O(N__19690),
            .I(N__19636));
    Span4Mux_h I__4390 (
            .O(N__19687),
            .I(N__19636));
    LocalMux I__4389 (
            .O(N__19684),
            .I(N__19636));
    LocalMux I__4388 (
            .O(N__19681),
            .I(N__19633));
    SRMux I__4387 (
            .O(N__19680),
            .I(N__19630));
    Span4Mux_s3_v I__4386 (
            .O(N__19677),
            .I(N__19622));
    LocalMux I__4385 (
            .O(N__19674),
            .I(N__19622));
    LocalMux I__4384 (
            .O(N__19671),
            .I(N__19622));
    Span4Mux_v I__4383 (
            .O(N__19668),
            .I(N__19615));
    Span4Mux_h I__4382 (
            .O(N__19661),
            .I(N__19615));
    LocalMux I__4381 (
            .O(N__19658),
            .I(N__19615));
    IoInMux I__4380 (
            .O(N__19657),
            .I(N__19612));
    IoInMux I__4379 (
            .O(N__19656),
            .I(N__19609));
    LocalMux I__4378 (
            .O(N__19653),
            .I(N__19606));
    SRMux I__4377 (
            .O(N__19652),
            .I(N__19603));
    Span4Mux_s3_v I__4376 (
            .O(N__19649),
            .I(N__19595));
    LocalMux I__4375 (
            .O(N__19646),
            .I(N__19595));
    LocalMux I__4374 (
            .O(N__19643),
            .I(N__19595));
    Span4Mux_v I__4373 (
            .O(N__19636),
            .I(N__19588));
    Span4Mux_h I__4372 (
            .O(N__19633),
            .I(N__19588));
    LocalMux I__4371 (
            .O(N__19630),
            .I(N__19588));
    SRMux I__4370 (
            .O(N__19629),
            .I(N__19585));
    Span4Mux_v I__4369 (
            .O(N__19622),
            .I(N__19580));
    Span4Mux_v I__4368 (
            .O(N__19615),
            .I(N__19580));
    LocalMux I__4367 (
            .O(N__19612),
            .I(N__19575));
    LocalMux I__4366 (
            .O(N__19609),
            .I(N__19575));
    Span12Mux_s9_h I__4365 (
            .O(N__19606),
            .I(N__19572));
    LocalMux I__4364 (
            .O(N__19603),
            .I(N__19569));
    SRMux I__4363 (
            .O(N__19602),
            .I(N__19566));
    Span4Mux_v I__4362 (
            .O(N__19595),
            .I(N__19563));
    Span4Mux_v I__4361 (
            .O(N__19588),
            .I(N__19558));
    LocalMux I__4360 (
            .O(N__19585),
            .I(N__19558));
    Span4Mux_h I__4359 (
            .O(N__19580),
            .I(N__19555));
    Span4Mux_s3_v I__4358 (
            .O(N__19575),
            .I(N__19552));
    Span12Mux_v I__4357 (
            .O(N__19572),
            .I(N__19547));
    Span12Mux_s9_h I__4356 (
            .O(N__19569),
            .I(N__19547));
    LocalMux I__4355 (
            .O(N__19566),
            .I(N__19544));
    Span4Mux_h I__4354 (
            .O(N__19563),
            .I(N__19539));
    Span4Mux_h I__4353 (
            .O(N__19558),
            .I(N__19539));
    Span4Mux_h I__4352 (
            .O(N__19555),
            .I(N__19534));
    Span4Mux_v I__4351 (
            .O(N__19552),
            .I(N__19534));
    Span12Mux_v I__4350 (
            .O(N__19547),
            .I(N__19529));
    Span12Mux_s9_h I__4349 (
            .O(N__19544),
            .I(N__19529));
    Span4Mux_h I__4348 (
            .O(N__19539),
            .I(N__19526));
    Odrv4 I__4347 (
            .O(N__19534),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__4346 (
            .O(N__19529),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__4345 (
            .O(N__19526),
            .I(CONSTANT_ONE_NET));
    InMux I__4344 (
            .O(N__19519),
            .I(N__19516));
    LocalMux I__4343 (
            .O(N__19516),
            .I(N__19513));
    Span4Mux_h I__4342 (
            .O(N__19513),
            .I(N__19510));
    Span4Mux_h I__4341 (
            .O(N__19510),
            .I(N__19507));
    Odrv4 I__4340 (
            .O(N__19507),
            .I(\transmit_module.Y_DELTA_PATTERN_33 ));
    InMux I__4339 (
            .O(N__19504),
            .I(N__19501));
    LocalMux I__4338 (
            .O(N__19501),
            .I(N__19498));
    Odrv4 I__4337 (
            .O(N__19498),
            .I(\transmit_module.Y_DELTA_PATTERN_27 ));
    InMux I__4336 (
            .O(N__19495),
            .I(N__19492));
    LocalMux I__4335 (
            .O(N__19492),
            .I(\transmit_module.Y_DELTA_PATTERN_28 ));
    InMux I__4334 (
            .O(N__19489),
            .I(N__19486));
    LocalMux I__4333 (
            .O(N__19486),
            .I(\transmit_module.Y_DELTA_PATTERN_29 ));
    InMux I__4332 (
            .O(N__19483),
            .I(N__19480));
    LocalMux I__4331 (
            .O(N__19480),
            .I(\transmit_module.Y_DELTA_PATTERN_30 ));
    InMux I__4330 (
            .O(N__19477),
            .I(N__19474));
    LocalMux I__4329 (
            .O(N__19474),
            .I(\transmit_module.Y_DELTA_PATTERN_12 ));
    InMux I__4328 (
            .O(N__19471),
            .I(N__19468));
    LocalMux I__4327 (
            .O(N__19468),
            .I(N__19465));
    Span4Mux_h I__4326 (
            .O(N__19465),
            .I(N__19462));
    Odrv4 I__4325 (
            .O(N__19462),
            .I(\transmit_module.Y_DELTA_PATTERN_11 ));
    InMux I__4324 (
            .O(N__19459),
            .I(N__19456));
    LocalMux I__4323 (
            .O(N__19456),
            .I(\transmit_module.Y_DELTA_PATTERN_25 ));
    InMux I__4322 (
            .O(N__19453),
            .I(N__19450));
    LocalMux I__4321 (
            .O(N__19450),
            .I(\transmit_module.Y_DELTA_PATTERN_26 ));
    InMux I__4320 (
            .O(N__19447),
            .I(N__19444));
    LocalMux I__4319 (
            .O(N__19444),
            .I(\transmit_module.Y_DELTA_PATTERN_13 ));
    InMux I__4318 (
            .O(N__19441),
            .I(N__19438));
    LocalMux I__4317 (
            .O(N__19438),
            .I(N__19435));
    Span12Mux_h I__4316 (
            .O(N__19435),
            .I(N__19432));
    Odrv12 I__4315 (
            .O(N__19432),
            .I(\line_buffer.n539 ));
    InMux I__4314 (
            .O(N__19429),
            .I(N__19426));
    LocalMux I__4313 (
            .O(N__19426),
            .I(N__19423));
    Span4Mux_h I__4312 (
            .O(N__19423),
            .I(N__19420));
    Span4Mux_h I__4311 (
            .O(N__19420),
            .I(N__19417));
    Odrv4 I__4310 (
            .O(N__19417),
            .I(\line_buffer.n531 ));
    InMux I__4309 (
            .O(N__19414),
            .I(N__19411));
    LocalMux I__4308 (
            .O(N__19411),
            .I(\line_buffer.n3746 ));
    InMux I__4307 (
            .O(N__19408),
            .I(N__19405));
    LocalMux I__4306 (
            .O(N__19405),
            .I(N__19402));
    Span4Mux_v I__4305 (
            .O(N__19402),
            .I(N__19399));
    Sp12to4 I__4304 (
            .O(N__19399),
            .I(N__19396));
    Odrv12 I__4303 (
            .O(N__19396),
            .I(\line_buffer.n573 ));
    InMux I__4302 (
            .O(N__19393),
            .I(N__19390));
    LocalMux I__4301 (
            .O(N__19390),
            .I(N__19387));
    Sp12to4 I__4300 (
            .O(N__19387),
            .I(N__19384));
    Span12Mux_v I__4299 (
            .O(N__19384),
            .I(N__19381));
    Odrv12 I__4298 (
            .O(N__19381),
            .I(\line_buffer.n565 ));
    InMux I__4297 (
            .O(N__19378),
            .I(N__19375));
    LocalMux I__4296 (
            .O(N__19375),
            .I(\line_buffer.n3677 ));
    InMux I__4295 (
            .O(N__19372),
            .I(N__19369));
    LocalMux I__4294 (
            .O(N__19369),
            .I(N__19366));
    Span12Mux_v I__4293 (
            .O(N__19366),
            .I(N__19363));
    Odrv12 I__4292 (
            .O(N__19363),
            .I(\line_buffer.n567 ));
    InMux I__4291 (
            .O(N__19360),
            .I(N__19357));
    LocalMux I__4290 (
            .O(N__19357),
            .I(N__19354));
    Span4Mux_v I__4289 (
            .O(N__19354),
            .I(N__19351));
    Sp12to4 I__4288 (
            .O(N__19351),
            .I(N__19348));
    Odrv12 I__4287 (
            .O(N__19348),
            .I(\line_buffer.n575 ));
    InMux I__4286 (
            .O(N__19345),
            .I(N__19342));
    LocalMux I__4285 (
            .O(N__19342),
            .I(\line_buffer.n3635 ));
    InMux I__4284 (
            .O(N__19339),
            .I(N__19334));
    InMux I__4283 (
            .O(N__19338),
            .I(N__19329));
    InMux I__4282 (
            .O(N__19337),
            .I(N__19329));
    LocalMux I__4281 (
            .O(N__19334),
            .I(\receive_module.rx_counter.X_4 ));
    LocalMux I__4280 (
            .O(N__19329),
            .I(\receive_module.rx_counter.X_4 ));
    InMux I__4279 (
            .O(N__19324),
            .I(\receive_module.rx_counter.n3304 ));
    InMux I__4278 (
            .O(N__19321),
            .I(N__19316));
    InMux I__4277 (
            .O(N__19320),
            .I(N__19311));
    InMux I__4276 (
            .O(N__19319),
            .I(N__19311));
    LocalMux I__4275 (
            .O(N__19316),
            .I(\receive_module.rx_counter.X_5 ));
    LocalMux I__4274 (
            .O(N__19311),
            .I(\receive_module.rx_counter.X_5 ));
    InMux I__4273 (
            .O(N__19306),
            .I(\receive_module.rx_counter.n3305 ));
    InMux I__4272 (
            .O(N__19303),
            .I(N__19298));
    InMux I__4271 (
            .O(N__19302),
            .I(N__19293));
    InMux I__4270 (
            .O(N__19301),
            .I(N__19293));
    LocalMux I__4269 (
            .O(N__19298),
            .I(\receive_module.rx_counter.X_6 ));
    LocalMux I__4268 (
            .O(N__19293),
            .I(\receive_module.rx_counter.X_6 ));
    InMux I__4267 (
            .O(N__19288),
            .I(\receive_module.rx_counter.n3306 ));
    InMux I__4266 (
            .O(N__19285),
            .I(N__19280));
    InMux I__4265 (
            .O(N__19284),
            .I(N__19275));
    InMux I__4264 (
            .O(N__19283),
            .I(N__19275));
    LocalMux I__4263 (
            .O(N__19280),
            .I(\receive_module.rx_counter.X_7 ));
    LocalMux I__4262 (
            .O(N__19275),
            .I(\receive_module.rx_counter.X_7 ));
    InMux I__4261 (
            .O(N__19270),
            .I(\receive_module.rx_counter.n3307 ));
    InMux I__4260 (
            .O(N__19267),
            .I(N__19263));
    InMux I__4259 (
            .O(N__19266),
            .I(N__19260));
    LocalMux I__4258 (
            .O(N__19263),
            .I(\receive_module.rx_counter.X_8 ));
    LocalMux I__4257 (
            .O(N__19260),
            .I(\receive_module.rx_counter.X_8 ));
    InMux I__4256 (
            .O(N__19255),
            .I(bfn_17_11_0_));
    InMux I__4255 (
            .O(N__19252),
            .I(\receive_module.rx_counter.n3309 ));
    CascadeMux I__4254 (
            .O(N__19249),
            .I(N__19245));
    InMux I__4253 (
            .O(N__19248),
            .I(N__19242));
    InMux I__4252 (
            .O(N__19245),
            .I(N__19239));
    LocalMux I__4251 (
            .O(N__19242),
            .I(\receive_module.rx_counter.X_9 ));
    LocalMux I__4250 (
            .O(N__19239),
            .I(\receive_module.rx_counter.X_9 ));
    SRMux I__4249 (
            .O(N__19234),
            .I(N__19230));
    SRMux I__4248 (
            .O(N__19233),
            .I(N__19227));
    LocalMux I__4247 (
            .O(N__19230),
            .I(N__19224));
    LocalMux I__4246 (
            .O(N__19227),
            .I(N__19221));
    Span4Mux_h I__4245 (
            .O(N__19224),
            .I(N__19218));
    Odrv4 I__4244 (
            .O(N__19221),
            .I(\receive_module.rx_counter.n3790 ));
    Odrv4 I__4243 (
            .O(N__19218),
            .I(\receive_module.rx_counter.n3790 ));
    InMux I__4242 (
            .O(N__19213),
            .I(N__19210));
    LocalMux I__4241 (
            .O(N__19210),
            .I(N__19207));
    Odrv12 I__4240 (
            .O(N__19207),
            .I(\line_buffer.n576 ));
    InMux I__4239 (
            .O(N__19204),
            .I(N__19201));
    LocalMux I__4238 (
            .O(N__19201),
            .I(N__19198));
    Span12Mux_v I__4237 (
            .O(N__19198),
            .I(N__19195));
    Span12Mux_v I__4236 (
            .O(N__19195),
            .I(N__19192));
    Odrv12 I__4235 (
            .O(N__19192),
            .I(\line_buffer.n568 ));
    InMux I__4234 (
            .O(N__19189),
            .I(N__19186));
    LocalMux I__4233 (
            .O(N__19186),
            .I(N__19183));
    Sp12to4 I__4232 (
            .O(N__19183),
            .I(N__19180));
    Span12Mux_v I__4231 (
            .O(N__19180),
            .I(N__19177));
    Odrv12 I__4230 (
            .O(N__19177),
            .I(\line_buffer.n504 ));
    InMux I__4229 (
            .O(N__19174),
            .I(N__19171));
    LocalMux I__4228 (
            .O(N__19171),
            .I(N__19168));
    Span12Mux_h I__4227 (
            .O(N__19168),
            .I(N__19165));
    Span12Mux_v I__4226 (
            .O(N__19165),
            .I(N__19162));
    Odrv12 I__4225 (
            .O(N__19162),
            .I(\line_buffer.n512 ));
    CascadeMux I__4224 (
            .O(N__19159),
            .I(\line_buffer.n3734_cascade_ ));
    InMux I__4223 (
            .O(N__19156),
            .I(N__19153));
    LocalMux I__4222 (
            .O(N__19153),
            .I(N__19150));
    Span4Mux_v I__4221 (
            .O(N__19150),
            .I(N__19147));
    Sp12to4 I__4220 (
            .O(N__19147),
            .I(N__19144));
    Odrv12 I__4219 (
            .O(N__19144),
            .I(\line_buffer.n444 ));
    InMux I__4218 (
            .O(N__19141),
            .I(N__19138));
    LocalMux I__4217 (
            .O(N__19138),
            .I(N__19135));
    Span4Mux_v I__4216 (
            .O(N__19135),
            .I(N__19132));
    Sp12to4 I__4215 (
            .O(N__19132),
            .I(N__19129));
    Span12Mux_h I__4214 (
            .O(N__19129),
            .I(N__19126));
    Odrv12 I__4213 (
            .O(N__19126),
            .I(\line_buffer.n436 ));
    InMux I__4212 (
            .O(N__19123),
            .I(N__19120));
    LocalMux I__4211 (
            .O(N__19120),
            .I(N__19117));
    Odrv12 I__4210 (
            .O(N__19117),
            .I(\line_buffer.n3673 ));
    InMux I__4209 (
            .O(N__19114),
            .I(N__19110));
    InMux I__4208 (
            .O(N__19113),
            .I(N__19106));
    LocalMux I__4207 (
            .O(N__19110),
            .I(N__19103));
    InMux I__4206 (
            .O(N__19109),
            .I(N__19100));
    LocalMux I__4205 (
            .O(N__19106),
            .I(N__19094));
    Span4Mux_h I__4204 (
            .O(N__19103),
            .I(N__19090));
    LocalMux I__4203 (
            .O(N__19100),
            .I(N__19087));
    CascadeMux I__4202 (
            .O(N__19099),
            .I(N__19083));
    InMux I__4201 (
            .O(N__19098),
            .I(N__19072));
    InMux I__4200 (
            .O(N__19097),
            .I(N__19072));
    Span4Mux_h I__4199 (
            .O(N__19094),
            .I(N__19069));
    InMux I__4198 (
            .O(N__19093),
            .I(N__19061));
    Span4Mux_v I__4197 (
            .O(N__19090),
            .I(N__19054));
    Span4Mux_h I__4196 (
            .O(N__19087),
            .I(N__19054));
    InMux I__4195 (
            .O(N__19086),
            .I(N__19051));
    InMux I__4194 (
            .O(N__19083),
            .I(N__19048));
    InMux I__4193 (
            .O(N__19082),
            .I(N__19043));
    InMux I__4192 (
            .O(N__19081),
            .I(N__19043));
    InMux I__4191 (
            .O(N__19080),
            .I(N__19034));
    InMux I__4190 (
            .O(N__19079),
            .I(N__19034));
    InMux I__4189 (
            .O(N__19078),
            .I(N__19034));
    InMux I__4188 (
            .O(N__19077),
            .I(N__19034));
    LocalMux I__4187 (
            .O(N__19072),
            .I(N__19031));
    Span4Mux_v I__4186 (
            .O(N__19069),
            .I(N__19028));
    InMux I__4185 (
            .O(N__19068),
            .I(N__19025));
    InMux I__4184 (
            .O(N__19067),
            .I(N__19019));
    InMux I__4183 (
            .O(N__19066),
            .I(N__19014));
    InMux I__4182 (
            .O(N__19065),
            .I(N__19014));
    InMux I__4181 (
            .O(N__19064),
            .I(N__19011));
    LocalMux I__4180 (
            .O(N__19061),
            .I(N__19008));
    InMux I__4179 (
            .O(N__19060),
            .I(N__19003));
    InMux I__4178 (
            .O(N__19059),
            .I(N__19003));
    Span4Mux_v I__4177 (
            .O(N__19054),
            .I(N__18998));
    LocalMux I__4176 (
            .O(N__19051),
            .I(N__18998));
    LocalMux I__4175 (
            .O(N__19048),
            .I(N__18993));
    LocalMux I__4174 (
            .O(N__19043),
            .I(N__18993));
    LocalMux I__4173 (
            .O(N__19034),
            .I(N__18990));
    Span4Mux_h I__4172 (
            .O(N__19031),
            .I(N__18982));
    Span4Mux_v I__4171 (
            .O(N__19028),
            .I(N__18982));
    LocalMux I__4170 (
            .O(N__19025),
            .I(N__18979));
    InMux I__4169 (
            .O(N__19024),
            .I(N__18976));
    InMux I__4168 (
            .O(N__19023),
            .I(N__18971));
    InMux I__4167 (
            .O(N__19022),
            .I(N__18971));
    LocalMux I__4166 (
            .O(N__19019),
            .I(N__18966));
    LocalMux I__4165 (
            .O(N__19014),
            .I(N__18966));
    LocalMux I__4164 (
            .O(N__19011),
            .I(N__18957));
    Span4Mux_h I__4163 (
            .O(N__19008),
            .I(N__18957));
    LocalMux I__4162 (
            .O(N__19003),
            .I(N__18957));
    Span4Mux_v I__4161 (
            .O(N__18998),
            .I(N__18957));
    Span4Mux_v I__4160 (
            .O(N__18993),
            .I(N__18954));
    Span4Mux_h I__4159 (
            .O(N__18990),
            .I(N__18951));
    InMux I__4158 (
            .O(N__18989),
            .I(N__18948));
    InMux I__4157 (
            .O(N__18988),
            .I(N__18943));
    InMux I__4156 (
            .O(N__18987),
            .I(N__18943));
    Span4Mux_v I__4155 (
            .O(N__18982),
            .I(N__18940));
    Span4Mux_v I__4154 (
            .O(N__18979),
            .I(N__18929));
    LocalMux I__4153 (
            .O(N__18976),
            .I(N__18929));
    LocalMux I__4152 (
            .O(N__18971),
            .I(N__18929));
    Span4Mux_h I__4151 (
            .O(N__18966),
            .I(N__18929));
    Span4Mux_v I__4150 (
            .O(N__18957),
            .I(N__18929));
    Odrv4 I__4149 (
            .O(N__18954),
            .I(\transmit_module.n3787 ));
    Odrv4 I__4148 (
            .O(N__18951),
            .I(\transmit_module.n3787 ));
    LocalMux I__4147 (
            .O(N__18948),
            .I(\transmit_module.n3787 ));
    LocalMux I__4146 (
            .O(N__18943),
            .I(\transmit_module.n3787 ));
    Odrv4 I__4145 (
            .O(N__18940),
            .I(\transmit_module.n3787 ));
    Odrv4 I__4144 (
            .O(N__18929),
            .I(\transmit_module.n3787 ));
    InMux I__4143 (
            .O(N__18916),
            .I(N__18913));
    LocalMux I__4142 (
            .O(N__18913),
            .I(N__18909));
    InMux I__4141 (
            .O(N__18912),
            .I(N__18906));
    Span12Mux_v I__4140 (
            .O(N__18909),
            .I(N__18903));
    LocalMux I__4139 (
            .O(N__18906),
            .I(\transmit_module.n108 ));
    Odrv12 I__4138 (
            .O(N__18903),
            .I(\transmit_module.n108 ));
    InMux I__4137 (
            .O(N__18898),
            .I(N__18895));
    LocalMux I__4136 (
            .O(N__18895),
            .I(N__18892));
    Odrv12 I__4135 (
            .O(N__18892),
            .I(\transmit_module.n139 ));
    CascadeMux I__4134 (
            .O(N__18889),
            .I(N__18886));
    CascadeBuf I__4133 (
            .O(N__18886),
            .I(N__18882));
    CascadeMux I__4132 (
            .O(N__18885),
            .I(N__18879));
    CascadeMux I__4131 (
            .O(N__18882),
            .I(N__18876));
    CascadeBuf I__4130 (
            .O(N__18879),
            .I(N__18873));
    CascadeBuf I__4129 (
            .O(N__18876),
            .I(N__18870));
    CascadeMux I__4128 (
            .O(N__18873),
            .I(N__18867));
    CascadeMux I__4127 (
            .O(N__18870),
            .I(N__18864));
    CascadeBuf I__4126 (
            .O(N__18867),
            .I(N__18861));
    CascadeBuf I__4125 (
            .O(N__18864),
            .I(N__18858));
    CascadeMux I__4124 (
            .O(N__18861),
            .I(N__18855));
    CascadeMux I__4123 (
            .O(N__18858),
            .I(N__18852));
    CascadeBuf I__4122 (
            .O(N__18855),
            .I(N__18849));
    CascadeBuf I__4121 (
            .O(N__18852),
            .I(N__18846));
    CascadeMux I__4120 (
            .O(N__18849),
            .I(N__18843));
    CascadeMux I__4119 (
            .O(N__18846),
            .I(N__18840));
    CascadeBuf I__4118 (
            .O(N__18843),
            .I(N__18837));
    CascadeBuf I__4117 (
            .O(N__18840),
            .I(N__18834));
    CascadeMux I__4116 (
            .O(N__18837),
            .I(N__18831));
    CascadeMux I__4115 (
            .O(N__18834),
            .I(N__18828));
    CascadeBuf I__4114 (
            .O(N__18831),
            .I(N__18825));
    CascadeBuf I__4113 (
            .O(N__18828),
            .I(N__18822));
    CascadeMux I__4112 (
            .O(N__18825),
            .I(N__18819));
    CascadeMux I__4111 (
            .O(N__18822),
            .I(N__18816));
    CascadeBuf I__4110 (
            .O(N__18819),
            .I(N__18813));
    CascadeBuf I__4109 (
            .O(N__18816),
            .I(N__18810));
    CascadeMux I__4108 (
            .O(N__18813),
            .I(N__18807));
    CascadeMux I__4107 (
            .O(N__18810),
            .I(N__18804));
    CascadeBuf I__4106 (
            .O(N__18807),
            .I(N__18801));
    CascadeBuf I__4105 (
            .O(N__18804),
            .I(N__18798));
    CascadeMux I__4104 (
            .O(N__18801),
            .I(N__18795));
    CascadeMux I__4103 (
            .O(N__18798),
            .I(N__18792));
    CascadeBuf I__4102 (
            .O(N__18795),
            .I(N__18789));
    CascadeBuf I__4101 (
            .O(N__18792),
            .I(N__18786));
    CascadeMux I__4100 (
            .O(N__18789),
            .I(N__18783));
    CascadeMux I__4099 (
            .O(N__18786),
            .I(N__18780));
    CascadeBuf I__4098 (
            .O(N__18783),
            .I(N__18777));
    CascadeBuf I__4097 (
            .O(N__18780),
            .I(N__18774));
    CascadeMux I__4096 (
            .O(N__18777),
            .I(N__18771));
    CascadeMux I__4095 (
            .O(N__18774),
            .I(N__18768));
    CascadeBuf I__4094 (
            .O(N__18771),
            .I(N__18765));
    CascadeBuf I__4093 (
            .O(N__18768),
            .I(N__18762));
    CascadeMux I__4092 (
            .O(N__18765),
            .I(N__18759));
    CascadeMux I__4091 (
            .O(N__18762),
            .I(N__18756));
    CascadeBuf I__4090 (
            .O(N__18759),
            .I(N__18753));
    CascadeBuf I__4089 (
            .O(N__18756),
            .I(N__18750));
    CascadeMux I__4088 (
            .O(N__18753),
            .I(N__18747));
    CascadeMux I__4087 (
            .O(N__18750),
            .I(N__18744));
    CascadeBuf I__4086 (
            .O(N__18747),
            .I(N__18741));
    CascadeBuf I__4085 (
            .O(N__18744),
            .I(N__18738));
    CascadeMux I__4084 (
            .O(N__18741),
            .I(N__18735));
    CascadeMux I__4083 (
            .O(N__18738),
            .I(N__18732));
    CascadeBuf I__4082 (
            .O(N__18735),
            .I(N__18729));
    CascadeBuf I__4081 (
            .O(N__18732),
            .I(N__18726));
    CascadeMux I__4080 (
            .O(N__18729),
            .I(N__18723));
    CascadeMux I__4079 (
            .O(N__18726),
            .I(N__18720));
    CascadeBuf I__4078 (
            .O(N__18723),
            .I(N__18717));
    CascadeBuf I__4077 (
            .O(N__18720),
            .I(N__18714));
    CascadeMux I__4076 (
            .O(N__18717),
            .I(N__18711));
    CascadeMux I__4075 (
            .O(N__18714),
            .I(N__18708));
    CascadeBuf I__4074 (
            .O(N__18711),
            .I(N__18705));
    InMux I__4073 (
            .O(N__18708),
            .I(N__18702));
    CascadeMux I__4072 (
            .O(N__18705),
            .I(N__18699));
    LocalMux I__4071 (
            .O(N__18702),
            .I(N__18696));
    InMux I__4070 (
            .O(N__18699),
            .I(N__18693));
    Span4Mux_s3_v I__4069 (
            .O(N__18696),
            .I(N__18690));
    LocalMux I__4068 (
            .O(N__18693),
            .I(N__18687));
    Span4Mux_v I__4067 (
            .O(N__18690),
            .I(N__18684));
    Span4Mux_h I__4066 (
            .O(N__18687),
            .I(N__18681));
    Span4Mux_h I__4065 (
            .O(N__18684),
            .I(N__18678));
    Span4Mux_h I__4064 (
            .O(N__18681),
            .I(N__18675));
    Span4Mux_h I__4063 (
            .O(N__18678),
            .I(N__18672));
    Sp12to4 I__4062 (
            .O(N__18675),
            .I(N__18669));
    Odrv4 I__4061 (
            .O(N__18672),
            .I(n20));
    Odrv12 I__4060 (
            .O(N__18669),
            .I(n20));
    IoInMux I__4059 (
            .O(N__18664),
            .I(N__18661));
    LocalMux I__4058 (
            .O(N__18661),
            .I(N__18658));
    Span4Mux_s0_v I__4057 (
            .O(N__18658),
            .I(N__18655));
    Odrv4 I__4056 (
            .O(N__18655),
            .I(GB_BUFFER_TVP_CLK_c_THRU_CO));
    InMux I__4055 (
            .O(N__18652),
            .I(N__18646));
    InMux I__4054 (
            .O(N__18651),
            .I(N__18646));
    LocalMux I__4053 (
            .O(N__18646),
            .I(N__18642));
    InMux I__4052 (
            .O(N__18645),
            .I(N__18639));
    Span4Mux_v I__4051 (
            .O(N__18642),
            .I(N__18636));
    LocalMux I__4050 (
            .O(N__18639),
            .I(N__18633));
    Span4Mux_h I__4049 (
            .O(N__18636),
            .I(N__18628));
    Span4Mux_h I__4048 (
            .O(N__18633),
            .I(N__18628));
    Sp12to4 I__4047 (
            .O(N__18628),
            .I(N__18625));
    Odrv12 I__4046 (
            .O(N__18625),
            .I(TVP_HSYNC_c));
    InMux I__4045 (
            .O(N__18622),
            .I(N__18619));
    LocalMux I__4044 (
            .O(N__18619),
            .I(\receive_module.rx_counter.n10 ));
    InMux I__4043 (
            .O(N__18616),
            .I(bfn_17_10_0_));
    InMux I__4042 (
            .O(N__18613),
            .I(N__18610));
    LocalMux I__4041 (
            .O(N__18610),
            .I(\receive_module.rx_counter.n9 ));
    InMux I__4040 (
            .O(N__18607),
            .I(\receive_module.rx_counter.n3301 ));
    InMux I__4039 (
            .O(N__18604),
            .I(N__18601));
    LocalMux I__4038 (
            .O(N__18601),
            .I(\receive_module.rx_counter.n8 ));
    InMux I__4037 (
            .O(N__18598),
            .I(\receive_module.rx_counter.n3302 ));
    InMux I__4036 (
            .O(N__18595),
            .I(N__18590));
    InMux I__4035 (
            .O(N__18594),
            .I(N__18585));
    InMux I__4034 (
            .O(N__18593),
            .I(N__18585));
    LocalMux I__4033 (
            .O(N__18590),
            .I(\receive_module.rx_counter.X_3 ));
    LocalMux I__4032 (
            .O(N__18585),
            .I(\receive_module.rx_counter.X_3 ));
    InMux I__4031 (
            .O(N__18580),
            .I(\receive_module.rx_counter.n3303 ));
    InMux I__4030 (
            .O(N__18577),
            .I(N__18574));
    LocalMux I__4029 (
            .O(N__18574),
            .I(N__18571));
    Span4Mux_h I__4028 (
            .O(N__18571),
            .I(N__18568));
    Span4Mux_v I__4027 (
            .O(N__18568),
            .I(N__18564));
    InMux I__4026 (
            .O(N__18567),
            .I(N__18561));
    Odrv4 I__4025 (
            .O(N__18564),
            .I(\transmit_module.n114 ));
    LocalMux I__4024 (
            .O(N__18561),
            .I(\transmit_module.n114 ));
    InMux I__4023 (
            .O(N__18556),
            .I(N__18553));
    LocalMux I__4022 (
            .O(N__18553),
            .I(N__18550));
    Span4Mux_h I__4021 (
            .O(N__18550),
            .I(N__18546));
    InMux I__4020 (
            .O(N__18549),
            .I(N__18543));
    Odrv4 I__4019 (
            .O(N__18546),
            .I(\transmit_module.n145 ));
    LocalMux I__4018 (
            .O(N__18543),
            .I(\transmit_module.n145 ));
    CascadeMux I__4017 (
            .O(N__18538),
            .I(N__18535));
    CascadeBuf I__4016 (
            .O(N__18535),
            .I(N__18531));
    CascadeMux I__4015 (
            .O(N__18534),
            .I(N__18528));
    CascadeMux I__4014 (
            .O(N__18531),
            .I(N__18525));
    CascadeBuf I__4013 (
            .O(N__18528),
            .I(N__18522));
    CascadeBuf I__4012 (
            .O(N__18525),
            .I(N__18519));
    CascadeMux I__4011 (
            .O(N__18522),
            .I(N__18516));
    CascadeMux I__4010 (
            .O(N__18519),
            .I(N__18513));
    CascadeBuf I__4009 (
            .O(N__18516),
            .I(N__18510));
    CascadeBuf I__4008 (
            .O(N__18513),
            .I(N__18507));
    CascadeMux I__4007 (
            .O(N__18510),
            .I(N__18504));
    CascadeMux I__4006 (
            .O(N__18507),
            .I(N__18501));
    CascadeBuf I__4005 (
            .O(N__18504),
            .I(N__18498));
    CascadeBuf I__4004 (
            .O(N__18501),
            .I(N__18495));
    CascadeMux I__4003 (
            .O(N__18498),
            .I(N__18492));
    CascadeMux I__4002 (
            .O(N__18495),
            .I(N__18489));
    CascadeBuf I__4001 (
            .O(N__18492),
            .I(N__18486));
    CascadeBuf I__4000 (
            .O(N__18489),
            .I(N__18483));
    CascadeMux I__3999 (
            .O(N__18486),
            .I(N__18480));
    CascadeMux I__3998 (
            .O(N__18483),
            .I(N__18477));
    CascadeBuf I__3997 (
            .O(N__18480),
            .I(N__18474));
    CascadeBuf I__3996 (
            .O(N__18477),
            .I(N__18471));
    CascadeMux I__3995 (
            .O(N__18474),
            .I(N__18468));
    CascadeMux I__3994 (
            .O(N__18471),
            .I(N__18465));
    CascadeBuf I__3993 (
            .O(N__18468),
            .I(N__18462));
    CascadeBuf I__3992 (
            .O(N__18465),
            .I(N__18459));
    CascadeMux I__3991 (
            .O(N__18462),
            .I(N__18456));
    CascadeMux I__3990 (
            .O(N__18459),
            .I(N__18453));
    CascadeBuf I__3989 (
            .O(N__18456),
            .I(N__18450));
    CascadeBuf I__3988 (
            .O(N__18453),
            .I(N__18447));
    CascadeMux I__3987 (
            .O(N__18450),
            .I(N__18444));
    CascadeMux I__3986 (
            .O(N__18447),
            .I(N__18441));
    CascadeBuf I__3985 (
            .O(N__18444),
            .I(N__18438));
    CascadeBuf I__3984 (
            .O(N__18441),
            .I(N__18435));
    CascadeMux I__3983 (
            .O(N__18438),
            .I(N__18432));
    CascadeMux I__3982 (
            .O(N__18435),
            .I(N__18429));
    CascadeBuf I__3981 (
            .O(N__18432),
            .I(N__18426));
    CascadeBuf I__3980 (
            .O(N__18429),
            .I(N__18423));
    CascadeMux I__3979 (
            .O(N__18426),
            .I(N__18420));
    CascadeMux I__3978 (
            .O(N__18423),
            .I(N__18417));
    CascadeBuf I__3977 (
            .O(N__18420),
            .I(N__18414));
    CascadeBuf I__3976 (
            .O(N__18417),
            .I(N__18411));
    CascadeMux I__3975 (
            .O(N__18414),
            .I(N__18408));
    CascadeMux I__3974 (
            .O(N__18411),
            .I(N__18405));
    CascadeBuf I__3973 (
            .O(N__18408),
            .I(N__18402));
    CascadeBuf I__3972 (
            .O(N__18405),
            .I(N__18399));
    CascadeMux I__3971 (
            .O(N__18402),
            .I(N__18396));
    CascadeMux I__3970 (
            .O(N__18399),
            .I(N__18393));
    CascadeBuf I__3969 (
            .O(N__18396),
            .I(N__18390));
    CascadeBuf I__3968 (
            .O(N__18393),
            .I(N__18387));
    CascadeMux I__3967 (
            .O(N__18390),
            .I(N__18384));
    CascadeMux I__3966 (
            .O(N__18387),
            .I(N__18381));
    CascadeBuf I__3965 (
            .O(N__18384),
            .I(N__18378));
    CascadeBuf I__3964 (
            .O(N__18381),
            .I(N__18375));
    CascadeMux I__3963 (
            .O(N__18378),
            .I(N__18372));
    CascadeMux I__3962 (
            .O(N__18375),
            .I(N__18369));
    CascadeBuf I__3961 (
            .O(N__18372),
            .I(N__18366));
    CascadeBuf I__3960 (
            .O(N__18369),
            .I(N__18363));
    CascadeMux I__3959 (
            .O(N__18366),
            .I(N__18360));
    CascadeMux I__3958 (
            .O(N__18363),
            .I(N__18357));
    CascadeBuf I__3957 (
            .O(N__18360),
            .I(N__18354));
    InMux I__3956 (
            .O(N__18357),
            .I(N__18351));
    CascadeMux I__3955 (
            .O(N__18354),
            .I(N__18348));
    LocalMux I__3954 (
            .O(N__18351),
            .I(N__18345));
    InMux I__3953 (
            .O(N__18348),
            .I(N__18342));
    Span4Mux_v I__3952 (
            .O(N__18345),
            .I(N__18339));
    LocalMux I__3951 (
            .O(N__18342),
            .I(N__18336));
    Span4Mux_v I__3950 (
            .O(N__18339),
            .I(N__18333));
    Span4Mux_h I__3949 (
            .O(N__18336),
            .I(N__18330));
    Span4Mux_v I__3948 (
            .O(N__18333),
            .I(N__18327));
    Sp12to4 I__3947 (
            .O(N__18330),
            .I(N__18324));
    Sp12to4 I__3946 (
            .O(N__18327),
            .I(N__18319));
    Span12Mux_v I__3945 (
            .O(N__18324),
            .I(N__18319));
    Odrv12 I__3944 (
            .O(N__18319),
            .I(n26));
    InMux I__3943 (
            .O(N__18316),
            .I(N__18311));
    InMux I__3942 (
            .O(N__18315),
            .I(N__18308));
    InMux I__3941 (
            .O(N__18314),
            .I(N__18304));
    LocalMux I__3940 (
            .O(N__18311),
            .I(N__18295));
    LocalMux I__3939 (
            .O(N__18308),
            .I(N__18291));
    InMux I__3938 (
            .O(N__18307),
            .I(N__18288));
    LocalMux I__3937 (
            .O(N__18304),
            .I(N__18285));
    InMux I__3936 (
            .O(N__18303),
            .I(N__18280));
    InMux I__3935 (
            .O(N__18302),
            .I(N__18280));
    InMux I__3934 (
            .O(N__18301),
            .I(N__18275));
    InMux I__3933 (
            .O(N__18300),
            .I(N__18275));
    CascadeMux I__3932 (
            .O(N__18299),
            .I(N__18270));
    InMux I__3931 (
            .O(N__18298),
            .I(N__18266));
    Span12Mux_h I__3930 (
            .O(N__18295),
            .I(N__18263));
    InMux I__3929 (
            .O(N__18294),
            .I(N__18260));
    Span4Mux_h I__3928 (
            .O(N__18291),
            .I(N__18257));
    LocalMux I__3927 (
            .O(N__18288),
            .I(N__18250));
    Span4Mux_v I__3926 (
            .O(N__18285),
            .I(N__18250));
    LocalMux I__3925 (
            .O(N__18280),
            .I(N__18250));
    LocalMux I__3924 (
            .O(N__18275),
            .I(N__18247));
    InMux I__3923 (
            .O(N__18274),
            .I(N__18242));
    InMux I__3922 (
            .O(N__18273),
            .I(N__18242));
    InMux I__3921 (
            .O(N__18270),
            .I(N__18237));
    InMux I__3920 (
            .O(N__18269),
            .I(N__18237));
    LocalMux I__3919 (
            .O(N__18266),
            .I(\transmit_module.VGA_VISIBLE ));
    Odrv12 I__3918 (
            .O(N__18263),
            .I(\transmit_module.VGA_VISIBLE ));
    LocalMux I__3917 (
            .O(N__18260),
            .I(\transmit_module.VGA_VISIBLE ));
    Odrv4 I__3916 (
            .O(N__18257),
            .I(\transmit_module.VGA_VISIBLE ));
    Odrv4 I__3915 (
            .O(N__18250),
            .I(\transmit_module.VGA_VISIBLE ));
    Odrv4 I__3914 (
            .O(N__18247),
            .I(\transmit_module.VGA_VISIBLE ));
    LocalMux I__3913 (
            .O(N__18242),
            .I(\transmit_module.VGA_VISIBLE ));
    LocalMux I__3912 (
            .O(N__18237),
            .I(\transmit_module.VGA_VISIBLE ));
    InMux I__3911 (
            .O(N__18220),
            .I(N__18217));
    LocalMux I__3910 (
            .O(N__18217),
            .I(N__18214));
    Span4Mux_v I__3909 (
            .O(N__18214),
            .I(N__18211));
    Odrv4 I__3908 (
            .O(N__18211),
            .I(\transmit_module.n129 ));
    InMux I__3907 (
            .O(N__18208),
            .I(N__18205));
    LocalMux I__3906 (
            .O(N__18205),
            .I(N__18202));
    Span4Mux_v I__3905 (
            .O(N__18202),
            .I(N__18199));
    Odrv4 I__3904 (
            .O(N__18199),
            .I(\transmit_module.n144 ));
    CascadeMux I__3903 (
            .O(N__18196),
            .I(\transmit_module.n144_cascade_ ));
    CascadeMux I__3902 (
            .O(N__18193),
            .I(N__18189));
    CascadeMux I__3901 (
            .O(N__18192),
            .I(N__18186));
    CascadeBuf I__3900 (
            .O(N__18189),
            .I(N__18183));
    CascadeBuf I__3899 (
            .O(N__18186),
            .I(N__18180));
    CascadeMux I__3898 (
            .O(N__18183),
            .I(N__18177));
    CascadeMux I__3897 (
            .O(N__18180),
            .I(N__18174));
    CascadeBuf I__3896 (
            .O(N__18177),
            .I(N__18171));
    CascadeBuf I__3895 (
            .O(N__18174),
            .I(N__18168));
    CascadeMux I__3894 (
            .O(N__18171),
            .I(N__18165));
    CascadeMux I__3893 (
            .O(N__18168),
            .I(N__18162));
    CascadeBuf I__3892 (
            .O(N__18165),
            .I(N__18159));
    CascadeBuf I__3891 (
            .O(N__18162),
            .I(N__18156));
    CascadeMux I__3890 (
            .O(N__18159),
            .I(N__18153));
    CascadeMux I__3889 (
            .O(N__18156),
            .I(N__18150));
    CascadeBuf I__3888 (
            .O(N__18153),
            .I(N__18147));
    CascadeBuf I__3887 (
            .O(N__18150),
            .I(N__18144));
    CascadeMux I__3886 (
            .O(N__18147),
            .I(N__18141));
    CascadeMux I__3885 (
            .O(N__18144),
            .I(N__18138));
    CascadeBuf I__3884 (
            .O(N__18141),
            .I(N__18135));
    CascadeBuf I__3883 (
            .O(N__18138),
            .I(N__18132));
    CascadeMux I__3882 (
            .O(N__18135),
            .I(N__18129));
    CascadeMux I__3881 (
            .O(N__18132),
            .I(N__18126));
    CascadeBuf I__3880 (
            .O(N__18129),
            .I(N__18123));
    CascadeBuf I__3879 (
            .O(N__18126),
            .I(N__18120));
    CascadeMux I__3878 (
            .O(N__18123),
            .I(N__18117));
    CascadeMux I__3877 (
            .O(N__18120),
            .I(N__18114));
    CascadeBuf I__3876 (
            .O(N__18117),
            .I(N__18111));
    CascadeBuf I__3875 (
            .O(N__18114),
            .I(N__18108));
    CascadeMux I__3874 (
            .O(N__18111),
            .I(N__18105));
    CascadeMux I__3873 (
            .O(N__18108),
            .I(N__18102));
    CascadeBuf I__3872 (
            .O(N__18105),
            .I(N__18099));
    CascadeBuf I__3871 (
            .O(N__18102),
            .I(N__18096));
    CascadeMux I__3870 (
            .O(N__18099),
            .I(N__18093));
    CascadeMux I__3869 (
            .O(N__18096),
            .I(N__18090));
    CascadeBuf I__3868 (
            .O(N__18093),
            .I(N__18087));
    CascadeBuf I__3867 (
            .O(N__18090),
            .I(N__18084));
    CascadeMux I__3866 (
            .O(N__18087),
            .I(N__18081));
    CascadeMux I__3865 (
            .O(N__18084),
            .I(N__18078));
    CascadeBuf I__3864 (
            .O(N__18081),
            .I(N__18075));
    CascadeBuf I__3863 (
            .O(N__18078),
            .I(N__18072));
    CascadeMux I__3862 (
            .O(N__18075),
            .I(N__18069));
    CascadeMux I__3861 (
            .O(N__18072),
            .I(N__18066));
    CascadeBuf I__3860 (
            .O(N__18069),
            .I(N__18063));
    CascadeBuf I__3859 (
            .O(N__18066),
            .I(N__18060));
    CascadeMux I__3858 (
            .O(N__18063),
            .I(N__18057));
    CascadeMux I__3857 (
            .O(N__18060),
            .I(N__18054));
    CascadeBuf I__3856 (
            .O(N__18057),
            .I(N__18051));
    CascadeBuf I__3855 (
            .O(N__18054),
            .I(N__18048));
    CascadeMux I__3854 (
            .O(N__18051),
            .I(N__18045));
    CascadeMux I__3853 (
            .O(N__18048),
            .I(N__18042));
    CascadeBuf I__3852 (
            .O(N__18045),
            .I(N__18039));
    CascadeBuf I__3851 (
            .O(N__18042),
            .I(N__18036));
    CascadeMux I__3850 (
            .O(N__18039),
            .I(N__18033));
    CascadeMux I__3849 (
            .O(N__18036),
            .I(N__18030));
    CascadeBuf I__3848 (
            .O(N__18033),
            .I(N__18027));
    CascadeBuf I__3847 (
            .O(N__18030),
            .I(N__18024));
    CascadeMux I__3846 (
            .O(N__18027),
            .I(N__18021));
    CascadeMux I__3845 (
            .O(N__18024),
            .I(N__18018));
    CascadeBuf I__3844 (
            .O(N__18021),
            .I(N__18015));
    CascadeBuf I__3843 (
            .O(N__18018),
            .I(N__18012));
    CascadeMux I__3842 (
            .O(N__18015),
            .I(N__18009));
    CascadeMux I__3841 (
            .O(N__18012),
            .I(N__18006));
    InMux I__3840 (
            .O(N__18009),
            .I(N__18003));
    InMux I__3839 (
            .O(N__18006),
            .I(N__18000));
    LocalMux I__3838 (
            .O(N__18003),
            .I(N__17997));
    LocalMux I__3837 (
            .O(N__18000),
            .I(N__17994));
    Span12Mux_s11_h I__3836 (
            .O(N__17997),
            .I(N__17991));
    Sp12to4 I__3835 (
            .O(N__17994),
            .I(N__17988));
    Span12Mux_v I__3834 (
            .O(N__17991),
            .I(N__17983));
    Span12Mux_v I__3833 (
            .O(N__17988),
            .I(N__17983));
    Odrv12 I__3832 (
            .O(N__17983),
            .I(n25));
    InMux I__3831 (
            .O(N__17980),
            .I(N__17976));
    InMux I__3830 (
            .O(N__17979),
            .I(N__17973));
    LocalMux I__3829 (
            .O(N__17976),
            .I(N__17969));
    LocalMux I__3828 (
            .O(N__17973),
            .I(N__17966));
    InMux I__3827 (
            .O(N__17972),
            .I(N__17963));
    Span4Mux_v I__3826 (
            .O(N__17969),
            .I(N__17956));
    Span4Mux_h I__3825 (
            .O(N__17966),
            .I(N__17956));
    LocalMux I__3824 (
            .O(N__17963),
            .I(N__17956));
    Span4Mux_v I__3823 (
            .O(N__17956),
            .I(N__17952));
    InMux I__3822 (
            .O(N__17955),
            .I(N__17949));
    Odrv4 I__3821 (
            .O(N__17952),
            .I(\transmit_module.TX_ADDR_2 ));
    LocalMux I__3820 (
            .O(N__17949),
            .I(\transmit_module.TX_ADDR_2 ));
    InMux I__3819 (
            .O(N__17944),
            .I(N__17941));
    LocalMux I__3818 (
            .O(N__17941),
            .I(\transmit_module.ADDR_Y_COMPONENT_2 ));
    InMux I__3817 (
            .O(N__17938),
            .I(N__17934));
    InMux I__3816 (
            .O(N__17937),
            .I(N__17930));
    LocalMux I__3815 (
            .O(N__17934),
            .I(N__17924));
    InMux I__3814 (
            .O(N__17933),
            .I(N__17921));
    LocalMux I__3813 (
            .O(N__17930),
            .I(N__17918));
    InMux I__3812 (
            .O(N__17929),
            .I(N__17915));
    InMux I__3811 (
            .O(N__17928),
            .I(N__17912));
    InMux I__3810 (
            .O(N__17927),
            .I(N__17909));
    Span4Mux_h I__3809 (
            .O(N__17924),
            .I(N__17900));
    LocalMux I__3808 (
            .O(N__17921),
            .I(N__17900));
    Span4Mux_v I__3807 (
            .O(N__17918),
            .I(N__17897));
    LocalMux I__3806 (
            .O(N__17915),
            .I(N__17894));
    LocalMux I__3805 (
            .O(N__17912),
            .I(N__17891));
    LocalMux I__3804 (
            .O(N__17909),
            .I(N__17888));
    InMux I__3803 (
            .O(N__17908),
            .I(N__17885));
    InMux I__3802 (
            .O(N__17907),
            .I(N__17878));
    InMux I__3801 (
            .O(N__17906),
            .I(N__17875));
    InMux I__3800 (
            .O(N__17905),
            .I(N__17872));
    Span4Mux_v I__3799 (
            .O(N__17900),
            .I(N__17863));
    Span4Mux_h I__3798 (
            .O(N__17897),
            .I(N__17863));
    Span4Mux_v I__3797 (
            .O(N__17894),
            .I(N__17863));
    Span4Mux_v I__3796 (
            .O(N__17891),
            .I(N__17863));
    Sp12to4 I__3795 (
            .O(N__17888),
            .I(N__17858));
    LocalMux I__3794 (
            .O(N__17885),
            .I(N__17858));
    InMux I__3793 (
            .O(N__17884),
            .I(N__17855));
    InMux I__3792 (
            .O(N__17883),
            .I(N__17852));
    InMux I__3791 (
            .O(N__17882),
            .I(N__17849));
    InMux I__3790 (
            .O(N__17881),
            .I(N__17846));
    LocalMux I__3789 (
            .O(N__17878),
            .I(\transmit_module.Y_DELTA_PATTERN_0 ));
    LocalMux I__3788 (
            .O(N__17875),
            .I(\transmit_module.Y_DELTA_PATTERN_0 ));
    LocalMux I__3787 (
            .O(N__17872),
            .I(\transmit_module.Y_DELTA_PATTERN_0 ));
    Odrv4 I__3786 (
            .O(N__17863),
            .I(\transmit_module.Y_DELTA_PATTERN_0 ));
    Odrv12 I__3785 (
            .O(N__17858),
            .I(\transmit_module.Y_DELTA_PATTERN_0 ));
    LocalMux I__3784 (
            .O(N__17855),
            .I(\transmit_module.Y_DELTA_PATTERN_0 ));
    LocalMux I__3783 (
            .O(N__17852),
            .I(\transmit_module.Y_DELTA_PATTERN_0 ));
    LocalMux I__3782 (
            .O(N__17849),
            .I(\transmit_module.Y_DELTA_PATTERN_0 ));
    LocalMux I__3781 (
            .O(N__17846),
            .I(\transmit_module.Y_DELTA_PATTERN_0 ));
    InMux I__3780 (
            .O(N__17827),
            .I(N__17824));
    LocalMux I__3779 (
            .O(N__17824),
            .I(N__17821));
    Span4Mux_v I__3778 (
            .O(N__17821),
            .I(N__17817));
    InMux I__3777 (
            .O(N__17820),
            .I(N__17814));
    Odrv4 I__3776 (
            .O(N__17817),
            .I(\transmit_module.n113 ));
    LocalMux I__3775 (
            .O(N__17814),
            .I(\transmit_module.n113 ));
    InMux I__3774 (
            .O(N__17809),
            .I(N__17800));
    InMux I__3773 (
            .O(N__17808),
            .I(N__17800));
    InMux I__3772 (
            .O(N__17807),
            .I(N__17800));
    LocalMux I__3771 (
            .O(N__17800),
            .I(N__17797));
    Span4Mux_v I__3770 (
            .O(N__17797),
            .I(N__17793));
    InMux I__3769 (
            .O(N__17796),
            .I(N__17790));
    Odrv4 I__3768 (
            .O(N__17793),
            .I(\transmit_module.TX_ADDR_3 ));
    LocalMux I__3767 (
            .O(N__17790),
            .I(\transmit_module.TX_ADDR_3 ));
    InMux I__3766 (
            .O(N__17785),
            .I(N__17782));
    LocalMux I__3765 (
            .O(N__17782),
            .I(\transmit_module.ADDR_Y_COMPONENT_3 ));
    CEMux I__3764 (
            .O(N__17779),
            .I(N__17775));
    CEMux I__3763 (
            .O(N__17778),
            .I(N__17771));
    LocalMux I__3762 (
            .O(N__17775),
            .I(N__17767));
    CEMux I__3761 (
            .O(N__17774),
            .I(N__17763));
    LocalMux I__3760 (
            .O(N__17771),
            .I(N__17759));
    CEMux I__3759 (
            .O(N__17770),
            .I(N__17756));
    Span4Mux_v I__3758 (
            .O(N__17767),
            .I(N__17753));
    CEMux I__3757 (
            .O(N__17766),
            .I(N__17750));
    LocalMux I__3756 (
            .O(N__17763),
            .I(N__17747));
    CEMux I__3755 (
            .O(N__17762),
            .I(N__17744));
    Span4Mux_v I__3754 (
            .O(N__17759),
            .I(N__17738));
    LocalMux I__3753 (
            .O(N__17756),
            .I(N__17738));
    Span4Mux_h I__3752 (
            .O(N__17753),
            .I(N__17733));
    LocalMux I__3751 (
            .O(N__17750),
            .I(N__17733));
    Span4Mux_v I__3750 (
            .O(N__17747),
            .I(N__17728));
    LocalMux I__3749 (
            .O(N__17744),
            .I(N__17728));
    CEMux I__3748 (
            .O(N__17743),
            .I(N__17725));
    Span4Mux_h I__3747 (
            .O(N__17738),
            .I(N__17720));
    Span4Mux_h I__3746 (
            .O(N__17733),
            .I(N__17720));
    Span4Mux_v I__3745 (
            .O(N__17728),
            .I(N__17717));
    LocalMux I__3744 (
            .O(N__17725),
            .I(N__17714));
    Odrv4 I__3743 (
            .O(N__17720),
            .I(\transmit_module.n2061 ));
    Odrv4 I__3742 (
            .O(N__17717),
            .I(\transmit_module.n2061 ));
    Odrv4 I__3741 (
            .O(N__17714),
            .I(\transmit_module.n2061 ));
    InMux I__3740 (
            .O(N__17707),
            .I(N__17704));
    LocalMux I__3739 (
            .O(N__17704),
            .I(N__17701));
    Odrv4 I__3738 (
            .O(N__17701),
            .I(TX_DATA_4));
    IoInMux I__3737 (
            .O(N__17698),
            .I(N__17694));
    IoInMux I__3736 (
            .O(N__17697),
            .I(N__17690));
    LocalMux I__3735 (
            .O(N__17694),
            .I(N__17687));
    IoInMux I__3734 (
            .O(N__17693),
            .I(N__17684));
    LocalMux I__3733 (
            .O(N__17690),
            .I(N__17681));
    IoSpan4Mux I__3732 (
            .O(N__17687),
            .I(N__17678));
    LocalMux I__3731 (
            .O(N__17684),
            .I(N__17675));
    IoSpan4Mux I__3730 (
            .O(N__17681),
            .I(N__17672));
    Span4Mux_s3_h I__3729 (
            .O(N__17678),
            .I(N__17669));
    Span4Mux_s2_v I__3728 (
            .O(N__17675),
            .I(N__17666));
    Span4Mux_s2_v I__3727 (
            .O(N__17672),
            .I(N__17663));
    Span4Mux_h I__3726 (
            .O(N__17669),
            .I(N__17660));
    Sp12to4 I__3725 (
            .O(N__17666),
            .I(N__17657));
    Sp12to4 I__3724 (
            .O(N__17663),
            .I(N__17654));
    Span4Mux_h I__3723 (
            .O(N__17660),
            .I(N__17651));
    Span12Mux_h I__3722 (
            .O(N__17657),
            .I(N__17646));
    Span12Mux_h I__3721 (
            .O(N__17654),
            .I(N__17646));
    Span4Mux_h I__3720 (
            .O(N__17651),
            .I(N__17643));
    Odrv12 I__3719 (
            .O(N__17646),
            .I(n1794));
    Odrv4 I__3718 (
            .O(N__17643),
            .I(n1794));
    InMux I__3717 (
            .O(N__17638),
            .I(N__17635));
    LocalMux I__3716 (
            .O(N__17635),
            .I(N__17632));
    Odrv4 I__3715 (
            .O(N__17632),
            .I(TX_DATA_2));
    IoInMux I__3714 (
            .O(N__17629),
            .I(N__17625));
    IoInMux I__3713 (
            .O(N__17628),
            .I(N__17621));
    LocalMux I__3712 (
            .O(N__17625),
            .I(N__17618));
    IoInMux I__3711 (
            .O(N__17624),
            .I(N__17615));
    LocalMux I__3710 (
            .O(N__17621),
            .I(N__17612));
    Span4Mux_s3_h I__3709 (
            .O(N__17618),
            .I(N__17609));
    LocalMux I__3708 (
            .O(N__17615),
            .I(N__17606));
    Span12Mux_s5_v I__3707 (
            .O(N__17612),
            .I(N__17601));
    Sp12to4 I__3706 (
            .O(N__17609),
            .I(N__17601));
    IoSpan4Mux I__3705 (
            .O(N__17606),
            .I(N__17598));
    Span12Mux_v I__3704 (
            .O(N__17601),
            .I(N__17595));
    Sp12to4 I__3703 (
            .O(N__17598),
            .I(N__17592));
    Span12Mux_h I__3702 (
            .O(N__17595),
            .I(N__17589));
    Span12Mux_v I__3701 (
            .O(N__17592),
            .I(N__17586));
    Odrv12 I__3700 (
            .O(N__17589),
            .I(n1796));
    Odrv12 I__3699 (
            .O(N__17586),
            .I(n1796));
    InMux I__3698 (
            .O(N__17581),
            .I(N__17578));
    LocalMux I__3697 (
            .O(N__17578),
            .I(\transmit_module.ADDR_Y_COMPONENT_13 ));
    InMux I__3696 (
            .O(N__17575),
            .I(N__17572));
    LocalMux I__3695 (
            .O(N__17572),
            .I(N__17569));
    Span12Mux_v I__3694 (
            .O(N__17569),
            .I(N__17566));
    Odrv12 I__3693 (
            .O(N__17566),
            .I(\line_buffer.n3634 ));
    InMux I__3692 (
            .O(N__17563),
            .I(N__17560));
    LocalMux I__3691 (
            .O(N__17560),
            .I(N__17557));
    Span4Mux_v I__3690 (
            .O(N__17557),
            .I(N__17554));
    Span4Mux_h I__3689 (
            .O(N__17554),
            .I(N__17551));
    Span4Mux_h I__3688 (
            .O(N__17551),
            .I(N__17548));
    Odrv4 I__3687 (
            .O(N__17548),
            .I(\line_buffer.n442 ));
    CascadeMux I__3686 (
            .O(N__17545),
            .I(N__17542));
    InMux I__3685 (
            .O(N__17542),
            .I(N__17539));
    LocalMux I__3684 (
            .O(N__17539),
            .I(N__17536));
    Span4Mux_v I__3683 (
            .O(N__17536),
            .I(N__17533));
    Span4Mux_h I__3682 (
            .O(N__17533),
            .I(N__17530));
    Span4Mux_h I__3681 (
            .O(N__17530),
            .I(N__17527));
    Span4Mux_v I__3680 (
            .O(N__17527),
            .I(N__17524));
    Odrv4 I__3679 (
            .O(N__17524),
            .I(\line_buffer.n434 ));
    InMux I__3678 (
            .O(N__17521),
            .I(N__17518));
    LocalMux I__3677 (
            .O(N__17518),
            .I(\line_buffer.n3749 ));
    InMux I__3676 (
            .O(N__17515),
            .I(N__17512));
    LocalMux I__3675 (
            .O(N__17512),
            .I(N__17509));
    Span4Mux_v I__3674 (
            .O(N__17509),
            .I(N__17506));
    Span4Mux_h I__3673 (
            .O(N__17506),
            .I(N__17503));
    Span4Mux_h I__3672 (
            .O(N__17503),
            .I(N__17500));
    Odrv4 I__3671 (
            .O(N__17500),
            .I(\line_buffer.n541 ));
    InMux I__3670 (
            .O(N__17497),
            .I(N__17494));
    LocalMux I__3669 (
            .O(N__17494),
            .I(N__17491));
    Span4Mux_v I__3668 (
            .O(N__17491),
            .I(N__17488));
    Span4Mux_h I__3667 (
            .O(N__17488),
            .I(N__17485));
    Span4Mux_h I__3666 (
            .O(N__17485),
            .I(N__17482));
    Odrv4 I__3665 (
            .O(N__17482),
            .I(\line_buffer.n533 ));
    InMux I__3664 (
            .O(N__17479),
            .I(N__17476));
    LocalMux I__3663 (
            .O(N__17476),
            .I(N__17473));
    Span12Mux_v I__3662 (
            .O(N__17473),
            .I(N__17470));
    Odrv12 I__3661 (
            .O(N__17470),
            .I(\line_buffer.n3676 ));
    InMux I__3660 (
            .O(N__17467),
            .I(N__17464));
    LocalMux I__3659 (
            .O(N__17464),
            .I(\line_buffer.n3674 ));
    InMux I__3658 (
            .O(N__17461),
            .I(N__17458));
    LocalMux I__3657 (
            .O(N__17458),
            .I(\line_buffer.n3716 ));
    InMux I__3656 (
            .O(N__17455),
            .I(N__17452));
    LocalMux I__3655 (
            .O(N__17452),
            .I(N__17449));
    Span4Mux_v I__3654 (
            .O(N__17449),
            .I(N__17446));
    Sp12to4 I__3653 (
            .O(N__17446),
            .I(N__17443));
    Odrv12 I__3652 (
            .O(N__17443),
            .I(\line_buffer.n446 ));
    InMux I__3651 (
            .O(N__17440),
            .I(N__17437));
    LocalMux I__3650 (
            .O(N__17437),
            .I(N__17434));
    Span12Mux_h I__3649 (
            .O(N__17434),
            .I(N__17431));
    Span12Mux_v I__3648 (
            .O(N__17431),
            .I(N__17428));
    Odrv12 I__3647 (
            .O(N__17428),
            .I(\line_buffer.n438 ));
    InMux I__3646 (
            .O(N__17425),
            .I(N__17422));
    LocalMux I__3645 (
            .O(N__17422),
            .I(\line_buffer.n3728 ));
    CascadeMux I__3644 (
            .O(N__17419),
            .I(\line_buffer.n3640_cascade_ ));
    InMux I__3643 (
            .O(N__17416),
            .I(N__17413));
    LocalMux I__3642 (
            .O(N__17413),
            .I(N__17410));
    Span4Mux_v I__3641 (
            .O(N__17410),
            .I(N__17407));
    Span4Mux_v I__3640 (
            .O(N__17407),
            .I(N__17404));
    Odrv4 I__3639 (
            .O(N__17404),
            .I(\line_buffer.n3641 ));
    InMux I__3638 (
            .O(N__17401),
            .I(N__17398));
    LocalMux I__3637 (
            .O(N__17398),
            .I(N__17395));
    Odrv12 I__3636 (
            .O(N__17395),
            .I(RX_TX_SYNC_BUFF));
    InMux I__3635 (
            .O(N__17392),
            .I(N__17389));
    LocalMux I__3634 (
            .O(N__17389),
            .I(N__17386));
    Span4Mux_v I__3633 (
            .O(N__17386),
            .I(N__17383));
    Odrv4 I__3632 (
            .O(N__17383),
            .I(RX_TX_SYNC));
    InMux I__3631 (
            .O(N__17380),
            .I(N__17377));
    LocalMux I__3630 (
            .O(N__17377),
            .I(\sync_buffer.BUFFER_0 ));
    InMux I__3629 (
            .O(N__17374),
            .I(N__17371));
    LocalMux I__3628 (
            .O(N__17371),
            .I(\sync_buffer.BUFFER_1 ));
    InMux I__3627 (
            .O(N__17368),
            .I(N__17365));
    LocalMux I__3626 (
            .O(N__17365),
            .I(\transmit_module.n124 ));
    CascadeMux I__3625 (
            .O(N__17362),
            .I(\transmit_module.n139_cascade_ ));
    InMux I__3624 (
            .O(N__17359),
            .I(N__17356));
    LocalMux I__3623 (
            .O(N__17356),
            .I(\transmit_module.ADDR_Y_COMPONENT_8 ));
    CascadeMux I__3622 (
            .O(N__17353),
            .I(N__17347));
    InMux I__3621 (
            .O(N__17352),
            .I(N__17342));
    InMux I__3620 (
            .O(N__17351),
            .I(N__17342));
    InMux I__3619 (
            .O(N__17350),
            .I(N__17337));
    InMux I__3618 (
            .O(N__17347),
            .I(N__17337));
    LocalMux I__3617 (
            .O(N__17342),
            .I(\transmit_module.TX_ADDR_8 ));
    LocalMux I__3616 (
            .O(N__17337),
            .I(\transmit_module.TX_ADDR_8 ));
    CascadeMux I__3615 (
            .O(N__17332),
            .I(N__17326));
    InMux I__3614 (
            .O(N__17331),
            .I(N__17323));
    InMux I__3613 (
            .O(N__17330),
            .I(N__17320));
    InMux I__3612 (
            .O(N__17329),
            .I(N__17315));
    InMux I__3611 (
            .O(N__17326),
            .I(N__17315));
    LocalMux I__3610 (
            .O(N__17323),
            .I(\transmit_module.TX_ADDR_9 ));
    LocalMux I__3609 (
            .O(N__17320),
            .I(\transmit_module.TX_ADDR_9 ));
    LocalMux I__3608 (
            .O(N__17315),
            .I(\transmit_module.TX_ADDR_9 ));
    InMux I__3607 (
            .O(N__17308),
            .I(N__17305));
    LocalMux I__3606 (
            .O(N__17305),
            .I(\transmit_module.n123 ));
    InMux I__3605 (
            .O(N__17302),
            .I(N__17299));
    LocalMux I__3604 (
            .O(N__17299),
            .I(\transmit_module.n138 ));
    CascadeMux I__3603 (
            .O(N__17296),
            .I(\transmit_module.n138_cascade_ ));
    InMux I__3602 (
            .O(N__17293),
            .I(N__17287));
    InMux I__3601 (
            .O(N__17292),
            .I(N__17287));
    LocalMux I__3600 (
            .O(N__17287),
            .I(\transmit_module.n107 ));
    CascadeMux I__3599 (
            .O(N__17284),
            .I(N__17280));
    CascadeMux I__3598 (
            .O(N__17283),
            .I(N__17277));
    CascadeBuf I__3597 (
            .O(N__17280),
            .I(N__17274));
    CascadeBuf I__3596 (
            .O(N__17277),
            .I(N__17271));
    CascadeMux I__3595 (
            .O(N__17274),
            .I(N__17268));
    CascadeMux I__3594 (
            .O(N__17271),
            .I(N__17265));
    CascadeBuf I__3593 (
            .O(N__17268),
            .I(N__17262));
    CascadeBuf I__3592 (
            .O(N__17265),
            .I(N__17259));
    CascadeMux I__3591 (
            .O(N__17262),
            .I(N__17256));
    CascadeMux I__3590 (
            .O(N__17259),
            .I(N__17253));
    CascadeBuf I__3589 (
            .O(N__17256),
            .I(N__17250));
    CascadeBuf I__3588 (
            .O(N__17253),
            .I(N__17247));
    CascadeMux I__3587 (
            .O(N__17250),
            .I(N__17244));
    CascadeMux I__3586 (
            .O(N__17247),
            .I(N__17241));
    CascadeBuf I__3585 (
            .O(N__17244),
            .I(N__17238));
    CascadeBuf I__3584 (
            .O(N__17241),
            .I(N__17235));
    CascadeMux I__3583 (
            .O(N__17238),
            .I(N__17232));
    CascadeMux I__3582 (
            .O(N__17235),
            .I(N__17229));
    CascadeBuf I__3581 (
            .O(N__17232),
            .I(N__17226));
    CascadeBuf I__3580 (
            .O(N__17229),
            .I(N__17223));
    CascadeMux I__3579 (
            .O(N__17226),
            .I(N__17220));
    CascadeMux I__3578 (
            .O(N__17223),
            .I(N__17217));
    CascadeBuf I__3577 (
            .O(N__17220),
            .I(N__17214));
    CascadeBuf I__3576 (
            .O(N__17217),
            .I(N__17211));
    CascadeMux I__3575 (
            .O(N__17214),
            .I(N__17208));
    CascadeMux I__3574 (
            .O(N__17211),
            .I(N__17205));
    CascadeBuf I__3573 (
            .O(N__17208),
            .I(N__17202));
    CascadeBuf I__3572 (
            .O(N__17205),
            .I(N__17199));
    CascadeMux I__3571 (
            .O(N__17202),
            .I(N__17196));
    CascadeMux I__3570 (
            .O(N__17199),
            .I(N__17193));
    CascadeBuf I__3569 (
            .O(N__17196),
            .I(N__17190));
    CascadeBuf I__3568 (
            .O(N__17193),
            .I(N__17187));
    CascadeMux I__3567 (
            .O(N__17190),
            .I(N__17184));
    CascadeMux I__3566 (
            .O(N__17187),
            .I(N__17181));
    CascadeBuf I__3565 (
            .O(N__17184),
            .I(N__17178));
    CascadeBuf I__3564 (
            .O(N__17181),
            .I(N__17175));
    CascadeMux I__3563 (
            .O(N__17178),
            .I(N__17172));
    CascadeMux I__3562 (
            .O(N__17175),
            .I(N__17169));
    CascadeBuf I__3561 (
            .O(N__17172),
            .I(N__17166));
    CascadeBuf I__3560 (
            .O(N__17169),
            .I(N__17163));
    CascadeMux I__3559 (
            .O(N__17166),
            .I(N__17160));
    CascadeMux I__3558 (
            .O(N__17163),
            .I(N__17157));
    CascadeBuf I__3557 (
            .O(N__17160),
            .I(N__17154));
    CascadeBuf I__3556 (
            .O(N__17157),
            .I(N__17151));
    CascadeMux I__3555 (
            .O(N__17154),
            .I(N__17148));
    CascadeMux I__3554 (
            .O(N__17151),
            .I(N__17145));
    CascadeBuf I__3553 (
            .O(N__17148),
            .I(N__17142));
    CascadeBuf I__3552 (
            .O(N__17145),
            .I(N__17139));
    CascadeMux I__3551 (
            .O(N__17142),
            .I(N__17136));
    CascadeMux I__3550 (
            .O(N__17139),
            .I(N__17133));
    CascadeBuf I__3549 (
            .O(N__17136),
            .I(N__17130));
    CascadeBuf I__3548 (
            .O(N__17133),
            .I(N__17127));
    CascadeMux I__3547 (
            .O(N__17130),
            .I(N__17124));
    CascadeMux I__3546 (
            .O(N__17127),
            .I(N__17121));
    CascadeBuf I__3545 (
            .O(N__17124),
            .I(N__17118));
    CascadeBuf I__3544 (
            .O(N__17121),
            .I(N__17115));
    CascadeMux I__3543 (
            .O(N__17118),
            .I(N__17112));
    CascadeMux I__3542 (
            .O(N__17115),
            .I(N__17109));
    CascadeBuf I__3541 (
            .O(N__17112),
            .I(N__17106));
    CascadeBuf I__3540 (
            .O(N__17109),
            .I(N__17103));
    CascadeMux I__3539 (
            .O(N__17106),
            .I(N__17100));
    CascadeMux I__3538 (
            .O(N__17103),
            .I(N__17097));
    InMux I__3537 (
            .O(N__17100),
            .I(N__17094));
    InMux I__3536 (
            .O(N__17097),
            .I(N__17091));
    LocalMux I__3535 (
            .O(N__17094),
            .I(N__17088));
    LocalMux I__3534 (
            .O(N__17091),
            .I(N__17085));
    Span4Mux_v I__3533 (
            .O(N__17088),
            .I(N__17082));
    Span4Mux_v I__3532 (
            .O(N__17085),
            .I(N__17079));
    Span4Mux_v I__3531 (
            .O(N__17082),
            .I(N__17076));
    Span4Mux_v I__3530 (
            .O(N__17079),
            .I(N__17073));
    Span4Mux_v I__3529 (
            .O(N__17076),
            .I(N__17070));
    Sp12to4 I__3528 (
            .O(N__17073),
            .I(N__17067));
    Span4Mux_v I__3527 (
            .O(N__17070),
            .I(N__17064));
    Span12Mux_v I__3526 (
            .O(N__17067),
            .I(N__17061));
    Span4Mux_h I__3525 (
            .O(N__17064),
            .I(N__17058));
    Odrv12 I__3524 (
            .O(N__17061),
            .I(n19));
    Odrv4 I__3523 (
            .O(N__17058),
            .I(n19));
    CEMux I__3522 (
            .O(N__17053),
            .I(N__17050));
    LocalMux I__3521 (
            .O(N__17050),
            .I(N__17047));
    Span4Mux_v I__3520 (
            .O(N__17047),
            .I(N__17044));
    Odrv4 I__3519 (
            .O(N__17044),
            .I(\receive_module.n3795 ));
    SRMux I__3518 (
            .O(N__17041),
            .I(N__17037));
    SRMux I__3517 (
            .O(N__17040),
            .I(N__17034));
    LocalMux I__3516 (
            .O(N__17037),
            .I(N__17028));
    LocalMux I__3515 (
            .O(N__17034),
            .I(N__17028));
    SRMux I__3514 (
            .O(N__17033),
            .I(N__17025));
    Span4Mux_v I__3513 (
            .O(N__17028),
            .I(N__17019));
    LocalMux I__3512 (
            .O(N__17025),
            .I(N__17019));
    SRMux I__3511 (
            .O(N__17024),
            .I(N__17016));
    Span4Mux_h I__3510 (
            .O(N__17019),
            .I(N__17013));
    LocalMux I__3509 (
            .O(N__17016),
            .I(N__17010));
    Span4Mux_h I__3508 (
            .O(N__17013),
            .I(N__17007));
    Span4Mux_v I__3507 (
            .O(N__17010),
            .I(N__17004));
    Sp12to4 I__3506 (
            .O(N__17007),
            .I(N__17001));
    Span4Mux_h I__3505 (
            .O(N__17004),
            .I(N__16998));
    Span12Mux_s10_v I__3504 (
            .O(N__17001),
            .I(N__16995));
    Span4Mux_h I__3503 (
            .O(N__16998),
            .I(N__16992));
    Odrv12 I__3502 (
            .O(N__16995),
            .I(\line_buffer.n451 ));
    Odrv4 I__3501 (
            .O(N__16992),
            .I(\line_buffer.n451 ));
    SRMux I__3500 (
            .O(N__16987),
            .I(N__16983));
    SRMux I__3499 (
            .O(N__16986),
            .I(N__16980));
    LocalMux I__3498 (
            .O(N__16983),
            .I(N__16977));
    LocalMux I__3497 (
            .O(N__16980),
            .I(N__16973));
    Span4Mux_v I__3496 (
            .O(N__16977),
            .I(N__16969));
    SRMux I__3495 (
            .O(N__16976),
            .I(N__16966));
    Span4Mux_h I__3494 (
            .O(N__16973),
            .I(N__16963));
    SRMux I__3493 (
            .O(N__16972),
            .I(N__16960));
    Sp12to4 I__3492 (
            .O(N__16969),
            .I(N__16957));
    LocalMux I__3491 (
            .O(N__16966),
            .I(N__16954));
    Span4Mux_v I__3490 (
            .O(N__16963),
            .I(N__16949));
    LocalMux I__3489 (
            .O(N__16960),
            .I(N__16949));
    Span12Mux_v I__3488 (
            .O(N__16957),
            .I(N__16942));
    Span12Mux_s11_v I__3487 (
            .O(N__16954),
            .I(N__16942));
    Sp12to4 I__3486 (
            .O(N__16949),
            .I(N__16942));
    Odrv12 I__3485 (
            .O(N__16942),
            .I(\line_buffer.n549 ));
    SRMux I__3484 (
            .O(N__16939),
            .I(N__16936));
    LocalMux I__3483 (
            .O(N__16936),
            .I(N__16932));
    SRMux I__3482 (
            .O(N__16935),
            .I(N__16929));
    Span4Mux_s3_v I__3481 (
            .O(N__16932),
            .I(N__16925));
    LocalMux I__3480 (
            .O(N__16929),
            .I(N__16922));
    SRMux I__3479 (
            .O(N__16928),
            .I(N__16919));
    Span4Mux_v I__3478 (
            .O(N__16925),
            .I(N__16912));
    Span4Mux_h I__3477 (
            .O(N__16922),
            .I(N__16912));
    LocalMux I__3476 (
            .O(N__16919),
            .I(N__16912));
    Span4Mux_v I__3475 (
            .O(N__16912),
            .I(N__16909));
    Span4Mux_h I__3474 (
            .O(N__16909),
            .I(N__16905));
    SRMux I__3473 (
            .O(N__16908),
            .I(N__16902));
    Sp12to4 I__3472 (
            .O(N__16905),
            .I(N__16897));
    LocalMux I__3471 (
            .O(N__16902),
            .I(N__16897));
    Span12Mux_h I__3470 (
            .O(N__16897),
            .I(N__16894));
    Odrv12 I__3469 (
            .O(N__16894),
            .I(\line_buffer.n516 ));
    InMux I__3468 (
            .O(N__16891),
            .I(N__16888));
    LocalMux I__3467 (
            .O(N__16888),
            .I(N__16885));
    Span4Mux_h I__3466 (
            .O(N__16885),
            .I(N__16882));
    Odrv4 I__3465 (
            .O(N__16882),
            .I(\receive_module.rx_counter.n3575 ));
    InMux I__3464 (
            .O(N__16879),
            .I(N__16876));
    LocalMux I__3463 (
            .O(N__16876),
            .I(N__16873));
    Odrv4 I__3462 (
            .O(N__16873),
            .I(\receive_module.rx_counter.n4_adj_606 ));
    CascadeMux I__3461 (
            .O(N__16870),
            .I(N__16867));
    InMux I__3460 (
            .O(N__16867),
            .I(N__16864));
    LocalMux I__3459 (
            .O(N__16864),
            .I(N__16859));
    CascadeMux I__3458 (
            .O(N__16863),
            .I(N__16855));
    InMux I__3457 (
            .O(N__16862),
            .I(N__16852));
    Span4Mux_h I__3456 (
            .O(N__16859),
            .I(N__16849));
    InMux I__3455 (
            .O(N__16858),
            .I(N__16846));
    InMux I__3454 (
            .O(N__16855),
            .I(N__16843));
    LocalMux I__3453 (
            .O(N__16852),
            .I(\receive_module.rx_counter.Y_8 ));
    Odrv4 I__3452 (
            .O(N__16849),
            .I(\receive_module.rx_counter.Y_8 ));
    LocalMux I__3451 (
            .O(N__16846),
            .I(\receive_module.rx_counter.Y_8 ));
    LocalMux I__3450 (
            .O(N__16843),
            .I(\receive_module.rx_counter.Y_8 ));
    InMux I__3449 (
            .O(N__16834),
            .I(N__16831));
    LocalMux I__3448 (
            .O(N__16831),
            .I(\receive_module.rx_counter.n55_adj_607 ));
    SRMux I__3447 (
            .O(N__16828),
            .I(N__16825));
    LocalMux I__3446 (
            .O(N__16825),
            .I(N__16821));
    SRMux I__3445 (
            .O(N__16824),
            .I(N__16818));
    Span4Mux_v I__3444 (
            .O(N__16821),
            .I(N__16812));
    LocalMux I__3443 (
            .O(N__16818),
            .I(N__16812));
    SRMux I__3442 (
            .O(N__16817),
            .I(N__16809));
    Span4Mux_v I__3441 (
            .O(N__16812),
            .I(N__16803));
    LocalMux I__3440 (
            .O(N__16809),
            .I(N__16803));
    SRMux I__3439 (
            .O(N__16808),
            .I(N__16800));
    Span4Mux_v I__3438 (
            .O(N__16803),
            .I(N__16795));
    LocalMux I__3437 (
            .O(N__16800),
            .I(N__16795));
    Span4Mux_h I__3436 (
            .O(N__16795),
            .I(N__16792));
    Span4Mux_h I__3435 (
            .O(N__16792),
            .I(N__16789));
    Odrv4 I__3434 (
            .O(N__16789),
            .I(\line_buffer.n581 ));
    CascadeMux I__3433 (
            .O(N__16786),
            .I(N__16776));
    CascadeMux I__3432 (
            .O(N__16785),
            .I(N__16773));
    InMux I__3431 (
            .O(N__16784),
            .I(N__16769));
    InMux I__3430 (
            .O(N__16783),
            .I(N__16762));
    InMux I__3429 (
            .O(N__16782),
            .I(N__16762));
    InMux I__3428 (
            .O(N__16781),
            .I(N__16762));
    InMux I__3427 (
            .O(N__16780),
            .I(N__16757));
    InMux I__3426 (
            .O(N__16779),
            .I(N__16757));
    InMux I__3425 (
            .O(N__16776),
            .I(N__16750));
    InMux I__3424 (
            .O(N__16773),
            .I(N__16750));
    InMux I__3423 (
            .O(N__16772),
            .I(N__16750));
    LocalMux I__3422 (
            .O(N__16769),
            .I(RX_ADDR_12));
    LocalMux I__3421 (
            .O(N__16762),
            .I(RX_ADDR_12));
    LocalMux I__3420 (
            .O(N__16757),
            .I(RX_ADDR_12));
    LocalMux I__3419 (
            .O(N__16750),
            .I(RX_ADDR_12));
    CascadeMux I__3418 (
            .O(N__16741),
            .I(N__16732));
    CascadeMux I__3417 (
            .O(N__16740),
            .I(N__16729));
    CascadeMux I__3416 (
            .O(N__16739),
            .I(N__16726));
    CascadeMux I__3415 (
            .O(N__16738),
            .I(N__16721));
    InMux I__3414 (
            .O(N__16737),
            .I(N__16718));
    InMux I__3413 (
            .O(N__16736),
            .I(N__16711));
    InMux I__3412 (
            .O(N__16735),
            .I(N__16711));
    InMux I__3411 (
            .O(N__16732),
            .I(N__16711));
    InMux I__3410 (
            .O(N__16729),
            .I(N__16708));
    InMux I__3409 (
            .O(N__16726),
            .I(N__16705));
    InMux I__3408 (
            .O(N__16725),
            .I(N__16698));
    InMux I__3407 (
            .O(N__16724),
            .I(N__16698));
    InMux I__3406 (
            .O(N__16721),
            .I(N__16698));
    LocalMux I__3405 (
            .O(N__16718),
            .I(RX_ADDR_13));
    LocalMux I__3404 (
            .O(N__16711),
            .I(RX_ADDR_13));
    LocalMux I__3403 (
            .O(N__16708),
            .I(RX_ADDR_13));
    LocalMux I__3402 (
            .O(N__16705),
            .I(RX_ADDR_13));
    LocalMux I__3401 (
            .O(N__16698),
            .I(RX_ADDR_13));
    CascadeMux I__3400 (
            .O(N__16687),
            .I(N__16682));
    CascadeMux I__3399 (
            .O(N__16686),
            .I(N__16679));
    InMux I__3398 (
            .O(N__16685),
            .I(N__16670));
    InMux I__3397 (
            .O(N__16682),
            .I(N__16665));
    InMux I__3396 (
            .O(N__16679),
            .I(N__16665));
    InMux I__3395 (
            .O(N__16678),
            .I(N__16662));
    InMux I__3394 (
            .O(N__16677),
            .I(N__16657));
    InMux I__3393 (
            .O(N__16676),
            .I(N__16657));
    InMux I__3392 (
            .O(N__16675),
            .I(N__16650));
    InMux I__3391 (
            .O(N__16674),
            .I(N__16650));
    InMux I__3390 (
            .O(N__16673),
            .I(N__16650));
    LocalMux I__3389 (
            .O(N__16670),
            .I(RX_ADDR_11));
    LocalMux I__3388 (
            .O(N__16665),
            .I(RX_ADDR_11));
    LocalMux I__3387 (
            .O(N__16662),
            .I(RX_ADDR_11));
    LocalMux I__3386 (
            .O(N__16657),
            .I(RX_ADDR_11));
    LocalMux I__3385 (
            .O(N__16650),
            .I(RX_ADDR_11));
    SRMux I__3384 (
            .O(N__16639),
            .I(N__16635));
    SRMux I__3383 (
            .O(N__16638),
            .I(N__16631));
    LocalMux I__3382 (
            .O(N__16635),
            .I(N__16628));
    SRMux I__3381 (
            .O(N__16634),
            .I(N__16625));
    LocalMux I__3380 (
            .O(N__16631),
            .I(N__16621));
    Span4Mux_h I__3379 (
            .O(N__16628),
            .I(N__16618));
    LocalMux I__3378 (
            .O(N__16625),
            .I(N__16615));
    SRMux I__3377 (
            .O(N__16624),
            .I(N__16612));
    Span4Mux_h I__3376 (
            .O(N__16621),
            .I(N__16609));
    Span4Mux_v I__3375 (
            .O(N__16618),
            .I(N__16604));
    Span4Mux_h I__3374 (
            .O(N__16615),
            .I(N__16604));
    LocalMux I__3373 (
            .O(N__16612),
            .I(N__16601));
    Span4Mux_v I__3372 (
            .O(N__16609),
            .I(N__16598));
    Sp12to4 I__3371 (
            .O(N__16604),
            .I(N__16595));
    Span4Mux_v I__3370 (
            .O(N__16601),
            .I(N__16592));
    Sp12to4 I__3369 (
            .O(N__16598),
            .I(N__16587));
    Span12Mux_s7_v I__3368 (
            .O(N__16595),
            .I(N__16587));
    Span4Mux_h I__3367 (
            .O(N__16592),
            .I(N__16584));
    Span12Mux_v I__3366 (
            .O(N__16587),
            .I(N__16581));
    Span4Mux_h I__3365 (
            .O(N__16584),
            .I(N__16578));
    Odrv12 I__3364 (
            .O(N__16581),
            .I(\line_buffer.n580 ));
    Odrv4 I__3363 (
            .O(N__16578),
            .I(\line_buffer.n580 ));
    InMux I__3362 (
            .O(N__16573),
            .I(N__16570));
    LocalMux I__3361 (
            .O(N__16570),
            .I(N__16567));
    Span4Mux_v I__3360 (
            .O(N__16567),
            .I(N__16564));
    Span4Mux_h I__3359 (
            .O(N__16564),
            .I(N__16561));
    Span4Mux_h I__3358 (
            .O(N__16561),
            .I(N__16558));
    Odrv4 I__3357 (
            .O(N__16558),
            .I(\line_buffer.n511 ));
    InMux I__3356 (
            .O(N__16555),
            .I(N__16552));
    LocalMux I__3355 (
            .O(N__16552),
            .I(N__16549));
    Span12Mux_h I__3354 (
            .O(N__16549),
            .I(N__16546));
    Odrv12 I__3353 (
            .O(N__16546),
            .I(\line_buffer.n503 ));
    InMux I__3352 (
            .O(N__16543),
            .I(N__16540));
    LocalMux I__3351 (
            .O(N__16540),
            .I(N__16537));
    Span4Mux_v I__3350 (
            .O(N__16537),
            .I(N__16534));
    Span4Mux_h I__3349 (
            .O(N__16534),
            .I(N__16531));
    Span4Mux_h I__3348 (
            .O(N__16531),
            .I(N__16528));
    Odrv4 I__3347 (
            .O(N__16528),
            .I(\line_buffer.n509 ));
    InMux I__3346 (
            .O(N__16525),
            .I(N__16522));
    LocalMux I__3345 (
            .O(N__16522),
            .I(N__16519));
    Span4Mux_v I__3344 (
            .O(N__16519),
            .I(N__16516));
    Sp12to4 I__3343 (
            .O(N__16516),
            .I(N__16513));
    Odrv12 I__3342 (
            .O(N__16513),
            .I(\line_buffer.n501 ));
    CascadeMux I__3341 (
            .O(N__16510),
            .I(\receive_module.rx_counter.n4_cascade_ ));
    CascadeMux I__3340 (
            .O(N__16507),
            .I(\receive_module.rx_counter.n6_cascade_ ));
    InMux I__3339 (
            .O(N__16504),
            .I(N__16501));
    LocalMux I__3338 (
            .O(N__16501),
            .I(\receive_module.rx_counter.n3534 ));
    InMux I__3337 (
            .O(N__16498),
            .I(N__16495));
    LocalMux I__3336 (
            .O(N__16495),
            .I(\receive_module.rx_counter.n3581 ));
    SRMux I__3335 (
            .O(N__16492),
            .I(N__16487));
    SRMux I__3334 (
            .O(N__16491),
            .I(N__16484));
    SRMux I__3333 (
            .O(N__16490),
            .I(N__16480));
    LocalMux I__3332 (
            .O(N__16487),
            .I(N__16475));
    LocalMux I__3331 (
            .O(N__16484),
            .I(N__16475));
    SRMux I__3330 (
            .O(N__16483),
            .I(N__16472));
    LocalMux I__3329 (
            .O(N__16480),
            .I(N__16469));
    Span4Mux_s3_v I__3328 (
            .O(N__16475),
            .I(N__16464));
    LocalMux I__3327 (
            .O(N__16472),
            .I(N__16464));
    Sp12to4 I__3326 (
            .O(N__16469),
            .I(N__16461));
    Sp12to4 I__3325 (
            .O(N__16464),
            .I(N__16458));
    Span12Mux_h I__3324 (
            .O(N__16461),
            .I(N__16455));
    Span12Mux_s10_v I__3323 (
            .O(N__16458),
            .I(N__16452));
    Odrv12 I__3322 (
            .O(N__16455),
            .I(\line_buffer.n517 ));
    Odrv12 I__3321 (
            .O(N__16452),
            .I(\line_buffer.n517 ));
    SRMux I__3320 (
            .O(N__16447),
            .I(N__16443));
    SRMux I__3319 (
            .O(N__16446),
            .I(N__16440));
    LocalMux I__3318 (
            .O(N__16443),
            .I(N__16433));
    LocalMux I__3317 (
            .O(N__16440),
            .I(N__16433));
    SRMux I__3316 (
            .O(N__16439),
            .I(N__16430));
    SRMux I__3315 (
            .O(N__16438),
            .I(N__16427));
    Span4Mux_v I__3314 (
            .O(N__16433),
            .I(N__16420));
    LocalMux I__3313 (
            .O(N__16430),
            .I(N__16420));
    LocalMux I__3312 (
            .O(N__16427),
            .I(N__16420));
    Span4Mux_v I__3311 (
            .O(N__16420),
            .I(N__16417));
    Span4Mux_h I__3310 (
            .O(N__16417),
            .I(N__16414));
    Span4Mux_h I__3309 (
            .O(N__16414),
            .I(N__16411));
    Span4Mux_v I__3308 (
            .O(N__16411),
            .I(N__16408));
    Odrv4 I__3307 (
            .O(N__16408),
            .I(\line_buffer.n452 ));
    SRMux I__3306 (
            .O(N__16405),
            .I(N__16401));
    SRMux I__3305 (
            .O(N__16404),
            .I(N__16398));
    LocalMux I__3304 (
            .O(N__16401),
            .I(N__16391));
    LocalMux I__3303 (
            .O(N__16398),
            .I(N__16391));
    SRMux I__3302 (
            .O(N__16397),
            .I(N__16388));
    SRMux I__3301 (
            .O(N__16396),
            .I(N__16385));
    Span4Mux_v I__3300 (
            .O(N__16391),
            .I(N__16380));
    LocalMux I__3299 (
            .O(N__16388),
            .I(N__16380));
    LocalMux I__3298 (
            .O(N__16385),
            .I(N__16377));
    Span4Mux_h I__3297 (
            .O(N__16380),
            .I(N__16374));
    Sp12to4 I__3296 (
            .O(N__16377),
            .I(N__16371));
    Span4Mux_h I__3295 (
            .O(N__16374),
            .I(N__16368));
    Span12Mux_h I__3294 (
            .O(N__16371),
            .I(N__16365));
    Span4Mux_h I__3293 (
            .O(N__16368),
            .I(N__16362));
    Odrv12 I__3292 (
            .O(N__16365),
            .I(\line_buffer.n548 ));
    Odrv4 I__3291 (
            .O(N__16362),
            .I(\line_buffer.n548 ));
    InMux I__3290 (
            .O(N__16357),
            .I(N__16353));
    InMux I__3289 (
            .O(N__16356),
            .I(N__16350));
    LocalMux I__3288 (
            .O(N__16353),
            .I(\receive_module.rx_counter.FRAME_COUNTER_0 ));
    LocalMux I__3287 (
            .O(N__16350),
            .I(\receive_module.rx_counter.FRAME_COUNTER_0 ));
    InMux I__3286 (
            .O(N__16345),
            .I(bfn_16_5_0_));
    InMux I__3285 (
            .O(N__16342),
            .I(N__16338));
    InMux I__3284 (
            .O(N__16341),
            .I(N__16335));
    LocalMux I__3283 (
            .O(N__16338),
            .I(\receive_module.rx_counter.FRAME_COUNTER_1 ));
    LocalMux I__3282 (
            .O(N__16335),
            .I(\receive_module.rx_counter.FRAME_COUNTER_1 ));
    InMux I__3281 (
            .O(N__16330),
            .I(\receive_module.rx_counter.n3310 ));
    InMux I__3280 (
            .O(N__16327),
            .I(N__16323));
    InMux I__3279 (
            .O(N__16326),
            .I(N__16320));
    LocalMux I__3278 (
            .O(N__16323),
            .I(\receive_module.rx_counter.FRAME_COUNTER_2 ));
    LocalMux I__3277 (
            .O(N__16320),
            .I(\receive_module.rx_counter.FRAME_COUNTER_2 ));
    InMux I__3276 (
            .O(N__16315),
            .I(\receive_module.rx_counter.n3311 ));
    InMux I__3275 (
            .O(N__16312),
            .I(N__16308));
    InMux I__3274 (
            .O(N__16311),
            .I(N__16305));
    LocalMux I__3273 (
            .O(N__16308),
            .I(\receive_module.rx_counter.FRAME_COUNTER_3 ));
    LocalMux I__3272 (
            .O(N__16305),
            .I(\receive_module.rx_counter.FRAME_COUNTER_3 ));
    InMux I__3271 (
            .O(N__16300),
            .I(\receive_module.rx_counter.n3312 ));
    InMux I__3270 (
            .O(N__16297),
            .I(N__16293));
    InMux I__3269 (
            .O(N__16296),
            .I(N__16290));
    LocalMux I__3268 (
            .O(N__16293),
            .I(\receive_module.rx_counter.FRAME_COUNTER_4 ));
    LocalMux I__3267 (
            .O(N__16290),
            .I(\receive_module.rx_counter.FRAME_COUNTER_4 ));
    InMux I__3266 (
            .O(N__16285),
            .I(\receive_module.rx_counter.n3313 ));
    InMux I__3265 (
            .O(N__16282),
            .I(\receive_module.rx_counter.n3314 ));
    InMux I__3264 (
            .O(N__16279),
            .I(N__16275));
    InMux I__3263 (
            .O(N__16278),
            .I(N__16272));
    LocalMux I__3262 (
            .O(N__16275),
            .I(\receive_module.rx_counter.FRAME_COUNTER_5 ));
    LocalMux I__3261 (
            .O(N__16272),
            .I(\receive_module.rx_counter.FRAME_COUNTER_5 ));
    CEMux I__3260 (
            .O(N__16267),
            .I(N__16263));
    CEMux I__3259 (
            .O(N__16266),
            .I(N__16260));
    LocalMux I__3258 (
            .O(N__16263),
            .I(N__16257));
    LocalMux I__3257 (
            .O(N__16260),
            .I(N__16254));
    Span4Mux_v I__3256 (
            .O(N__16257),
            .I(N__16251));
    Span4Mux_h I__3255 (
            .O(N__16254),
            .I(N__16248));
    Odrv4 I__3254 (
            .O(N__16251),
            .I(\receive_module.rx_counter.n3792 ));
    Odrv4 I__3253 (
            .O(N__16248),
            .I(\receive_module.rx_counter.n3792 ));
    SRMux I__3252 (
            .O(N__16243),
            .I(N__16240));
    LocalMux I__3251 (
            .O(N__16240),
            .I(N__16237));
    Span4Mux_h I__3250 (
            .O(N__16237),
            .I(N__16234));
    Odrv4 I__3249 (
            .O(N__16234),
            .I(\receive_module.rx_counter.n2517 ));
    InMux I__3248 (
            .O(N__16231),
            .I(N__16228));
    LocalMux I__3247 (
            .O(N__16228),
            .I(N__16225));
    Span4Mux_h I__3246 (
            .O(N__16225),
            .I(N__16222));
    Odrv4 I__3245 (
            .O(N__16222),
            .I(\receive_module.n136 ));
    CascadeMux I__3244 (
            .O(N__16219),
            .I(N__16216));
    CascadeBuf I__3243 (
            .O(N__16216),
            .I(N__16212));
    CascadeMux I__3242 (
            .O(N__16215),
            .I(N__16209));
    CascadeMux I__3241 (
            .O(N__16212),
            .I(N__16206));
    CascadeBuf I__3240 (
            .O(N__16209),
            .I(N__16203));
    CascadeBuf I__3239 (
            .O(N__16206),
            .I(N__16200));
    CascadeMux I__3238 (
            .O(N__16203),
            .I(N__16197));
    CascadeMux I__3237 (
            .O(N__16200),
            .I(N__16194));
    CascadeBuf I__3236 (
            .O(N__16197),
            .I(N__16191));
    CascadeBuf I__3235 (
            .O(N__16194),
            .I(N__16188));
    CascadeMux I__3234 (
            .O(N__16191),
            .I(N__16185));
    CascadeMux I__3233 (
            .O(N__16188),
            .I(N__16182));
    CascadeBuf I__3232 (
            .O(N__16185),
            .I(N__16179));
    CascadeBuf I__3231 (
            .O(N__16182),
            .I(N__16176));
    CascadeMux I__3230 (
            .O(N__16179),
            .I(N__16173));
    CascadeMux I__3229 (
            .O(N__16176),
            .I(N__16170));
    CascadeBuf I__3228 (
            .O(N__16173),
            .I(N__16167));
    CascadeBuf I__3227 (
            .O(N__16170),
            .I(N__16164));
    CascadeMux I__3226 (
            .O(N__16167),
            .I(N__16161));
    CascadeMux I__3225 (
            .O(N__16164),
            .I(N__16158));
    CascadeBuf I__3224 (
            .O(N__16161),
            .I(N__16155));
    CascadeBuf I__3223 (
            .O(N__16158),
            .I(N__16152));
    CascadeMux I__3222 (
            .O(N__16155),
            .I(N__16149));
    CascadeMux I__3221 (
            .O(N__16152),
            .I(N__16146));
    CascadeBuf I__3220 (
            .O(N__16149),
            .I(N__16143));
    CascadeBuf I__3219 (
            .O(N__16146),
            .I(N__16140));
    CascadeMux I__3218 (
            .O(N__16143),
            .I(N__16137));
    CascadeMux I__3217 (
            .O(N__16140),
            .I(N__16134));
    CascadeBuf I__3216 (
            .O(N__16137),
            .I(N__16131));
    CascadeBuf I__3215 (
            .O(N__16134),
            .I(N__16128));
    CascadeMux I__3214 (
            .O(N__16131),
            .I(N__16125));
    CascadeMux I__3213 (
            .O(N__16128),
            .I(N__16122));
    CascadeBuf I__3212 (
            .O(N__16125),
            .I(N__16119));
    CascadeBuf I__3211 (
            .O(N__16122),
            .I(N__16116));
    CascadeMux I__3210 (
            .O(N__16119),
            .I(N__16113));
    CascadeMux I__3209 (
            .O(N__16116),
            .I(N__16110));
    CascadeBuf I__3208 (
            .O(N__16113),
            .I(N__16107));
    CascadeBuf I__3207 (
            .O(N__16110),
            .I(N__16104));
    CascadeMux I__3206 (
            .O(N__16107),
            .I(N__16101));
    CascadeMux I__3205 (
            .O(N__16104),
            .I(N__16098));
    CascadeBuf I__3204 (
            .O(N__16101),
            .I(N__16095));
    CascadeBuf I__3203 (
            .O(N__16098),
            .I(N__16092));
    CascadeMux I__3202 (
            .O(N__16095),
            .I(N__16089));
    CascadeMux I__3201 (
            .O(N__16092),
            .I(N__16086));
    CascadeBuf I__3200 (
            .O(N__16089),
            .I(N__16083));
    CascadeBuf I__3199 (
            .O(N__16086),
            .I(N__16080));
    CascadeMux I__3198 (
            .O(N__16083),
            .I(N__16077));
    CascadeMux I__3197 (
            .O(N__16080),
            .I(N__16074));
    CascadeBuf I__3196 (
            .O(N__16077),
            .I(N__16071));
    CascadeBuf I__3195 (
            .O(N__16074),
            .I(N__16068));
    CascadeMux I__3194 (
            .O(N__16071),
            .I(N__16065));
    CascadeMux I__3193 (
            .O(N__16068),
            .I(N__16062));
    CascadeBuf I__3192 (
            .O(N__16065),
            .I(N__16059));
    CascadeBuf I__3191 (
            .O(N__16062),
            .I(N__16056));
    CascadeMux I__3190 (
            .O(N__16059),
            .I(N__16053));
    CascadeMux I__3189 (
            .O(N__16056),
            .I(N__16050));
    CascadeBuf I__3188 (
            .O(N__16053),
            .I(N__16047));
    CascadeBuf I__3187 (
            .O(N__16050),
            .I(N__16044));
    CascadeMux I__3186 (
            .O(N__16047),
            .I(N__16041));
    CascadeMux I__3185 (
            .O(N__16044),
            .I(N__16038));
    CascadeBuf I__3184 (
            .O(N__16041),
            .I(N__16035));
    InMux I__3183 (
            .O(N__16038),
            .I(N__16032));
    CascadeMux I__3182 (
            .O(N__16035),
            .I(N__16029));
    LocalMux I__3181 (
            .O(N__16032),
            .I(N__16026));
    InMux I__3180 (
            .O(N__16029),
            .I(N__16023));
    Span4Mux_s1_v I__3179 (
            .O(N__16026),
            .I(N__16020));
    LocalMux I__3178 (
            .O(N__16023),
            .I(N__16017));
    Span4Mux_h I__3177 (
            .O(N__16020),
            .I(N__16014));
    Span4Mux_s1_v I__3176 (
            .O(N__16017),
            .I(N__16011));
    Span4Mux_h I__3175 (
            .O(N__16014),
            .I(N__16007));
    Span4Mux_v I__3174 (
            .O(N__16011),
            .I(N__16004));
    InMux I__3173 (
            .O(N__16010),
            .I(N__16001));
    Span4Mux_v I__3172 (
            .O(N__16007),
            .I(N__15998));
    Sp12to4 I__3171 (
            .O(N__16004),
            .I(N__15995));
    LocalMux I__3170 (
            .O(N__16001),
            .I(N__15991));
    Sp12to4 I__3169 (
            .O(N__15998),
            .I(N__15986));
    Span12Mux_h I__3168 (
            .O(N__15995),
            .I(N__15986));
    InMux I__3167 (
            .O(N__15994),
            .I(N__15983));
    Sp12to4 I__3166 (
            .O(N__15991),
            .I(N__15978));
    Span12Mux_v I__3165 (
            .O(N__15986),
            .I(N__15978));
    LocalMux I__3164 (
            .O(N__15983),
            .I(RX_ADDR_0));
    Odrv12 I__3163 (
            .O(N__15978),
            .I(RX_ADDR_0));
    CascadeMux I__3162 (
            .O(N__15973),
            .I(N__15970));
    InMux I__3161 (
            .O(N__15970),
            .I(N__15967));
    LocalMux I__3160 (
            .O(N__15967),
            .I(N__15964));
    Span4Mux_h I__3159 (
            .O(N__15964),
            .I(N__15961));
    Odrv4 I__3158 (
            .O(N__15961),
            .I(\receive_module.n135 ));
    CascadeMux I__3157 (
            .O(N__15958),
            .I(N__15954));
    CascadeMux I__3156 (
            .O(N__15957),
            .I(N__15951));
    CascadeBuf I__3155 (
            .O(N__15954),
            .I(N__15948));
    CascadeBuf I__3154 (
            .O(N__15951),
            .I(N__15945));
    CascadeMux I__3153 (
            .O(N__15948),
            .I(N__15942));
    CascadeMux I__3152 (
            .O(N__15945),
            .I(N__15939));
    CascadeBuf I__3151 (
            .O(N__15942),
            .I(N__15936));
    CascadeBuf I__3150 (
            .O(N__15939),
            .I(N__15933));
    CascadeMux I__3149 (
            .O(N__15936),
            .I(N__15930));
    CascadeMux I__3148 (
            .O(N__15933),
            .I(N__15927));
    CascadeBuf I__3147 (
            .O(N__15930),
            .I(N__15924));
    CascadeBuf I__3146 (
            .O(N__15927),
            .I(N__15921));
    CascadeMux I__3145 (
            .O(N__15924),
            .I(N__15918));
    CascadeMux I__3144 (
            .O(N__15921),
            .I(N__15915));
    CascadeBuf I__3143 (
            .O(N__15918),
            .I(N__15912));
    CascadeBuf I__3142 (
            .O(N__15915),
            .I(N__15909));
    CascadeMux I__3141 (
            .O(N__15912),
            .I(N__15906));
    CascadeMux I__3140 (
            .O(N__15909),
            .I(N__15903));
    CascadeBuf I__3139 (
            .O(N__15906),
            .I(N__15900));
    CascadeBuf I__3138 (
            .O(N__15903),
            .I(N__15897));
    CascadeMux I__3137 (
            .O(N__15900),
            .I(N__15894));
    CascadeMux I__3136 (
            .O(N__15897),
            .I(N__15891));
    CascadeBuf I__3135 (
            .O(N__15894),
            .I(N__15888));
    CascadeBuf I__3134 (
            .O(N__15891),
            .I(N__15885));
    CascadeMux I__3133 (
            .O(N__15888),
            .I(N__15882));
    CascadeMux I__3132 (
            .O(N__15885),
            .I(N__15879));
    CascadeBuf I__3131 (
            .O(N__15882),
            .I(N__15876));
    CascadeBuf I__3130 (
            .O(N__15879),
            .I(N__15873));
    CascadeMux I__3129 (
            .O(N__15876),
            .I(N__15870));
    CascadeMux I__3128 (
            .O(N__15873),
            .I(N__15867));
    CascadeBuf I__3127 (
            .O(N__15870),
            .I(N__15864));
    CascadeBuf I__3126 (
            .O(N__15867),
            .I(N__15861));
    CascadeMux I__3125 (
            .O(N__15864),
            .I(N__15858));
    CascadeMux I__3124 (
            .O(N__15861),
            .I(N__15855));
    CascadeBuf I__3123 (
            .O(N__15858),
            .I(N__15852));
    CascadeBuf I__3122 (
            .O(N__15855),
            .I(N__15849));
    CascadeMux I__3121 (
            .O(N__15852),
            .I(N__15846));
    CascadeMux I__3120 (
            .O(N__15849),
            .I(N__15843));
    CascadeBuf I__3119 (
            .O(N__15846),
            .I(N__15840));
    CascadeBuf I__3118 (
            .O(N__15843),
            .I(N__15837));
    CascadeMux I__3117 (
            .O(N__15840),
            .I(N__15834));
    CascadeMux I__3116 (
            .O(N__15837),
            .I(N__15831));
    CascadeBuf I__3115 (
            .O(N__15834),
            .I(N__15828));
    CascadeBuf I__3114 (
            .O(N__15831),
            .I(N__15825));
    CascadeMux I__3113 (
            .O(N__15828),
            .I(N__15822));
    CascadeMux I__3112 (
            .O(N__15825),
            .I(N__15819));
    CascadeBuf I__3111 (
            .O(N__15822),
            .I(N__15816));
    CascadeBuf I__3110 (
            .O(N__15819),
            .I(N__15813));
    CascadeMux I__3109 (
            .O(N__15816),
            .I(N__15810));
    CascadeMux I__3108 (
            .O(N__15813),
            .I(N__15807));
    CascadeBuf I__3107 (
            .O(N__15810),
            .I(N__15804));
    CascadeBuf I__3106 (
            .O(N__15807),
            .I(N__15801));
    CascadeMux I__3105 (
            .O(N__15804),
            .I(N__15798));
    CascadeMux I__3104 (
            .O(N__15801),
            .I(N__15795));
    CascadeBuf I__3103 (
            .O(N__15798),
            .I(N__15792));
    CascadeBuf I__3102 (
            .O(N__15795),
            .I(N__15789));
    CascadeMux I__3101 (
            .O(N__15792),
            .I(N__15786));
    CascadeMux I__3100 (
            .O(N__15789),
            .I(N__15783));
    CascadeBuf I__3099 (
            .O(N__15786),
            .I(N__15780));
    CascadeBuf I__3098 (
            .O(N__15783),
            .I(N__15777));
    CascadeMux I__3097 (
            .O(N__15780),
            .I(N__15774));
    CascadeMux I__3096 (
            .O(N__15777),
            .I(N__15771));
    InMux I__3095 (
            .O(N__15774),
            .I(N__15768));
    InMux I__3094 (
            .O(N__15771),
            .I(N__15765));
    LocalMux I__3093 (
            .O(N__15768),
            .I(N__15762));
    LocalMux I__3092 (
            .O(N__15765),
            .I(N__15759));
    Span4Mux_h I__3091 (
            .O(N__15762),
            .I(N__15755));
    Span4Mux_h I__3090 (
            .O(N__15759),
            .I(N__15752));
    InMux I__3089 (
            .O(N__15758),
            .I(N__15748));
    Sp12to4 I__3088 (
            .O(N__15755),
            .I(N__15745));
    Sp12to4 I__3087 (
            .O(N__15752),
            .I(N__15742));
    InMux I__3086 (
            .O(N__15751),
            .I(N__15739));
    LocalMux I__3085 (
            .O(N__15748),
            .I(N__15736));
    Span12Mux_v I__3084 (
            .O(N__15745),
            .I(N__15733));
    Span12Mux_v I__3083 (
            .O(N__15742),
            .I(N__15730));
    LocalMux I__3082 (
            .O(N__15739),
            .I(N__15725));
    Span4Mux_v I__3081 (
            .O(N__15736),
            .I(N__15725));
    Span12Mux_v I__3080 (
            .O(N__15733),
            .I(N__15720));
    Span12Mux_v I__3079 (
            .O(N__15730),
            .I(N__15720));
    Odrv4 I__3078 (
            .O(N__15725),
            .I(RX_ADDR_1));
    Odrv12 I__3077 (
            .O(N__15720),
            .I(RX_ADDR_1));
    InMux I__3076 (
            .O(N__15715),
            .I(N__15712));
    LocalMux I__3075 (
            .O(N__15712),
            .I(N__15709));
    Span4Mux_v I__3074 (
            .O(N__15709),
            .I(N__15706));
    Span4Mux_h I__3073 (
            .O(N__15706),
            .I(N__15703));
    Odrv4 I__3072 (
            .O(N__15703),
            .I(\line_buffer.n545 ));
    InMux I__3071 (
            .O(N__15700),
            .I(N__15697));
    LocalMux I__3070 (
            .O(N__15697),
            .I(N__15694));
    Span4Mux_v I__3069 (
            .O(N__15694),
            .I(N__15691));
    Sp12to4 I__3068 (
            .O(N__15691),
            .I(N__15688));
    Span12Mux_h I__3067 (
            .O(N__15688),
            .I(N__15685));
    Span12Mux_v I__3066 (
            .O(N__15685),
            .I(N__15682));
    Odrv12 I__3065 (
            .O(N__15682),
            .I(\line_buffer.n537 ));
    InMux I__3064 (
            .O(N__15679),
            .I(N__15676));
    LocalMux I__3063 (
            .O(N__15676),
            .I(\line_buffer.n3680 ));
    InMux I__3062 (
            .O(N__15673),
            .I(N__15670));
    LocalMux I__3061 (
            .O(N__15670),
            .I(N__15667));
    Span12Mux_s10_v I__3060 (
            .O(N__15667),
            .I(N__15664));
    Odrv12 I__3059 (
            .O(N__15664),
            .I(\receive_module.n126 ));
    CascadeMux I__3058 (
            .O(N__15661),
            .I(N__15658));
    CascadeBuf I__3057 (
            .O(N__15658),
            .I(N__15654));
    CascadeMux I__3056 (
            .O(N__15657),
            .I(N__15651));
    CascadeMux I__3055 (
            .O(N__15654),
            .I(N__15648));
    CascadeBuf I__3054 (
            .O(N__15651),
            .I(N__15645));
    CascadeBuf I__3053 (
            .O(N__15648),
            .I(N__15642));
    CascadeMux I__3052 (
            .O(N__15645),
            .I(N__15639));
    CascadeMux I__3051 (
            .O(N__15642),
            .I(N__15636));
    CascadeBuf I__3050 (
            .O(N__15639),
            .I(N__15633));
    CascadeBuf I__3049 (
            .O(N__15636),
            .I(N__15630));
    CascadeMux I__3048 (
            .O(N__15633),
            .I(N__15627));
    CascadeMux I__3047 (
            .O(N__15630),
            .I(N__15624));
    CascadeBuf I__3046 (
            .O(N__15627),
            .I(N__15621));
    CascadeBuf I__3045 (
            .O(N__15624),
            .I(N__15618));
    CascadeMux I__3044 (
            .O(N__15621),
            .I(N__15615));
    CascadeMux I__3043 (
            .O(N__15618),
            .I(N__15612));
    CascadeBuf I__3042 (
            .O(N__15615),
            .I(N__15609));
    CascadeBuf I__3041 (
            .O(N__15612),
            .I(N__15606));
    CascadeMux I__3040 (
            .O(N__15609),
            .I(N__15603));
    CascadeMux I__3039 (
            .O(N__15606),
            .I(N__15600));
    CascadeBuf I__3038 (
            .O(N__15603),
            .I(N__15597));
    CascadeBuf I__3037 (
            .O(N__15600),
            .I(N__15594));
    CascadeMux I__3036 (
            .O(N__15597),
            .I(N__15591));
    CascadeMux I__3035 (
            .O(N__15594),
            .I(N__15588));
    CascadeBuf I__3034 (
            .O(N__15591),
            .I(N__15585));
    CascadeBuf I__3033 (
            .O(N__15588),
            .I(N__15582));
    CascadeMux I__3032 (
            .O(N__15585),
            .I(N__15579));
    CascadeMux I__3031 (
            .O(N__15582),
            .I(N__15576));
    CascadeBuf I__3030 (
            .O(N__15579),
            .I(N__15573));
    CascadeBuf I__3029 (
            .O(N__15576),
            .I(N__15570));
    CascadeMux I__3028 (
            .O(N__15573),
            .I(N__15567));
    CascadeMux I__3027 (
            .O(N__15570),
            .I(N__15564));
    CascadeBuf I__3026 (
            .O(N__15567),
            .I(N__15561));
    CascadeBuf I__3025 (
            .O(N__15564),
            .I(N__15558));
    CascadeMux I__3024 (
            .O(N__15561),
            .I(N__15555));
    CascadeMux I__3023 (
            .O(N__15558),
            .I(N__15552));
    CascadeBuf I__3022 (
            .O(N__15555),
            .I(N__15549));
    CascadeBuf I__3021 (
            .O(N__15552),
            .I(N__15546));
    CascadeMux I__3020 (
            .O(N__15549),
            .I(N__15543));
    CascadeMux I__3019 (
            .O(N__15546),
            .I(N__15540));
    CascadeBuf I__3018 (
            .O(N__15543),
            .I(N__15537));
    CascadeBuf I__3017 (
            .O(N__15540),
            .I(N__15534));
    CascadeMux I__3016 (
            .O(N__15537),
            .I(N__15531));
    CascadeMux I__3015 (
            .O(N__15534),
            .I(N__15528));
    CascadeBuf I__3014 (
            .O(N__15531),
            .I(N__15525));
    CascadeBuf I__3013 (
            .O(N__15528),
            .I(N__15522));
    CascadeMux I__3012 (
            .O(N__15525),
            .I(N__15519));
    CascadeMux I__3011 (
            .O(N__15522),
            .I(N__15516));
    CascadeBuf I__3010 (
            .O(N__15519),
            .I(N__15513));
    CascadeBuf I__3009 (
            .O(N__15516),
            .I(N__15510));
    CascadeMux I__3008 (
            .O(N__15513),
            .I(N__15507));
    CascadeMux I__3007 (
            .O(N__15510),
            .I(N__15504));
    CascadeBuf I__3006 (
            .O(N__15507),
            .I(N__15501));
    CascadeBuf I__3005 (
            .O(N__15504),
            .I(N__15498));
    CascadeMux I__3004 (
            .O(N__15501),
            .I(N__15495));
    CascadeMux I__3003 (
            .O(N__15498),
            .I(N__15492));
    CascadeBuf I__3002 (
            .O(N__15495),
            .I(N__15489));
    CascadeBuf I__3001 (
            .O(N__15492),
            .I(N__15486));
    CascadeMux I__3000 (
            .O(N__15489),
            .I(N__15483));
    CascadeMux I__2999 (
            .O(N__15486),
            .I(N__15480));
    CascadeBuf I__2998 (
            .O(N__15483),
            .I(N__15476));
    InMux I__2997 (
            .O(N__15480),
            .I(N__15473));
    InMux I__2996 (
            .O(N__15479),
            .I(N__15470));
    CascadeMux I__2995 (
            .O(N__15476),
            .I(N__15467));
    LocalMux I__2994 (
            .O(N__15473),
            .I(N__15464));
    LocalMux I__2993 (
            .O(N__15470),
            .I(N__15461));
    InMux I__2992 (
            .O(N__15467),
            .I(N__15458));
    Span4Mux_s1_v I__2991 (
            .O(N__15464),
            .I(N__15455));
    Span4Mux_h I__2990 (
            .O(N__15461),
            .I(N__15452));
    LocalMux I__2989 (
            .O(N__15458),
            .I(N__15449));
    Span4Mux_h I__2988 (
            .O(N__15455),
            .I(N__15446));
    Span4Mux_v I__2987 (
            .O(N__15452),
            .I(N__15443));
    Sp12to4 I__2986 (
            .O(N__15449),
            .I(N__15439));
    Span4Mux_v I__2985 (
            .O(N__15446),
            .I(N__15436));
    Span4Mux_v I__2984 (
            .O(N__15443),
            .I(N__15433));
    InMux I__2983 (
            .O(N__15442),
            .I(N__15430));
    Span12Mux_s9_v I__2982 (
            .O(N__15439),
            .I(N__15427));
    Span4Mux_v I__2981 (
            .O(N__15436),
            .I(N__15424));
    Odrv4 I__2980 (
            .O(N__15433),
            .I(RX_ADDR_10));
    LocalMux I__2979 (
            .O(N__15430),
            .I(RX_ADDR_10));
    Odrv12 I__2978 (
            .O(N__15427),
            .I(RX_ADDR_10));
    Odrv4 I__2977 (
            .O(N__15424),
            .I(RX_ADDR_10));
    InMux I__2976 (
            .O(N__15415),
            .I(N__15412));
    LocalMux I__2975 (
            .O(N__15412),
            .I(N__15409));
    Span12Mux_s5_v I__2974 (
            .O(N__15409),
            .I(N__15406));
    Span12Mux_v I__2973 (
            .O(N__15406),
            .I(N__15403));
    Odrv12 I__2972 (
            .O(N__15403),
            .I(\receive_module.n132 ));
    CascadeMux I__2971 (
            .O(N__15400),
            .I(N__15396));
    CascadeMux I__2970 (
            .O(N__15399),
            .I(N__15393));
    CascadeBuf I__2969 (
            .O(N__15396),
            .I(N__15390));
    CascadeBuf I__2968 (
            .O(N__15393),
            .I(N__15387));
    CascadeMux I__2967 (
            .O(N__15390),
            .I(N__15384));
    CascadeMux I__2966 (
            .O(N__15387),
            .I(N__15381));
    CascadeBuf I__2965 (
            .O(N__15384),
            .I(N__15378));
    CascadeBuf I__2964 (
            .O(N__15381),
            .I(N__15375));
    CascadeMux I__2963 (
            .O(N__15378),
            .I(N__15372));
    CascadeMux I__2962 (
            .O(N__15375),
            .I(N__15369));
    CascadeBuf I__2961 (
            .O(N__15372),
            .I(N__15366));
    CascadeBuf I__2960 (
            .O(N__15369),
            .I(N__15363));
    CascadeMux I__2959 (
            .O(N__15366),
            .I(N__15360));
    CascadeMux I__2958 (
            .O(N__15363),
            .I(N__15357));
    CascadeBuf I__2957 (
            .O(N__15360),
            .I(N__15354));
    CascadeBuf I__2956 (
            .O(N__15357),
            .I(N__15351));
    CascadeMux I__2955 (
            .O(N__15354),
            .I(N__15348));
    CascadeMux I__2954 (
            .O(N__15351),
            .I(N__15345));
    CascadeBuf I__2953 (
            .O(N__15348),
            .I(N__15342));
    CascadeBuf I__2952 (
            .O(N__15345),
            .I(N__15339));
    CascadeMux I__2951 (
            .O(N__15342),
            .I(N__15336));
    CascadeMux I__2950 (
            .O(N__15339),
            .I(N__15333));
    CascadeBuf I__2949 (
            .O(N__15336),
            .I(N__15330));
    CascadeBuf I__2948 (
            .O(N__15333),
            .I(N__15327));
    CascadeMux I__2947 (
            .O(N__15330),
            .I(N__15324));
    CascadeMux I__2946 (
            .O(N__15327),
            .I(N__15321));
    CascadeBuf I__2945 (
            .O(N__15324),
            .I(N__15318));
    CascadeBuf I__2944 (
            .O(N__15321),
            .I(N__15315));
    CascadeMux I__2943 (
            .O(N__15318),
            .I(N__15312));
    CascadeMux I__2942 (
            .O(N__15315),
            .I(N__15309));
    CascadeBuf I__2941 (
            .O(N__15312),
            .I(N__15306));
    CascadeBuf I__2940 (
            .O(N__15309),
            .I(N__15303));
    CascadeMux I__2939 (
            .O(N__15306),
            .I(N__15300));
    CascadeMux I__2938 (
            .O(N__15303),
            .I(N__15297));
    CascadeBuf I__2937 (
            .O(N__15300),
            .I(N__15294));
    CascadeBuf I__2936 (
            .O(N__15297),
            .I(N__15291));
    CascadeMux I__2935 (
            .O(N__15294),
            .I(N__15288));
    CascadeMux I__2934 (
            .O(N__15291),
            .I(N__15285));
    CascadeBuf I__2933 (
            .O(N__15288),
            .I(N__15282));
    CascadeBuf I__2932 (
            .O(N__15285),
            .I(N__15279));
    CascadeMux I__2931 (
            .O(N__15282),
            .I(N__15276));
    CascadeMux I__2930 (
            .O(N__15279),
            .I(N__15273));
    CascadeBuf I__2929 (
            .O(N__15276),
            .I(N__15270));
    CascadeBuf I__2928 (
            .O(N__15273),
            .I(N__15267));
    CascadeMux I__2927 (
            .O(N__15270),
            .I(N__15264));
    CascadeMux I__2926 (
            .O(N__15267),
            .I(N__15261));
    CascadeBuf I__2925 (
            .O(N__15264),
            .I(N__15258));
    CascadeBuf I__2924 (
            .O(N__15261),
            .I(N__15255));
    CascadeMux I__2923 (
            .O(N__15258),
            .I(N__15252));
    CascadeMux I__2922 (
            .O(N__15255),
            .I(N__15249));
    CascadeBuf I__2921 (
            .O(N__15252),
            .I(N__15246));
    CascadeBuf I__2920 (
            .O(N__15249),
            .I(N__15243));
    CascadeMux I__2919 (
            .O(N__15246),
            .I(N__15240));
    CascadeMux I__2918 (
            .O(N__15243),
            .I(N__15237));
    CascadeBuf I__2917 (
            .O(N__15240),
            .I(N__15234));
    CascadeBuf I__2916 (
            .O(N__15237),
            .I(N__15231));
    CascadeMux I__2915 (
            .O(N__15234),
            .I(N__15228));
    CascadeMux I__2914 (
            .O(N__15231),
            .I(N__15225));
    CascadeBuf I__2913 (
            .O(N__15228),
            .I(N__15222));
    CascadeBuf I__2912 (
            .O(N__15225),
            .I(N__15219));
    CascadeMux I__2911 (
            .O(N__15222),
            .I(N__15215));
    CascadeMux I__2910 (
            .O(N__15219),
            .I(N__15212));
    InMux I__2909 (
            .O(N__15218),
            .I(N__15209));
    InMux I__2908 (
            .O(N__15215),
            .I(N__15206));
    InMux I__2907 (
            .O(N__15212),
            .I(N__15203));
    LocalMux I__2906 (
            .O(N__15209),
            .I(N__15199));
    LocalMux I__2905 (
            .O(N__15206),
            .I(N__15196));
    LocalMux I__2904 (
            .O(N__15203),
            .I(N__15193));
    InMux I__2903 (
            .O(N__15202),
            .I(N__15190));
    Span12Mux_v I__2902 (
            .O(N__15199),
            .I(N__15183));
    Span12Mux_h I__2901 (
            .O(N__15196),
            .I(N__15183));
    Span12Mux_h I__2900 (
            .O(N__15193),
            .I(N__15183));
    LocalMux I__2899 (
            .O(N__15190),
            .I(RX_ADDR_4));
    Odrv12 I__2898 (
            .O(N__15183),
            .I(RX_ADDR_4));
    InMux I__2897 (
            .O(N__15178),
            .I(N__15175));
    LocalMux I__2896 (
            .O(N__15175),
            .I(N__15172));
    Span12Mux_s4_v I__2895 (
            .O(N__15172),
            .I(N__15169));
    Span12Mux_v I__2894 (
            .O(N__15169),
            .I(N__15166));
    Odrv12 I__2893 (
            .O(N__15166),
            .I(\receive_module.n131 ));
    CascadeMux I__2892 (
            .O(N__15163),
            .I(N__15159));
    CascadeMux I__2891 (
            .O(N__15162),
            .I(N__15156));
    CascadeBuf I__2890 (
            .O(N__15159),
            .I(N__15153));
    CascadeBuf I__2889 (
            .O(N__15156),
            .I(N__15150));
    CascadeMux I__2888 (
            .O(N__15153),
            .I(N__15147));
    CascadeMux I__2887 (
            .O(N__15150),
            .I(N__15144));
    CascadeBuf I__2886 (
            .O(N__15147),
            .I(N__15141));
    CascadeBuf I__2885 (
            .O(N__15144),
            .I(N__15138));
    CascadeMux I__2884 (
            .O(N__15141),
            .I(N__15135));
    CascadeMux I__2883 (
            .O(N__15138),
            .I(N__15132));
    CascadeBuf I__2882 (
            .O(N__15135),
            .I(N__15129));
    CascadeBuf I__2881 (
            .O(N__15132),
            .I(N__15126));
    CascadeMux I__2880 (
            .O(N__15129),
            .I(N__15123));
    CascadeMux I__2879 (
            .O(N__15126),
            .I(N__15120));
    CascadeBuf I__2878 (
            .O(N__15123),
            .I(N__15117));
    CascadeBuf I__2877 (
            .O(N__15120),
            .I(N__15114));
    CascadeMux I__2876 (
            .O(N__15117),
            .I(N__15111));
    CascadeMux I__2875 (
            .O(N__15114),
            .I(N__15108));
    CascadeBuf I__2874 (
            .O(N__15111),
            .I(N__15105));
    CascadeBuf I__2873 (
            .O(N__15108),
            .I(N__15102));
    CascadeMux I__2872 (
            .O(N__15105),
            .I(N__15099));
    CascadeMux I__2871 (
            .O(N__15102),
            .I(N__15096));
    CascadeBuf I__2870 (
            .O(N__15099),
            .I(N__15093));
    CascadeBuf I__2869 (
            .O(N__15096),
            .I(N__15090));
    CascadeMux I__2868 (
            .O(N__15093),
            .I(N__15087));
    CascadeMux I__2867 (
            .O(N__15090),
            .I(N__15084));
    CascadeBuf I__2866 (
            .O(N__15087),
            .I(N__15081));
    CascadeBuf I__2865 (
            .O(N__15084),
            .I(N__15078));
    CascadeMux I__2864 (
            .O(N__15081),
            .I(N__15075));
    CascadeMux I__2863 (
            .O(N__15078),
            .I(N__15072));
    CascadeBuf I__2862 (
            .O(N__15075),
            .I(N__15069));
    CascadeBuf I__2861 (
            .O(N__15072),
            .I(N__15066));
    CascadeMux I__2860 (
            .O(N__15069),
            .I(N__15063));
    CascadeMux I__2859 (
            .O(N__15066),
            .I(N__15060));
    CascadeBuf I__2858 (
            .O(N__15063),
            .I(N__15057));
    CascadeBuf I__2857 (
            .O(N__15060),
            .I(N__15054));
    CascadeMux I__2856 (
            .O(N__15057),
            .I(N__15051));
    CascadeMux I__2855 (
            .O(N__15054),
            .I(N__15048));
    CascadeBuf I__2854 (
            .O(N__15051),
            .I(N__15045));
    CascadeBuf I__2853 (
            .O(N__15048),
            .I(N__15042));
    CascadeMux I__2852 (
            .O(N__15045),
            .I(N__15039));
    CascadeMux I__2851 (
            .O(N__15042),
            .I(N__15036));
    CascadeBuf I__2850 (
            .O(N__15039),
            .I(N__15033));
    CascadeBuf I__2849 (
            .O(N__15036),
            .I(N__15030));
    CascadeMux I__2848 (
            .O(N__15033),
            .I(N__15027));
    CascadeMux I__2847 (
            .O(N__15030),
            .I(N__15024));
    CascadeBuf I__2846 (
            .O(N__15027),
            .I(N__15021));
    CascadeBuf I__2845 (
            .O(N__15024),
            .I(N__15018));
    CascadeMux I__2844 (
            .O(N__15021),
            .I(N__15015));
    CascadeMux I__2843 (
            .O(N__15018),
            .I(N__15012));
    CascadeBuf I__2842 (
            .O(N__15015),
            .I(N__15009));
    CascadeBuf I__2841 (
            .O(N__15012),
            .I(N__15006));
    CascadeMux I__2840 (
            .O(N__15009),
            .I(N__15003));
    CascadeMux I__2839 (
            .O(N__15006),
            .I(N__15000));
    CascadeBuf I__2838 (
            .O(N__15003),
            .I(N__14997));
    CascadeBuf I__2837 (
            .O(N__15000),
            .I(N__14994));
    CascadeMux I__2836 (
            .O(N__14997),
            .I(N__14991));
    CascadeMux I__2835 (
            .O(N__14994),
            .I(N__14987));
    CascadeBuf I__2834 (
            .O(N__14991),
            .I(N__14984));
    InMux I__2833 (
            .O(N__14990),
            .I(N__14981));
    CascadeBuf I__2832 (
            .O(N__14987),
            .I(N__14978));
    CascadeMux I__2831 (
            .O(N__14984),
            .I(N__14975));
    LocalMux I__2830 (
            .O(N__14981),
            .I(N__14972));
    CascadeMux I__2829 (
            .O(N__14978),
            .I(N__14969));
    InMux I__2828 (
            .O(N__14975),
            .I(N__14966));
    Span4Mux_v I__2827 (
            .O(N__14972),
            .I(N__14963));
    InMux I__2826 (
            .O(N__14969),
            .I(N__14960));
    LocalMux I__2825 (
            .O(N__14966),
            .I(N__14957));
    Span4Mux_v I__2824 (
            .O(N__14963),
            .I(N__14953));
    LocalMux I__2823 (
            .O(N__14960),
            .I(N__14950));
    Span4Mux_s1_v I__2822 (
            .O(N__14957),
            .I(N__14947));
    CascadeMux I__2821 (
            .O(N__14956),
            .I(N__14944));
    Span4Mux_v I__2820 (
            .O(N__14953),
            .I(N__14941));
    Span4Mux_s1_v I__2819 (
            .O(N__14950),
            .I(N__14938));
    Span4Mux_h I__2818 (
            .O(N__14947),
            .I(N__14935));
    InMux I__2817 (
            .O(N__14944),
            .I(N__14932));
    Sp12to4 I__2816 (
            .O(N__14941),
            .I(N__14929));
    Span4Mux_h I__2815 (
            .O(N__14938),
            .I(N__14926));
    Span4Mux_h I__2814 (
            .O(N__14935),
            .I(N__14923));
    LocalMux I__2813 (
            .O(N__14932),
            .I(RX_ADDR_5));
    Odrv12 I__2812 (
            .O(N__14929),
            .I(RX_ADDR_5));
    Odrv4 I__2811 (
            .O(N__14926),
            .I(RX_ADDR_5));
    Odrv4 I__2810 (
            .O(N__14923),
            .I(RX_ADDR_5));
    InMux I__2809 (
            .O(N__14914),
            .I(N__14911));
    LocalMux I__2808 (
            .O(N__14911),
            .I(N__14908));
    Span12Mux_s3_v I__2807 (
            .O(N__14908),
            .I(N__14905));
    Span12Mux_v I__2806 (
            .O(N__14905),
            .I(N__14902));
    Odrv12 I__2805 (
            .O(N__14902),
            .I(\receive_module.n130 ));
    CascadeMux I__2804 (
            .O(N__14899),
            .I(N__14896));
    CascadeBuf I__2803 (
            .O(N__14896),
            .I(N__14892));
    CascadeMux I__2802 (
            .O(N__14895),
            .I(N__14889));
    CascadeMux I__2801 (
            .O(N__14892),
            .I(N__14886));
    CascadeBuf I__2800 (
            .O(N__14889),
            .I(N__14883));
    CascadeBuf I__2799 (
            .O(N__14886),
            .I(N__14880));
    CascadeMux I__2798 (
            .O(N__14883),
            .I(N__14877));
    CascadeMux I__2797 (
            .O(N__14880),
            .I(N__14874));
    CascadeBuf I__2796 (
            .O(N__14877),
            .I(N__14871));
    CascadeBuf I__2795 (
            .O(N__14874),
            .I(N__14868));
    CascadeMux I__2794 (
            .O(N__14871),
            .I(N__14865));
    CascadeMux I__2793 (
            .O(N__14868),
            .I(N__14862));
    CascadeBuf I__2792 (
            .O(N__14865),
            .I(N__14859));
    CascadeBuf I__2791 (
            .O(N__14862),
            .I(N__14856));
    CascadeMux I__2790 (
            .O(N__14859),
            .I(N__14853));
    CascadeMux I__2789 (
            .O(N__14856),
            .I(N__14850));
    CascadeBuf I__2788 (
            .O(N__14853),
            .I(N__14847));
    CascadeBuf I__2787 (
            .O(N__14850),
            .I(N__14844));
    CascadeMux I__2786 (
            .O(N__14847),
            .I(N__14841));
    CascadeMux I__2785 (
            .O(N__14844),
            .I(N__14838));
    CascadeBuf I__2784 (
            .O(N__14841),
            .I(N__14835));
    CascadeBuf I__2783 (
            .O(N__14838),
            .I(N__14832));
    CascadeMux I__2782 (
            .O(N__14835),
            .I(N__14829));
    CascadeMux I__2781 (
            .O(N__14832),
            .I(N__14826));
    CascadeBuf I__2780 (
            .O(N__14829),
            .I(N__14823));
    CascadeBuf I__2779 (
            .O(N__14826),
            .I(N__14820));
    CascadeMux I__2778 (
            .O(N__14823),
            .I(N__14817));
    CascadeMux I__2777 (
            .O(N__14820),
            .I(N__14814));
    CascadeBuf I__2776 (
            .O(N__14817),
            .I(N__14811));
    CascadeBuf I__2775 (
            .O(N__14814),
            .I(N__14808));
    CascadeMux I__2774 (
            .O(N__14811),
            .I(N__14805));
    CascadeMux I__2773 (
            .O(N__14808),
            .I(N__14802));
    CascadeBuf I__2772 (
            .O(N__14805),
            .I(N__14799));
    CascadeBuf I__2771 (
            .O(N__14802),
            .I(N__14796));
    CascadeMux I__2770 (
            .O(N__14799),
            .I(N__14793));
    CascadeMux I__2769 (
            .O(N__14796),
            .I(N__14790));
    CascadeBuf I__2768 (
            .O(N__14793),
            .I(N__14787));
    CascadeBuf I__2767 (
            .O(N__14790),
            .I(N__14784));
    CascadeMux I__2766 (
            .O(N__14787),
            .I(N__14781));
    CascadeMux I__2765 (
            .O(N__14784),
            .I(N__14778));
    CascadeBuf I__2764 (
            .O(N__14781),
            .I(N__14775));
    CascadeBuf I__2763 (
            .O(N__14778),
            .I(N__14772));
    CascadeMux I__2762 (
            .O(N__14775),
            .I(N__14769));
    CascadeMux I__2761 (
            .O(N__14772),
            .I(N__14766));
    CascadeBuf I__2760 (
            .O(N__14769),
            .I(N__14763));
    CascadeBuf I__2759 (
            .O(N__14766),
            .I(N__14760));
    CascadeMux I__2758 (
            .O(N__14763),
            .I(N__14757));
    CascadeMux I__2757 (
            .O(N__14760),
            .I(N__14754));
    CascadeBuf I__2756 (
            .O(N__14757),
            .I(N__14751));
    CascadeBuf I__2755 (
            .O(N__14754),
            .I(N__14748));
    CascadeMux I__2754 (
            .O(N__14751),
            .I(N__14745));
    CascadeMux I__2753 (
            .O(N__14748),
            .I(N__14742));
    CascadeBuf I__2752 (
            .O(N__14745),
            .I(N__14739));
    CascadeBuf I__2751 (
            .O(N__14742),
            .I(N__14736));
    CascadeMux I__2750 (
            .O(N__14739),
            .I(N__14733));
    CascadeMux I__2749 (
            .O(N__14736),
            .I(N__14730));
    CascadeBuf I__2748 (
            .O(N__14733),
            .I(N__14727));
    CascadeBuf I__2747 (
            .O(N__14730),
            .I(N__14724));
    CascadeMux I__2746 (
            .O(N__14727),
            .I(N__14721));
    CascadeMux I__2745 (
            .O(N__14724),
            .I(N__14718));
    CascadeBuf I__2744 (
            .O(N__14721),
            .I(N__14715));
    InMux I__2743 (
            .O(N__14718),
            .I(N__14711));
    CascadeMux I__2742 (
            .O(N__14715),
            .I(N__14708));
    CascadeMux I__2741 (
            .O(N__14714),
            .I(N__14705));
    LocalMux I__2740 (
            .O(N__14711),
            .I(N__14702));
    InMux I__2739 (
            .O(N__14708),
            .I(N__14699));
    InMux I__2738 (
            .O(N__14705),
            .I(N__14696));
    Span4Mux_h I__2737 (
            .O(N__14702),
            .I(N__14693));
    LocalMux I__2736 (
            .O(N__14699),
            .I(N__14690));
    LocalMux I__2735 (
            .O(N__14696),
            .I(N__14687));
    Span4Mux_h I__2734 (
            .O(N__14693),
            .I(N__14683));
    Span4Mux_h I__2733 (
            .O(N__14690),
            .I(N__14680));
    Span12Mux_v I__2732 (
            .O(N__14687),
            .I(N__14677));
    InMux I__2731 (
            .O(N__14686),
            .I(N__14674));
    Span4Mux_h I__2730 (
            .O(N__14683),
            .I(N__14669));
    Span4Mux_h I__2729 (
            .O(N__14680),
            .I(N__14669));
    Odrv12 I__2728 (
            .O(N__14677),
            .I(RX_ADDR_6));
    LocalMux I__2727 (
            .O(N__14674),
            .I(RX_ADDR_6));
    Odrv4 I__2726 (
            .O(N__14669),
            .I(RX_ADDR_6));
    InMux I__2725 (
            .O(N__14662),
            .I(N__14659));
    LocalMux I__2724 (
            .O(N__14659),
            .I(N__14656));
    Span12Mux_s2_v I__2723 (
            .O(N__14656),
            .I(N__14653));
    Span12Mux_v I__2722 (
            .O(N__14653),
            .I(N__14650));
    Odrv12 I__2721 (
            .O(N__14650),
            .I(\receive_module.n129 ));
    CascadeMux I__2720 (
            .O(N__14647),
            .I(N__14643));
    CascadeMux I__2719 (
            .O(N__14646),
            .I(N__14640));
    CascadeBuf I__2718 (
            .O(N__14643),
            .I(N__14637));
    CascadeBuf I__2717 (
            .O(N__14640),
            .I(N__14634));
    CascadeMux I__2716 (
            .O(N__14637),
            .I(N__14631));
    CascadeMux I__2715 (
            .O(N__14634),
            .I(N__14628));
    CascadeBuf I__2714 (
            .O(N__14631),
            .I(N__14625));
    CascadeBuf I__2713 (
            .O(N__14628),
            .I(N__14622));
    CascadeMux I__2712 (
            .O(N__14625),
            .I(N__14619));
    CascadeMux I__2711 (
            .O(N__14622),
            .I(N__14616));
    CascadeBuf I__2710 (
            .O(N__14619),
            .I(N__14613));
    CascadeBuf I__2709 (
            .O(N__14616),
            .I(N__14610));
    CascadeMux I__2708 (
            .O(N__14613),
            .I(N__14607));
    CascadeMux I__2707 (
            .O(N__14610),
            .I(N__14604));
    CascadeBuf I__2706 (
            .O(N__14607),
            .I(N__14601));
    CascadeBuf I__2705 (
            .O(N__14604),
            .I(N__14598));
    CascadeMux I__2704 (
            .O(N__14601),
            .I(N__14595));
    CascadeMux I__2703 (
            .O(N__14598),
            .I(N__14592));
    CascadeBuf I__2702 (
            .O(N__14595),
            .I(N__14589));
    CascadeBuf I__2701 (
            .O(N__14592),
            .I(N__14586));
    CascadeMux I__2700 (
            .O(N__14589),
            .I(N__14583));
    CascadeMux I__2699 (
            .O(N__14586),
            .I(N__14580));
    CascadeBuf I__2698 (
            .O(N__14583),
            .I(N__14577));
    CascadeBuf I__2697 (
            .O(N__14580),
            .I(N__14574));
    CascadeMux I__2696 (
            .O(N__14577),
            .I(N__14571));
    CascadeMux I__2695 (
            .O(N__14574),
            .I(N__14568));
    CascadeBuf I__2694 (
            .O(N__14571),
            .I(N__14565));
    CascadeBuf I__2693 (
            .O(N__14568),
            .I(N__14562));
    CascadeMux I__2692 (
            .O(N__14565),
            .I(N__14559));
    CascadeMux I__2691 (
            .O(N__14562),
            .I(N__14556));
    CascadeBuf I__2690 (
            .O(N__14559),
            .I(N__14553));
    CascadeBuf I__2689 (
            .O(N__14556),
            .I(N__14550));
    CascadeMux I__2688 (
            .O(N__14553),
            .I(N__14547));
    CascadeMux I__2687 (
            .O(N__14550),
            .I(N__14544));
    CascadeBuf I__2686 (
            .O(N__14547),
            .I(N__14541));
    CascadeBuf I__2685 (
            .O(N__14544),
            .I(N__14538));
    CascadeMux I__2684 (
            .O(N__14541),
            .I(N__14535));
    CascadeMux I__2683 (
            .O(N__14538),
            .I(N__14532));
    CascadeBuf I__2682 (
            .O(N__14535),
            .I(N__14529));
    CascadeBuf I__2681 (
            .O(N__14532),
            .I(N__14526));
    CascadeMux I__2680 (
            .O(N__14529),
            .I(N__14523));
    CascadeMux I__2679 (
            .O(N__14526),
            .I(N__14520));
    CascadeBuf I__2678 (
            .O(N__14523),
            .I(N__14517));
    CascadeBuf I__2677 (
            .O(N__14520),
            .I(N__14514));
    CascadeMux I__2676 (
            .O(N__14517),
            .I(N__14511));
    CascadeMux I__2675 (
            .O(N__14514),
            .I(N__14508));
    CascadeBuf I__2674 (
            .O(N__14511),
            .I(N__14505));
    CascadeBuf I__2673 (
            .O(N__14508),
            .I(N__14502));
    CascadeMux I__2672 (
            .O(N__14505),
            .I(N__14499));
    CascadeMux I__2671 (
            .O(N__14502),
            .I(N__14496));
    CascadeBuf I__2670 (
            .O(N__14499),
            .I(N__14493));
    CascadeBuf I__2669 (
            .O(N__14496),
            .I(N__14490));
    CascadeMux I__2668 (
            .O(N__14493),
            .I(N__14487));
    CascadeMux I__2667 (
            .O(N__14490),
            .I(N__14484));
    CascadeBuf I__2666 (
            .O(N__14487),
            .I(N__14481));
    CascadeBuf I__2665 (
            .O(N__14484),
            .I(N__14478));
    CascadeMux I__2664 (
            .O(N__14481),
            .I(N__14475));
    CascadeMux I__2663 (
            .O(N__14478),
            .I(N__14472));
    CascadeBuf I__2662 (
            .O(N__14475),
            .I(N__14469));
    CascadeBuf I__2661 (
            .O(N__14472),
            .I(N__14466));
    CascadeMux I__2660 (
            .O(N__14469),
            .I(N__14463));
    CascadeMux I__2659 (
            .O(N__14466),
            .I(N__14459));
    InMux I__2658 (
            .O(N__14463),
            .I(N__14456));
    InMux I__2657 (
            .O(N__14462),
            .I(N__14453));
    InMux I__2656 (
            .O(N__14459),
            .I(N__14450));
    LocalMux I__2655 (
            .O(N__14456),
            .I(N__14447));
    LocalMux I__2654 (
            .O(N__14453),
            .I(N__14443));
    LocalMux I__2653 (
            .O(N__14450),
            .I(N__14440));
    Span4Mux_s1_v I__2652 (
            .O(N__14447),
            .I(N__14437));
    CascadeMux I__2651 (
            .O(N__14446),
            .I(N__14434));
    Span12Mux_v I__2650 (
            .O(N__14443),
            .I(N__14431));
    Span4Mux_s1_v I__2649 (
            .O(N__14440),
            .I(N__14428));
    Span4Mux_h I__2648 (
            .O(N__14437),
            .I(N__14425));
    InMux I__2647 (
            .O(N__14434),
            .I(N__14422));
    Span12Mux_v I__2646 (
            .O(N__14431),
            .I(N__14419));
    Span4Mux_h I__2645 (
            .O(N__14428),
            .I(N__14414));
    Span4Mux_h I__2644 (
            .O(N__14425),
            .I(N__14414));
    LocalMux I__2643 (
            .O(N__14422),
            .I(RX_ADDR_7));
    Odrv12 I__2642 (
            .O(N__14419),
            .I(RX_ADDR_7));
    Odrv4 I__2641 (
            .O(N__14414),
            .I(RX_ADDR_7));
    InMux I__2640 (
            .O(N__14407),
            .I(N__14404));
    LocalMux I__2639 (
            .O(N__14404),
            .I(N__14401));
    Span12Mux_v I__2638 (
            .O(N__14401),
            .I(N__14398));
    Odrv12 I__2637 (
            .O(N__14398),
            .I(\receive_module.n128 ));
    CascadeMux I__2636 (
            .O(N__14395),
            .I(N__14392));
    CascadeBuf I__2635 (
            .O(N__14392),
            .I(N__14388));
    CascadeMux I__2634 (
            .O(N__14391),
            .I(N__14385));
    CascadeMux I__2633 (
            .O(N__14388),
            .I(N__14382));
    CascadeBuf I__2632 (
            .O(N__14385),
            .I(N__14379));
    CascadeBuf I__2631 (
            .O(N__14382),
            .I(N__14376));
    CascadeMux I__2630 (
            .O(N__14379),
            .I(N__14373));
    CascadeMux I__2629 (
            .O(N__14376),
            .I(N__14370));
    CascadeBuf I__2628 (
            .O(N__14373),
            .I(N__14367));
    CascadeBuf I__2627 (
            .O(N__14370),
            .I(N__14364));
    CascadeMux I__2626 (
            .O(N__14367),
            .I(N__14361));
    CascadeMux I__2625 (
            .O(N__14364),
            .I(N__14358));
    CascadeBuf I__2624 (
            .O(N__14361),
            .I(N__14355));
    CascadeBuf I__2623 (
            .O(N__14358),
            .I(N__14352));
    CascadeMux I__2622 (
            .O(N__14355),
            .I(N__14349));
    CascadeMux I__2621 (
            .O(N__14352),
            .I(N__14346));
    CascadeBuf I__2620 (
            .O(N__14349),
            .I(N__14343));
    CascadeBuf I__2619 (
            .O(N__14346),
            .I(N__14340));
    CascadeMux I__2618 (
            .O(N__14343),
            .I(N__14337));
    CascadeMux I__2617 (
            .O(N__14340),
            .I(N__14334));
    CascadeBuf I__2616 (
            .O(N__14337),
            .I(N__14331));
    CascadeBuf I__2615 (
            .O(N__14334),
            .I(N__14328));
    CascadeMux I__2614 (
            .O(N__14331),
            .I(N__14325));
    CascadeMux I__2613 (
            .O(N__14328),
            .I(N__14322));
    CascadeBuf I__2612 (
            .O(N__14325),
            .I(N__14319));
    CascadeBuf I__2611 (
            .O(N__14322),
            .I(N__14316));
    CascadeMux I__2610 (
            .O(N__14319),
            .I(N__14313));
    CascadeMux I__2609 (
            .O(N__14316),
            .I(N__14310));
    CascadeBuf I__2608 (
            .O(N__14313),
            .I(N__14307));
    CascadeBuf I__2607 (
            .O(N__14310),
            .I(N__14304));
    CascadeMux I__2606 (
            .O(N__14307),
            .I(N__14301));
    CascadeMux I__2605 (
            .O(N__14304),
            .I(N__14298));
    CascadeBuf I__2604 (
            .O(N__14301),
            .I(N__14295));
    CascadeBuf I__2603 (
            .O(N__14298),
            .I(N__14292));
    CascadeMux I__2602 (
            .O(N__14295),
            .I(N__14289));
    CascadeMux I__2601 (
            .O(N__14292),
            .I(N__14286));
    CascadeBuf I__2600 (
            .O(N__14289),
            .I(N__14283));
    CascadeBuf I__2599 (
            .O(N__14286),
            .I(N__14280));
    CascadeMux I__2598 (
            .O(N__14283),
            .I(N__14277));
    CascadeMux I__2597 (
            .O(N__14280),
            .I(N__14274));
    CascadeBuf I__2596 (
            .O(N__14277),
            .I(N__14271));
    CascadeBuf I__2595 (
            .O(N__14274),
            .I(N__14268));
    CascadeMux I__2594 (
            .O(N__14271),
            .I(N__14265));
    CascadeMux I__2593 (
            .O(N__14268),
            .I(N__14262));
    CascadeBuf I__2592 (
            .O(N__14265),
            .I(N__14259));
    CascadeBuf I__2591 (
            .O(N__14262),
            .I(N__14256));
    CascadeMux I__2590 (
            .O(N__14259),
            .I(N__14253));
    CascadeMux I__2589 (
            .O(N__14256),
            .I(N__14250));
    CascadeBuf I__2588 (
            .O(N__14253),
            .I(N__14247));
    CascadeBuf I__2587 (
            .O(N__14250),
            .I(N__14244));
    CascadeMux I__2586 (
            .O(N__14247),
            .I(N__14241));
    CascadeMux I__2585 (
            .O(N__14244),
            .I(N__14238));
    CascadeBuf I__2584 (
            .O(N__14241),
            .I(N__14235));
    CascadeBuf I__2583 (
            .O(N__14238),
            .I(N__14232));
    CascadeMux I__2582 (
            .O(N__14235),
            .I(N__14229));
    CascadeMux I__2581 (
            .O(N__14232),
            .I(N__14226));
    CascadeBuf I__2580 (
            .O(N__14229),
            .I(N__14223));
    CascadeBuf I__2579 (
            .O(N__14226),
            .I(N__14220));
    CascadeMux I__2578 (
            .O(N__14223),
            .I(N__14217));
    CascadeMux I__2577 (
            .O(N__14220),
            .I(N__14214));
    CascadeBuf I__2576 (
            .O(N__14217),
            .I(N__14211));
    InMux I__2575 (
            .O(N__14214),
            .I(N__14207));
    CascadeMux I__2574 (
            .O(N__14211),
            .I(N__14204));
    InMux I__2573 (
            .O(N__14210),
            .I(N__14201));
    LocalMux I__2572 (
            .O(N__14207),
            .I(N__14198));
    InMux I__2571 (
            .O(N__14204),
            .I(N__14195));
    LocalMux I__2570 (
            .O(N__14201),
            .I(N__14192));
    Span4Mux_s1_v I__2569 (
            .O(N__14198),
            .I(N__14189));
    LocalMux I__2568 (
            .O(N__14195),
            .I(N__14186));
    Span12Mux_h I__2567 (
            .O(N__14192),
            .I(N__14183));
    Span4Mux_h I__2566 (
            .O(N__14189),
            .I(N__14179));
    Span4Mux_s1_v I__2565 (
            .O(N__14186),
            .I(N__14176));
    Span12Mux_v I__2564 (
            .O(N__14183),
            .I(N__14173));
    InMux I__2563 (
            .O(N__14182),
            .I(N__14170));
    Span4Mux_h I__2562 (
            .O(N__14179),
            .I(N__14165));
    Span4Mux_h I__2561 (
            .O(N__14176),
            .I(N__14165));
    Odrv12 I__2560 (
            .O(N__14173),
            .I(RX_ADDR_8));
    LocalMux I__2559 (
            .O(N__14170),
            .I(RX_ADDR_8));
    Odrv4 I__2558 (
            .O(N__14165),
            .I(RX_ADDR_8));
    InMux I__2557 (
            .O(N__14158),
            .I(N__14155));
    LocalMux I__2556 (
            .O(N__14155),
            .I(N__14152));
    Span12Mux_s7_v I__2555 (
            .O(N__14152),
            .I(N__14149));
    Span12Mux_v I__2554 (
            .O(N__14149),
            .I(N__14146));
    Odrv12 I__2553 (
            .O(N__14146),
            .I(\receive_module.n127 ));
    CascadeMux I__2552 (
            .O(N__14143),
            .I(N__14140));
    CascadeBuf I__2551 (
            .O(N__14140),
            .I(N__14136));
    CascadeMux I__2550 (
            .O(N__14139),
            .I(N__14133));
    CascadeMux I__2549 (
            .O(N__14136),
            .I(N__14130));
    CascadeBuf I__2548 (
            .O(N__14133),
            .I(N__14127));
    CascadeBuf I__2547 (
            .O(N__14130),
            .I(N__14124));
    CascadeMux I__2546 (
            .O(N__14127),
            .I(N__14121));
    CascadeMux I__2545 (
            .O(N__14124),
            .I(N__14118));
    CascadeBuf I__2544 (
            .O(N__14121),
            .I(N__14115));
    CascadeBuf I__2543 (
            .O(N__14118),
            .I(N__14112));
    CascadeMux I__2542 (
            .O(N__14115),
            .I(N__14109));
    CascadeMux I__2541 (
            .O(N__14112),
            .I(N__14106));
    CascadeBuf I__2540 (
            .O(N__14109),
            .I(N__14103));
    CascadeBuf I__2539 (
            .O(N__14106),
            .I(N__14100));
    CascadeMux I__2538 (
            .O(N__14103),
            .I(N__14097));
    CascadeMux I__2537 (
            .O(N__14100),
            .I(N__14094));
    CascadeBuf I__2536 (
            .O(N__14097),
            .I(N__14091));
    CascadeBuf I__2535 (
            .O(N__14094),
            .I(N__14088));
    CascadeMux I__2534 (
            .O(N__14091),
            .I(N__14085));
    CascadeMux I__2533 (
            .O(N__14088),
            .I(N__14082));
    CascadeBuf I__2532 (
            .O(N__14085),
            .I(N__14079));
    CascadeBuf I__2531 (
            .O(N__14082),
            .I(N__14076));
    CascadeMux I__2530 (
            .O(N__14079),
            .I(N__14073));
    CascadeMux I__2529 (
            .O(N__14076),
            .I(N__14070));
    CascadeBuf I__2528 (
            .O(N__14073),
            .I(N__14067));
    CascadeBuf I__2527 (
            .O(N__14070),
            .I(N__14064));
    CascadeMux I__2526 (
            .O(N__14067),
            .I(N__14061));
    CascadeMux I__2525 (
            .O(N__14064),
            .I(N__14058));
    CascadeBuf I__2524 (
            .O(N__14061),
            .I(N__14055));
    CascadeBuf I__2523 (
            .O(N__14058),
            .I(N__14052));
    CascadeMux I__2522 (
            .O(N__14055),
            .I(N__14049));
    CascadeMux I__2521 (
            .O(N__14052),
            .I(N__14046));
    CascadeBuf I__2520 (
            .O(N__14049),
            .I(N__14043));
    CascadeBuf I__2519 (
            .O(N__14046),
            .I(N__14040));
    CascadeMux I__2518 (
            .O(N__14043),
            .I(N__14037));
    CascadeMux I__2517 (
            .O(N__14040),
            .I(N__14034));
    CascadeBuf I__2516 (
            .O(N__14037),
            .I(N__14031));
    CascadeBuf I__2515 (
            .O(N__14034),
            .I(N__14028));
    CascadeMux I__2514 (
            .O(N__14031),
            .I(N__14025));
    CascadeMux I__2513 (
            .O(N__14028),
            .I(N__14022));
    CascadeBuf I__2512 (
            .O(N__14025),
            .I(N__14019));
    CascadeBuf I__2511 (
            .O(N__14022),
            .I(N__14016));
    CascadeMux I__2510 (
            .O(N__14019),
            .I(N__14013));
    CascadeMux I__2509 (
            .O(N__14016),
            .I(N__14010));
    CascadeBuf I__2508 (
            .O(N__14013),
            .I(N__14007));
    CascadeBuf I__2507 (
            .O(N__14010),
            .I(N__14004));
    CascadeMux I__2506 (
            .O(N__14007),
            .I(N__14001));
    CascadeMux I__2505 (
            .O(N__14004),
            .I(N__13998));
    CascadeBuf I__2504 (
            .O(N__14001),
            .I(N__13995));
    CascadeBuf I__2503 (
            .O(N__13998),
            .I(N__13992));
    CascadeMux I__2502 (
            .O(N__13995),
            .I(N__13989));
    CascadeMux I__2501 (
            .O(N__13992),
            .I(N__13986));
    CascadeBuf I__2500 (
            .O(N__13989),
            .I(N__13983));
    CascadeBuf I__2499 (
            .O(N__13986),
            .I(N__13980));
    CascadeMux I__2498 (
            .O(N__13983),
            .I(N__13977));
    CascadeMux I__2497 (
            .O(N__13980),
            .I(N__13973));
    CascadeBuf I__2496 (
            .O(N__13977),
            .I(N__13970));
    InMux I__2495 (
            .O(N__13976),
            .I(N__13967));
    CascadeBuf I__2494 (
            .O(N__13973),
            .I(N__13964));
    CascadeMux I__2493 (
            .O(N__13970),
            .I(N__13961));
    LocalMux I__2492 (
            .O(N__13967),
            .I(N__13958));
    CascadeMux I__2491 (
            .O(N__13964),
            .I(N__13955));
    CascadeBuf I__2490 (
            .O(N__13961),
            .I(N__13952));
    Span4Mux_v I__2489 (
            .O(N__13958),
            .I(N__13949));
    InMux I__2488 (
            .O(N__13955),
            .I(N__13946));
    CascadeMux I__2487 (
            .O(N__13952),
            .I(N__13943));
    Span4Mux_v I__2486 (
            .O(N__13949),
            .I(N__13939));
    LocalMux I__2485 (
            .O(N__13946),
            .I(N__13936));
    InMux I__2484 (
            .O(N__13943),
            .I(N__13933));
    CascadeMux I__2483 (
            .O(N__13942),
            .I(N__13930));
    Span4Mux_v I__2482 (
            .O(N__13939),
            .I(N__13927));
    Span4Mux_s1_v I__2481 (
            .O(N__13936),
            .I(N__13924));
    LocalMux I__2480 (
            .O(N__13933),
            .I(N__13921));
    InMux I__2479 (
            .O(N__13930),
            .I(N__13918));
    Sp12to4 I__2478 (
            .O(N__13927),
            .I(N__13915));
    Span4Mux_h I__2477 (
            .O(N__13924),
            .I(N__13912));
    Span12Mux_s1_v I__2476 (
            .O(N__13921),
            .I(N__13909));
    LocalMux I__2475 (
            .O(N__13918),
            .I(RX_ADDR_9));
    Odrv12 I__2474 (
            .O(N__13915),
            .I(RX_ADDR_9));
    Odrv4 I__2473 (
            .O(N__13912),
            .I(RX_ADDR_9));
    Odrv12 I__2472 (
            .O(N__13909),
            .I(RX_ADDR_9));
    InMux I__2471 (
            .O(N__13900),
            .I(N__13897));
    LocalMux I__2470 (
            .O(N__13897),
            .I(\transmit_module.ADDR_Y_COMPONENT_9 ));
    InMux I__2469 (
            .O(N__13894),
            .I(N__13891));
    LocalMux I__2468 (
            .O(N__13891),
            .I(N__13888));
    Odrv4 I__2467 (
            .O(N__13888),
            .I(\transmit_module.ADDR_Y_COMPONENT_12 ));
    InMux I__2466 (
            .O(N__13885),
            .I(N__13882));
    LocalMux I__2465 (
            .O(N__13882),
            .I(N__13879));
    Odrv4 I__2464 (
            .O(N__13879),
            .I(\transmit_module.n120 ));
    InMux I__2463 (
            .O(N__13876),
            .I(N__13873));
    LocalMux I__2462 (
            .O(N__13873),
            .I(N__13870));
    Odrv4 I__2461 (
            .O(N__13870),
            .I(\transmit_module.n119 ));
    InMux I__2460 (
            .O(N__13867),
            .I(N__13864));
    LocalMux I__2459 (
            .O(N__13864),
            .I(N__13861));
    Span4Mux_h I__2458 (
            .O(N__13861),
            .I(N__13858));
    Odrv4 I__2457 (
            .O(N__13858),
            .I(\transmit_module.ADDR_Y_COMPONENT_11 ));
    InMux I__2456 (
            .O(N__13855),
            .I(N__13852));
    LocalMux I__2455 (
            .O(N__13852),
            .I(N__13849));
    Odrv4 I__2454 (
            .O(N__13849),
            .I(\transmit_module.n121 ));
    CEMux I__2453 (
            .O(N__13846),
            .I(N__13843));
    LocalMux I__2452 (
            .O(N__13843),
            .I(N__13839));
    CEMux I__2451 (
            .O(N__13842),
            .I(N__13836));
    Span4Mux_v I__2450 (
            .O(N__13839),
            .I(N__13833));
    LocalMux I__2449 (
            .O(N__13836),
            .I(N__13830));
    Span4Mux_h I__2448 (
            .O(N__13833),
            .I(N__13827));
    Odrv4 I__2447 (
            .O(N__13830),
            .I(\transmit_module.n2039 ));
    Odrv4 I__2446 (
            .O(N__13827),
            .I(\transmit_module.n2039 ));
    InMux I__2445 (
            .O(N__13822),
            .I(N__13819));
    LocalMux I__2444 (
            .O(N__13819),
            .I(N__13816));
    Odrv12 I__2443 (
            .O(N__13816),
            .I(\transmit_module.n130 ));
    InMux I__2442 (
            .O(N__13813),
            .I(N__13810));
    LocalMux I__2441 (
            .O(N__13810),
            .I(\line_buffer.n3755 ));
    InMux I__2440 (
            .O(N__13807),
            .I(N__13804));
    LocalMux I__2439 (
            .O(N__13804),
            .I(N__13801));
    Span4Mux_v I__2438 (
            .O(N__13801),
            .I(N__13798));
    Odrv4 I__2437 (
            .O(N__13798),
            .I(TX_DATA_0));
    InMux I__2436 (
            .O(N__13795),
            .I(N__13792));
    LocalMux I__2435 (
            .O(N__13792),
            .I(N__13789));
    Span12Mux_v I__2434 (
            .O(N__13789),
            .I(N__13786));
    Odrv12 I__2433 (
            .O(N__13786),
            .I(\receive_module.n134 ));
    CascadeMux I__2432 (
            .O(N__13783),
            .I(N__13779));
    CascadeMux I__2431 (
            .O(N__13782),
            .I(N__13776));
    CascadeBuf I__2430 (
            .O(N__13779),
            .I(N__13773));
    CascadeBuf I__2429 (
            .O(N__13776),
            .I(N__13770));
    CascadeMux I__2428 (
            .O(N__13773),
            .I(N__13767));
    CascadeMux I__2427 (
            .O(N__13770),
            .I(N__13764));
    CascadeBuf I__2426 (
            .O(N__13767),
            .I(N__13761));
    CascadeBuf I__2425 (
            .O(N__13764),
            .I(N__13758));
    CascadeMux I__2424 (
            .O(N__13761),
            .I(N__13755));
    CascadeMux I__2423 (
            .O(N__13758),
            .I(N__13752));
    CascadeBuf I__2422 (
            .O(N__13755),
            .I(N__13749));
    CascadeBuf I__2421 (
            .O(N__13752),
            .I(N__13746));
    CascadeMux I__2420 (
            .O(N__13749),
            .I(N__13743));
    CascadeMux I__2419 (
            .O(N__13746),
            .I(N__13740));
    CascadeBuf I__2418 (
            .O(N__13743),
            .I(N__13737));
    CascadeBuf I__2417 (
            .O(N__13740),
            .I(N__13734));
    CascadeMux I__2416 (
            .O(N__13737),
            .I(N__13731));
    CascadeMux I__2415 (
            .O(N__13734),
            .I(N__13728));
    CascadeBuf I__2414 (
            .O(N__13731),
            .I(N__13725));
    CascadeBuf I__2413 (
            .O(N__13728),
            .I(N__13722));
    CascadeMux I__2412 (
            .O(N__13725),
            .I(N__13719));
    CascadeMux I__2411 (
            .O(N__13722),
            .I(N__13716));
    CascadeBuf I__2410 (
            .O(N__13719),
            .I(N__13713));
    CascadeBuf I__2409 (
            .O(N__13716),
            .I(N__13710));
    CascadeMux I__2408 (
            .O(N__13713),
            .I(N__13707));
    CascadeMux I__2407 (
            .O(N__13710),
            .I(N__13704));
    CascadeBuf I__2406 (
            .O(N__13707),
            .I(N__13701));
    CascadeBuf I__2405 (
            .O(N__13704),
            .I(N__13698));
    CascadeMux I__2404 (
            .O(N__13701),
            .I(N__13695));
    CascadeMux I__2403 (
            .O(N__13698),
            .I(N__13692));
    CascadeBuf I__2402 (
            .O(N__13695),
            .I(N__13689));
    CascadeBuf I__2401 (
            .O(N__13692),
            .I(N__13686));
    CascadeMux I__2400 (
            .O(N__13689),
            .I(N__13683));
    CascadeMux I__2399 (
            .O(N__13686),
            .I(N__13680));
    CascadeBuf I__2398 (
            .O(N__13683),
            .I(N__13677));
    CascadeBuf I__2397 (
            .O(N__13680),
            .I(N__13674));
    CascadeMux I__2396 (
            .O(N__13677),
            .I(N__13671));
    CascadeMux I__2395 (
            .O(N__13674),
            .I(N__13668));
    CascadeBuf I__2394 (
            .O(N__13671),
            .I(N__13665));
    CascadeBuf I__2393 (
            .O(N__13668),
            .I(N__13662));
    CascadeMux I__2392 (
            .O(N__13665),
            .I(N__13659));
    CascadeMux I__2391 (
            .O(N__13662),
            .I(N__13656));
    CascadeBuf I__2390 (
            .O(N__13659),
            .I(N__13653));
    CascadeBuf I__2389 (
            .O(N__13656),
            .I(N__13650));
    CascadeMux I__2388 (
            .O(N__13653),
            .I(N__13647));
    CascadeMux I__2387 (
            .O(N__13650),
            .I(N__13644));
    CascadeBuf I__2386 (
            .O(N__13647),
            .I(N__13641));
    CascadeBuf I__2385 (
            .O(N__13644),
            .I(N__13638));
    CascadeMux I__2384 (
            .O(N__13641),
            .I(N__13635));
    CascadeMux I__2383 (
            .O(N__13638),
            .I(N__13632));
    CascadeBuf I__2382 (
            .O(N__13635),
            .I(N__13629));
    CascadeBuf I__2381 (
            .O(N__13632),
            .I(N__13626));
    CascadeMux I__2380 (
            .O(N__13629),
            .I(N__13623));
    CascadeMux I__2379 (
            .O(N__13626),
            .I(N__13620));
    CascadeBuf I__2378 (
            .O(N__13623),
            .I(N__13617));
    CascadeBuf I__2377 (
            .O(N__13620),
            .I(N__13614));
    CascadeMux I__2376 (
            .O(N__13617),
            .I(N__13611));
    CascadeMux I__2375 (
            .O(N__13614),
            .I(N__13608));
    CascadeBuf I__2374 (
            .O(N__13611),
            .I(N__13605));
    CascadeBuf I__2373 (
            .O(N__13608),
            .I(N__13602));
    CascadeMux I__2372 (
            .O(N__13605),
            .I(N__13599));
    CascadeMux I__2371 (
            .O(N__13602),
            .I(N__13596));
    InMux I__2370 (
            .O(N__13599),
            .I(N__13593));
    InMux I__2369 (
            .O(N__13596),
            .I(N__13590));
    LocalMux I__2368 (
            .O(N__13593),
            .I(N__13586));
    LocalMux I__2367 (
            .O(N__13590),
            .I(N__13583));
    InMux I__2366 (
            .O(N__13589),
            .I(N__13580));
    Span4Mux_h I__2365 (
            .O(N__13586),
            .I(N__13577));
    Span4Mux_h I__2364 (
            .O(N__13583),
            .I(N__13574));
    LocalMux I__2363 (
            .O(N__13580),
            .I(N__13571));
    Sp12to4 I__2362 (
            .O(N__13577),
            .I(N__13567));
    Sp12to4 I__2361 (
            .O(N__13574),
            .I(N__13564));
    Span12Mux_v I__2360 (
            .O(N__13571),
            .I(N__13561));
    InMux I__2359 (
            .O(N__13570),
            .I(N__13558));
    Span12Mux_v I__2358 (
            .O(N__13567),
            .I(N__13553));
    Span12Mux_v I__2357 (
            .O(N__13564),
            .I(N__13553));
    Odrv12 I__2356 (
            .O(N__13561),
            .I(RX_ADDR_2));
    LocalMux I__2355 (
            .O(N__13558),
            .I(RX_ADDR_2));
    Odrv12 I__2354 (
            .O(N__13553),
            .I(RX_ADDR_2));
    CascadeMux I__2353 (
            .O(N__13546),
            .I(N__13540));
    InMux I__2352 (
            .O(N__13545),
            .I(N__13537));
    CascadeMux I__2351 (
            .O(N__13544),
            .I(N__13534));
    InMux I__2350 (
            .O(N__13543),
            .I(N__13531));
    InMux I__2349 (
            .O(N__13540),
            .I(N__13528));
    LocalMux I__2348 (
            .O(N__13537),
            .I(N__13525));
    InMux I__2347 (
            .O(N__13534),
            .I(N__13522));
    LocalMux I__2346 (
            .O(N__13531),
            .I(\transmit_module.TX_ADDR_7 ));
    LocalMux I__2345 (
            .O(N__13528),
            .I(\transmit_module.TX_ADDR_7 ));
    Odrv4 I__2344 (
            .O(N__13525),
            .I(\transmit_module.TX_ADDR_7 ));
    LocalMux I__2343 (
            .O(N__13522),
            .I(\transmit_module.TX_ADDR_7 ));
    InMux I__2342 (
            .O(N__13513),
            .I(N__13510));
    LocalMux I__2341 (
            .O(N__13510),
            .I(\transmit_module.n125 ));
    InMux I__2340 (
            .O(N__13507),
            .I(\transmit_module.n3264 ));
    InMux I__2339 (
            .O(N__13504),
            .I(bfn_15_14_0_));
    InMux I__2338 (
            .O(N__13501),
            .I(\transmit_module.n3266 ));
    InMux I__2337 (
            .O(N__13498),
            .I(N__13492));
    InMux I__2336 (
            .O(N__13497),
            .I(N__13487));
    InMux I__2335 (
            .O(N__13496),
            .I(N__13487));
    InMux I__2334 (
            .O(N__13495),
            .I(N__13484));
    LocalMux I__2333 (
            .O(N__13492),
            .I(\transmit_module.TX_ADDR_10 ));
    LocalMux I__2332 (
            .O(N__13487),
            .I(\transmit_module.TX_ADDR_10 ));
    LocalMux I__2331 (
            .O(N__13484),
            .I(\transmit_module.TX_ADDR_10 ));
    InMux I__2330 (
            .O(N__13477),
            .I(N__13474));
    LocalMux I__2329 (
            .O(N__13474),
            .I(\transmit_module.n122 ));
    InMux I__2328 (
            .O(N__13471),
            .I(\transmit_module.n3267 ));
    InMux I__2327 (
            .O(N__13468),
            .I(\transmit_module.n3268 ));
    InMux I__2326 (
            .O(N__13465),
            .I(\transmit_module.n3269 ));
    InMux I__2325 (
            .O(N__13462),
            .I(\transmit_module.n3270 ));
    InMux I__2324 (
            .O(N__13459),
            .I(\receive_module.n3257 ));
    InMux I__2323 (
            .O(N__13456),
            .I(N__13451));
    InMux I__2322 (
            .O(N__13455),
            .I(N__13448));
    InMux I__2321 (
            .O(N__13454),
            .I(N__13445));
    LocalMux I__2320 (
            .O(N__13451),
            .I(N__13440));
    LocalMux I__2319 (
            .O(N__13448),
            .I(N__13440));
    LocalMux I__2318 (
            .O(N__13445),
            .I(N__13434));
    Span4Mux_v I__2317 (
            .O(N__13440),
            .I(N__13434));
    InMux I__2316 (
            .O(N__13439),
            .I(N__13431));
    Odrv4 I__2315 (
            .O(N__13434),
            .I(\transmit_module.TX_ADDR_0 ));
    LocalMux I__2314 (
            .O(N__13431),
            .I(\transmit_module.TX_ADDR_0 ));
    InMux I__2313 (
            .O(N__13426),
            .I(N__13423));
    LocalMux I__2312 (
            .O(N__13423),
            .I(N__13419));
    CascadeMux I__2311 (
            .O(N__13422),
            .I(N__13416));
    Span4Mux_v I__2310 (
            .O(N__13419),
            .I(N__13413));
    InMux I__2309 (
            .O(N__13416),
            .I(N__13410));
    Span4Mux_h I__2308 (
            .O(N__13413),
            .I(N__13407));
    LocalMux I__2307 (
            .O(N__13410),
            .I(N__13404));
    Odrv4 I__2306 (
            .O(N__13407),
            .I(\transmit_module.X_DELTA_PATTERN_0 ));
    Odrv4 I__2305 (
            .O(N__13404),
            .I(\transmit_module.X_DELTA_PATTERN_0 ));
    InMux I__2304 (
            .O(N__13399),
            .I(N__13396));
    LocalMux I__2303 (
            .O(N__13396),
            .I(N__13393));
    Odrv4 I__2302 (
            .O(N__13393),
            .I(\transmit_module.n132 ));
    InMux I__2301 (
            .O(N__13390),
            .I(N__13386));
    CascadeMux I__2300 (
            .O(N__13389),
            .I(N__13381));
    LocalMux I__2299 (
            .O(N__13386),
            .I(N__13378));
    InMux I__2298 (
            .O(N__13385),
            .I(N__13373));
    InMux I__2297 (
            .O(N__13384),
            .I(N__13373));
    InMux I__2296 (
            .O(N__13381),
            .I(N__13370));
    Odrv4 I__2295 (
            .O(N__13378),
            .I(\transmit_module.TX_ADDR_1 ));
    LocalMux I__2294 (
            .O(N__13373),
            .I(\transmit_module.TX_ADDR_1 ));
    LocalMux I__2293 (
            .O(N__13370),
            .I(\transmit_module.TX_ADDR_1 ));
    CascadeMux I__2292 (
            .O(N__13363),
            .I(N__13360));
    InMux I__2291 (
            .O(N__13360),
            .I(N__13357));
    LocalMux I__2290 (
            .O(N__13357),
            .I(N__13354));
    Odrv4 I__2289 (
            .O(N__13354),
            .I(\transmit_module.n131 ));
    InMux I__2288 (
            .O(N__13351),
            .I(\transmit_module.n3258 ));
    InMux I__2287 (
            .O(N__13348),
            .I(\transmit_module.n3259 ));
    InMux I__2286 (
            .O(N__13345),
            .I(\transmit_module.n3260 ));
    InMux I__2285 (
            .O(N__13342),
            .I(N__13339));
    LocalMux I__2284 (
            .O(N__13339),
            .I(N__13333));
    InMux I__2283 (
            .O(N__13338),
            .I(N__13330));
    InMux I__2282 (
            .O(N__13337),
            .I(N__13327));
    InMux I__2281 (
            .O(N__13336),
            .I(N__13324));
    Odrv4 I__2280 (
            .O(N__13333),
            .I(\transmit_module.TX_ADDR_4 ));
    LocalMux I__2279 (
            .O(N__13330),
            .I(\transmit_module.TX_ADDR_4 ));
    LocalMux I__2278 (
            .O(N__13327),
            .I(\transmit_module.TX_ADDR_4 ));
    LocalMux I__2277 (
            .O(N__13324),
            .I(\transmit_module.TX_ADDR_4 ));
    InMux I__2276 (
            .O(N__13315),
            .I(N__13312));
    LocalMux I__2275 (
            .O(N__13312),
            .I(\transmit_module.n128 ));
    InMux I__2274 (
            .O(N__13309),
            .I(\transmit_module.n3261 ));
    InMux I__2273 (
            .O(N__13306),
            .I(N__13301));
    InMux I__2272 (
            .O(N__13305),
            .I(N__13298));
    CascadeMux I__2271 (
            .O(N__13304),
            .I(N__13294));
    LocalMux I__2270 (
            .O(N__13301),
            .I(N__13289));
    LocalMux I__2269 (
            .O(N__13298),
            .I(N__13289));
    InMux I__2268 (
            .O(N__13297),
            .I(N__13286));
    InMux I__2267 (
            .O(N__13294),
            .I(N__13283));
    Odrv4 I__2266 (
            .O(N__13289),
            .I(\transmit_module.TX_ADDR_5 ));
    LocalMux I__2265 (
            .O(N__13286),
            .I(\transmit_module.TX_ADDR_5 ));
    LocalMux I__2264 (
            .O(N__13283),
            .I(\transmit_module.TX_ADDR_5 ));
    InMux I__2263 (
            .O(N__13276),
            .I(N__13273));
    LocalMux I__2262 (
            .O(N__13273),
            .I(\transmit_module.n127 ));
    InMux I__2261 (
            .O(N__13270),
            .I(\transmit_module.n3262 ));
    InMux I__2260 (
            .O(N__13267),
            .I(N__13262));
    InMux I__2259 (
            .O(N__13266),
            .I(N__13259));
    CascadeMux I__2258 (
            .O(N__13265),
            .I(N__13255));
    LocalMux I__2257 (
            .O(N__13262),
            .I(N__13252));
    LocalMux I__2256 (
            .O(N__13259),
            .I(N__13249));
    InMux I__2255 (
            .O(N__13258),
            .I(N__13246));
    InMux I__2254 (
            .O(N__13255),
            .I(N__13243));
    Odrv12 I__2253 (
            .O(N__13252),
            .I(\transmit_module.TX_ADDR_6 ));
    Odrv4 I__2252 (
            .O(N__13249),
            .I(\transmit_module.TX_ADDR_6 ));
    LocalMux I__2251 (
            .O(N__13246),
            .I(\transmit_module.TX_ADDR_6 ));
    LocalMux I__2250 (
            .O(N__13243),
            .I(\transmit_module.TX_ADDR_6 ));
    InMux I__2249 (
            .O(N__13234),
            .I(N__13231));
    LocalMux I__2248 (
            .O(N__13231),
            .I(\transmit_module.n126 ));
    InMux I__2247 (
            .O(N__13228),
            .I(\transmit_module.n3263 ));
    InMux I__2246 (
            .O(N__13225),
            .I(\receive_module.n3248 ));
    InMux I__2245 (
            .O(N__13222),
            .I(\receive_module.n3249 ));
    InMux I__2244 (
            .O(N__13219),
            .I(\receive_module.n3250 ));
    InMux I__2243 (
            .O(N__13216),
            .I(\receive_module.n3251 ));
    InMux I__2242 (
            .O(N__13213),
            .I(bfn_15_12_0_));
    InMux I__2241 (
            .O(N__13210),
            .I(\receive_module.n3253 ));
    InMux I__2240 (
            .O(N__13207),
            .I(\receive_module.n3254 ));
    InMux I__2239 (
            .O(N__13204),
            .I(\receive_module.n3255 ));
    InMux I__2238 (
            .O(N__13201),
            .I(\receive_module.n3256 ));
    InMux I__2237 (
            .O(N__13198),
            .I(N__13195));
    LocalMux I__2236 (
            .O(N__13195),
            .I(N__13192));
    Span4Mux_h I__2235 (
            .O(N__13192),
            .I(N__13189));
    Span4Mux_h I__2234 (
            .O(N__13189),
            .I(N__13186));
    Odrv4 I__2233 (
            .O(N__13186),
            .I(\line_buffer.n543 ));
    InMux I__2232 (
            .O(N__13183),
            .I(N__13180));
    LocalMux I__2231 (
            .O(N__13180),
            .I(N__13177));
    Span4Mux_h I__2230 (
            .O(N__13177),
            .I(N__13174));
    Span4Mux_h I__2229 (
            .O(N__13174),
            .I(N__13171));
    Span4Mux_h I__2228 (
            .O(N__13171),
            .I(N__13168));
    Odrv4 I__2227 (
            .O(N__13168),
            .I(\line_buffer.n535 ));
    InMux I__2226 (
            .O(N__13165),
            .I(N__13161));
    InMux I__2225 (
            .O(N__13164),
            .I(N__13156));
    LocalMux I__2224 (
            .O(N__13161),
            .I(N__13153));
    InMux I__2223 (
            .O(N__13160),
            .I(N__13148));
    InMux I__2222 (
            .O(N__13159),
            .I(N__13148));
    LocalMux I__2221 (
            .O(N__13156),
            .I(\receive_module.rx_counter.Y_7 ));
    Odrv4 I__2220 (
            .O(N__13153),
            .I(\receive_module.rx_counter.Y_7 ));
    LocalMux I__2219 (
            .O(N__13148),
            .I(\receive_module.rx_counter.Y_7 ));
    InMux I__2218 (
            .O(N__13141),
            .I(N__13137));
    InMux I__2217 (
            .O(N__13140),
            .I(N__13134));
    LocalMux I__2216 (
            .O(N__13137),
            .I(\receive_module.rx_counter.n3791 ));
    LocalMux I__2215 (
            .O(N__13134),
            .I(\receive_module.rx_counter.n3791 ));
    CascadeMux I__2214 (
            .O(N__13129),
            .I(N__13126));
    InMux I__2213 (
            .O(N__13126),
            .I(N__13123));
    LocalMux I__2212 (
            .O(N__13123),
            .I(N__13117));
    InMux I__2211 (
            .O(N__13122),
            .I(N__13114));
    InMux I__2210 (
            .O(N__13121),
            .I(N__13109));
    InMux I__2209 (
            .O(N__13120),
            .I(N__13109));
    Odrv4 I__2208 (
            .O(N__13117),
            .I(\receive_module.rx_counter.Y_4 ));
    LocalMux I__2207 (
            .O(N__13114),
            .I(\receive_module.rx_counter.Y_4 ));
    LocalMux I__2206 (
            .O(N__13109),
            .I(\receive_module.rx_counter.Y_4 ));
    InMux I__2205 (
            .O(N__13102),
            .I(N__13099));
    LocalMux I__2204 (
            .O(N__13099),
            .I(\receive_module.rx_counter.n3551 ));
    CEMux I__2203 (
            .O(N__13096),
            .I(N__13093));
    LocalMux I__2202 (
            .O(N__13093),
            .I(N__13089));
    CEMux I__2201 (
            .O(N__13092),
            .I(N__13086));
    Span4Mux_h I__2200 (
            .O(N__13089),
            .I(N__13083));
    LocalMux I__2199 (
            .O(N__13086),
            .I(N__13080));
    Odrv4 I__2198 (
            .O(N__13083),
            .I(\receive_module.rx_counter.n2045 ));
    Odrv12 I__2197 (
            .O(N__13080),
            .I(\receive_module.rx_counter.n2045 ));
    InMux I__2196 (
            .O(N__13075),
            .I(N__13072));
    LocalMux I__2195 (
            .O(N__13072),
            .I(\receive_module.rx_counter.old_HS ));
    InMux I__2194 (
            .O(N__13069),
            .I(bfn_15_11_0_));
    InMux I__2193 (
            .O(N__13066),
            .I(\receive_module.n3245 ));
    InMux I__2192 (
            .O(N__13063),
            .I(\receive_module.n3246 ));
    InMux I__2191 (
            .O(N__13060),
            .I(\receive_module.n3247 ));
    InMux I__2190 (
            .O(N__13057),
            .I(N__13054));
    LocalMux I__2189 (
            .O(N__13054),
            .I(N__13050));
    InMux I__2188 (
            .O(N__13053),
            .I(N__13047));
    Span4Mux_v I__2187 (
            .O(N__13050),
            .I(N__13044));
    LocalMux I__2186 (
            .O(N__13047),
            .I(N__13041));
    Span4Mux_v I__2185 (
            .O(N__13044),
            .I(N__13038));
    Odrv4 I__2184 (
            .O(N__13041),
            .I(\transmit_module.n110 ));
    Odrv4 I__2183 (
            .O(N__13038),
            .I(\transmit_module.n110 ));
    InMux I__2182 (
            .O(N__13033),
            .I(N__13030));
    LocalMux I__2181 (
            .O(N__13030),
            .I(N__13027));
    Span12Mux_v I__2180 (
            .O(N__13027),
            .I(N__13024));
    Odrv12 I__2179 (
            .O(N__13024),
            .I(\transmit_module.n141 ));
    CascadeMux I__2178 (
            .O(N__13021),
            .I(N__13018));
    CascadeBuf I__2177 (
            .O(N__13018),
            .I(N__13015));
    CascadeMux I__2176 (
            .O(N__13015),
            .I(N__13011));
    CascadeMux I__2175 (
            .O(N__13014),
            .I(N__13008));
    CascadeBuf I__2174 (
            .O(N__13011),
            .I(N__13005));
    CascadeBuf I__2173 (
            .O(N__13008),
            .I(N__13002));
    CascadeMux I__2172 (
            .O(N__13005),
            .I(N__12999));
    CascadeMux I__2171 (
            .O(N__13002),
            .I(N__12996));
    CascadeBuf I__2170 (
            .O(N__12999),
            .I(N__12993));
    CascadeBuf I__2169 (
            .O(N__12996),
            .I(N__12990));
    CascadeMux I__2168 (
            .O(N__12993),
            .I(N__12987));
    CascadeMux I__2167 (
            .O(N__12990),
            .I(N__12984));
    CascadeBuf I__2166 (
            .O(N__12987),
            .I(N__12981));
    CascadeBuf I__2165 (
            .O(N__12984),
            .I(N__12978));
    CascadeMux I__2164 (
            .O(N__12981),
            .I(N__12975));
    CascadeMux I__2163 (
            .O(N__12978),
            .I(N__12972));
    CascadeBuf I__2162 (
            .O(N__12975),
            .I(N__12969));
    CascadeBuf I__2161 (
            .O(N__12972),
            .I(N__12966));
    CascadeMux I__2160 (
            .O(N__12969),
            .I(N__12963));
    CascadeMux I__2159 (
            .O(N__12966),
            .I(N__12960));
    CascadeBuf I__2158 (
            .O(N__12963),
            .I(N__12957));
    CascadeBuf I__2157 (
            .O(N__12960),
            .I(N__12954));
    CascadeMux I__2156 (
            .O(N__12957),
            .I(N__12951));
    CascadeMux I__2155 (
            .O(N__12954),
            .I(N__12948));
    CascadeBuf I__2154 (
            .O(N__12951),
            .I(N__12945));
    CascadeBuf I__2153 (
            .O(N__12948),
            .I(N__12942));
    CascadeMux I__2152 (
            .O(N__12945),
            .I(N__12939));
    CascadeMux I__2151 (
            .O(N__12942),
            .I(N__12936));
    CascadeBuf I__2150 (
            .O(N__12939),
            .I(N__12933));
    CascadeBuf I__2149 (
            .O(N__12936),
            .I(N__12930));
    CascadeMux I__2148 (
            .O(N__12933),
            .I(N__12927));
    CascadeMux I__2147 (
            .O(N__12930),
            .I(N__12924));
    CascadeBuf I__2146 (
            .O(N__12927),
            .I(N__12921));
    CascadeBuf I__2145 (
            .O(N__12924),
            .I(N__12918));
    CascadeMux I__2144 (
            .O(N__12921),
            .I(N__12915));
    CascadeMux I__2143 (
            .O(N__12918),
            .I(N__12912));
    CascadeBuf I__2142 (
            .O(N__12915),
            .I(N__12909));
    CascadeBuf I__2141 (
            .O(N__12912),
            .I(N__12906));
    CascadeMux I__2140 (
            .O(N__12909),
            .I(N__12903));
    CascadeMux I__2139 (
            .O(N__12906),
            .I(N__12900));
    CascadeBuf I__2138 (
            .O(N__12903),
            .I(N__12897));
    CascadeBuf I__2137 (
            .O(N__12900),
            .I(N__12894));
    CascadeMux I__2136 (
            .O(N__12897),
            .I(N__12891));
    CascadeMux I__2135 (
            .O(N__12894),
            .I(N__12888));
    CascadeBuf I__2134 (
            .O(N__12891),
            .I(N__12885));
    CascadeBuf I__2133 (
            .O(N__12888),
            .I(N__12882));
    CascadeMux I__2132 (
            .O(N__12885),
            .I(N__12879));
    CascadeMux I__2131 (
            .O(N__12882),
            .I(N__12876));
    CascadeBuf I__2130 (
            .O(N__12879),
            .I(N__12873));
    CascadeBuf I__2129 (
            .O(N__12876),
            .I(N__12870));
    CascadeMux I__2128 (
            .O(N__12873),
            .I(N__12867));
    CascadeMux I__2127 (
            .O(N__12870),
            .I(N__12864));
    CascadeBuf I__2126 (
            .O(N__12867),
            .I(N__12861));
    CascadeBuf I__2125 (
            .O(N__12864),
            .I(N__12858));
    CascadeMux I__2124 (
            .O(N__12861),
            .I(N__12855));
    CascadeMux I__2123 (
            .O(N__12858),
            .I(N__12852));
    CascadeBuf I__2122 (
            .O(N__12855),
            .I(N__12849));
    CascadeBuf I__2121 (
            .O(N__12852),
            .I(N__12846));
    CascadeMux I__2120 (
            .O(N__12849),
            .I(N__12843));
    CascadeMux I__2119 (
            .O(N__12846),
            .I(N__12840));
    InMux I__2118 (
            .O(N__12843),
            .I(N__12837));
    CascadeBuf I__2117 (
            .O(N__12840),
            .I(N__12834));
    LocalMux I__2116 (
            .O(N__12837),
            .I(N__12831));
    CascadeMux I__2115 (
            .O(N__12834),
            .I(N__12828));
    Span4Mux_h I__2114 (
            .O(N__12831),
            .I(N__12825));
    InMux I__2113 (
            .O(N__12828),
            .I(N__12822));
    Span4Mux_h I__2112 (
            .O(N__12825),
            .I(N__12819));
    LocalMux I__2111 (
            .O(N__12822),
            .I(N__12816));
    Span4Mux_h I__2110 (
            .O(N__12819),
            .I(N__12813));
    Span12Mux_s4_v I__2109 (
            .O(N__12816),
            .I(N__12810));
    Odrv4 I__2108 (
            .O(N__12813),
            .I(n22));
    Odrv12 I__2107 (
            .O(N__12810),
            .I(n22));
    InMux I__2106 (
            .O(N__12805),
            .I(N__12802));
    LocalMux I__2105 (
            .O(N__12802),
            .I(N__12798));
    InMux I__2104 (
            .O(N__12801),
            .I(N__12795));
    Span12Mux_s4_v I__2103 (
            .O(N__12798),
            .I(N__12792));
    LocalMux I__2102 (
            .O(N__12795),
            .I(N__12789));
    Span12Mux_v I__2101 (
            .O(N__12792),
            .I(N__12786));
    Odrv4 I__2100 (
            .O(N__12789),
            .I(\transmit_module.n109 ));
    Odrv12 I__2099 (
            .O(N__12786),
            .I(\transmit_module.n109 ));
    InMux I__2098 (
            .O(N__12781),
            .I(N__12778));
    LocalMux I__2097 (
            .O(N__12778),
            .I(N__12774));
    InMux I__2096 (
            .O(N__12777),
            .I(N__12771));
    Span12Mux_s11_v I__2095 (
            .O(N__12774),
            .I(N__12768));
    LocalMux I__2094 (
            .O(N__12771),
            .I(\transmit_module.n140 ));
    Odrv12 I__2093 (
            .O(N__12768),
            .I(\transmit_module.n140 ));
    CascadeMux I__2092 (
            .O(N__12763),
            .I(N__12759));
    CascadeMux I__2091 (
            .O(N__12762),
            .I(N__12756));
    CascadeBuf I__2090 (
            .O(N__12759),
            .I(N__12753));
    CascadeBuf I__2089 (
            .O(N__12756),
            .I(N__12750));
    CascadeMux I__2088 (
            .O(N__12753),
            .I(N__12747));
    CascadeMux I__2087 (
            .O(N__12750),
            .I(N__12744));
    CascadeBuf I__2086 (
            .O(N__12747),
            .I(N__12741));
    CascadeBuf I__2085 (
            .O(N__12744),
            .I(N__12738));
    CascadeMux I__2084 (
            .O(N__12741),
            .I(N__12735));
    CascadeMux I__2083 (
            .O(N__12738),
            .I(N__12732));
    CascadeBuf I__2082 (
            .O(N__12735),
            .I(N__12729));
    CascadeBuf I__2081 (
            .O(N__12732),
            .I(N__12726));
    CascadeMux I__2080 (
            .O(N__12729),
            .I(N__12723));
    CascadeMux I__2079 (
            .O(N__12726),
            .I(N__12720));
    CascadeBuf I__2078 (
            .O(N__12723),
            .I(N__12717));
    CascadeBuf I__2077 (
            .O(N__12720),
            .I(N__12714));
    CascadeMux I__2076 (
            .O(N__12717),
            .I(N__12711));
    CascadeMux I__2075 (
            .O(N__12714),
            .I(N__12708));
    CascadeBuf I__2074 (
            .O(N__12711),
            .I(N__12705));
    CascadeBuf I__2073 (
            .O(N__12708),
            .I(N__12702));
    CascadeMux I__2072 (
            .O(N__12705),
            .I(N__12699));
    CascadeMux I__2071 (
            .O(N__12702),
            .I(N__12696));
    CascadeBuf I__2070 (
            .O(N__12699),
            .I(N__12693));
    CascadeBuf I__2069 (
            .O(N__12696),
            .I(N__12690));
    CascadeMux I__2068 (
            .O(N__12693),
            .I(N__12687));
    CascadeMux I__2067 (
            .O(N__12690),
            .I(N__12684));
    CascadeBuf I__2066 (
            .O(N__12687),
            .I(N__12681));
    CascadeBuf I__2065 (
            .O(N__12684),
            .I(N__12678));
    CascadeMux I__2064 (
            .O(N__12681),
            .I(N__12675));
    CascadeMux I__2063 (
            .O(N__12678),
            .I(N__12672));
    CascadeBuf I__2062 (
            .O(N__12675),
            .I(N__12669));
    CascadeBuf I__2061 (
            .O(N__12672),
            .I(N__12666));
    CascadeMux I__2060 (
            .O(N__12669),
            .I(N__12663));
    CascadeMux I__2059 (
            .O(N__12666),
            .I(N__12660));
    CascadeBuf I__2058 (
            .O(N__12663),
            .I(N__12657));
    CascadeBuf I__2057 (
            .O(N__12660),
            .I(N__12654));
    CascadeMux I__2056 (
            .O(N__12657),
            .I(N__12651));
    CascadeMux I__2055 (
            .O(N__12654),
            .I(N__12648));
    CascadeBuf I__2054 (
            .O(N__12651),
            .I(N__12645));
    CascadeBuf I__2053 (
            .O(N__12648),
            .I(N__12642));
    CascadeMux I__2052 (
            .O(N__12645),
            .I(N__12639));
    CascadeMux I__2051 (
            .O(N__12642),
            .I(N__12636));
    CascadeBuf I__2050 (
            .O(N__12639),
            .I(N__12633));
    CascadeBuf I__2049 (
            .O(N__12636),
            .I(N__12630));
    CascadeMux I__2048 (
            .O(N__12633),
            .I(N__12627));
    CascadeMux I__2047 (
            .O(N__12630),
            .I(N__12624));
    CascadeBuf I__2046 (
            .O(N__12627),
            .I(N__12621));
    CascadeBuf I__2045 (
            .O(N__12624),
            .I(N__12618));
    CascadeMux I__2044 (
            .O(N__12621),
            .I(N__12615));
    CascadeMux I__2043 (
            .O(N__12618),
            .I(N__12612));
    CascadeBuf I__2042 (
            .O(N__12615),
            .I(N__12609));
    CascadeBuf I__2041 (
            .O(N__12612),
            .I(N__12606));
    CascadeMux I__2040 (
            .O(N__12609),
            .I(N__12603));
    CascadeMux I__2039 (
            .O(N__12606),
            .I(N__12600));
    CascadeBuf I__2038 (
            .O(N__12603),
            .I(N__12597));
    CascadeBuf I__2037 (
            .O(N__12600),
            .I(N__12594));
    CascadeMux I__2036 (
            .O(N__12597),
            .I(N__12591));
    CascadeMux I__2035 (
            .O(N__12594),
            .I(N__12588));
    CascadeBuf I__2034 (
            .O(N__12591),
            .I(N__12585));
    CascadeBuf I__2033 (
            .O(N__12588),
            .I(N__12582));
    CascadeMux I__2032 (
            .O(N__12585),
            .I(N__12579));
    CascadeMux I__2031 (
            .O(N__12582),
            .I(N__12576));
    InMux I__2030 (
            .O(N__12579),
            .I(N__12573));
    InMux I__2029 (
            .O(N__12576),
            .I(N__12570));
    LocalMux I__2028 (
            .O(N__12573),
            .I(N__12567));
    LocalMux I__2027 (
            .O(N__12570),
            .I(N__12564));
    Span12Mux_s9_h I__2026 (
            .O(N__12567),
            .I(N__12561));
    Span4Mux_h I__2025 (
            .O(N__12564),
            .I(N__12558));
    Odrv12 I__2024 (
            .O(N__12561),
            .I(n21));
    Odrv4 I__2023 (
            .O(N__12558),
            .I(n21));
    IoInMux I__2022 (
            .O(N__12553),
            .I(N__12550));
    LocalMux I__2021 (
            .O(N__12550),
            .I(N__12547));
    Span4Mux_s3_v I__2020 (
            .O(N__12547),
            .I(N__12544));
    Span4Mux_h I__2019 (
            .O(N__12544),
            .I(N__12540));
    InMux I__2018 (
            .O(N__12543),
            .I(N__12537));
    Odrv4 I__2017 (
            .O(N__12540),
            .I(LED_c));
    LocalMux I__2016 (
            .O(N__12537),
            .I(LED_c));
    CascadeMux I__2015 (
            .O(N__12532),
            .I(\receive_module.rx_counter.n3628_cascade_ ));
    InMux I__2014 (
            .O(N__12529),
            .I(N__12526));
    LocalMux I__2013 (
            .O(N__12526),
            .I(\receive_module.rx_counter.n7_adj_609 ));
    InMux I__2012 (
            .O(N__12523),
            .I(N__12520));
    LocalMux I__2011 (
            .O(N__12520),
            .I(\receive_module.rx_counter.n11 ));
    CascadeMux I__2010 (
            .O(N__12517),
            .I(\receive_module.rx_counter.n11_cascade_ ));
    InMux I__2009 (
            .O(N__12514),
            .I(N__12508));
    InMux I__2008 (
            .O(N__12513),
            .I(N__12508));
    LocalMux I__2007 (
            .O(N__12508),
            .I(\receive_module.rx_counter.old_VS ));
    InMux I__2006 (
            .O(N__12505),
            .I(N__12502));
    LocalMux I__2005 (
            .O(N__12502),
            .I(N__12499));
    Odrv4 I__2004 (
            .O(N__12499),
            .I(\transmit_module.ADDR_Y_COMPONENT_6 ));
    InMux I__2003 (
            .O(N__12496),
            .I(N__12492));
    InMux I__2002 (
            .O(N__12495),
            .I(N__12489));
    LocalMux I__2001 (
            .O(N__12492),
            .I(N__12486));
    LocalMux I__2000 (
            .O(N__12489),
            .I(\transmit_module.n106 ));
    Odrv12 I__1999 (
            .O(N__12486),
            .I(\transmit_module.n106 ));
    InMux I__1998 (
            .O(N__12481),
            .I(N__12478));
    LocalMux I__1997 (
            .O(N__12478),
            .I(N__12475));
    Odrv12 I__1996 (
            .O(N__12475),
            .I(\transmit_module.n137 ));
    CascadeMux I__1995 (
            .O(N__12472),
            .I(N__12469));
    CascadeBuf I__1994 (
            .O(N__12469),
            .I(N__12465));
    CascadeMux I__1993 (
            .O(N__12468),
            .I(N__12462));
    CascadeMux I__1992 (
            .O(N__12465),
            .I(N__12459));
    CascadeBuf I__1991 (
            .O(N__12462),
            .I(N__12456));
    CascadeBuf I__1990 (
            .O(N__12459),
            .I(N__12453));
    CascadeMux I__1989 (
            .O(N__12456),
            .I(N__12450));
    CascadeMux I__1988 (
            .O(N__12453),
            .I(N__12447));
    CascadeBuf I__1987 (
            .O(N__12450),
            .I(N__12444));
    CascadeBuf I__1986 (
            .O(N__12447),
            .I(N__12441));
    CascadeMux I__1985 (
            .O(N__12444),
            .I(N__12438));
    CascadeMux I__1984 (
            .O(N__12441),
            .I(N__12435));
    CascadeBuf I__1983 (
            .O(N__12438),
            .I(N__12432));
    CascadeBuf I__1982 (
            .O(N__12435),
            .I(N__12429));
    CascadeMux I__1981 (
            .O(N__12432),
            .I(N__12426));
    CascadeMux I__1980 (
            .O(N__12429),
            .I(N__12423));
    CascadeBuf I__1979 (
            .O(N__12426),
            .I(N__12420));
    CascadeBuf I__1978 (
            .O(N__12423),
            .I(N__12417));
    CascadeMux I__1977 (
            .O(N__12420),
            .I(N__12414));
    CascadeMux I__1976 (
            .O(N__12417),
            .I(N__12411));
    CascadeBuf I__1975 (
            .O(N__12414),
            .I(N__12408));
    CascadeBuf I__1974 (
            .O(N__12411),
            .I(N__12405));
    CascadeMux I__1973 (
            .O(N__12408),
            .I(N__12402));
    CascadeMux I__1972 (
            .O(N__12405),
            .I(N__12399));
    CascadeBuf I__1971 (
            .O(N__12402),
            .I(N__12396));
    CascadeBuf I__1970 (
            .O(N__12399),
            .I(N__12393));
    CascadeMux I__1969 (
            .O(N__12396),
            .I(N__12390));
    CascadeMux I__1968 (
            .O(N__12393),
            .I(N__12387));
    CascadeBuf I__1967 (
            .O(N__12390),
            .I(N__12384));
    CascadeBuf I__1966 (
            .O(N__12387),
            .I(N__12381));
    CascadeMux I__1965 (
            .O(N__12384),
            .I(N__12378));
    CascadeMux I__1964 (
            .O(N__12381),
            .I(N__12375));
    CascadeBuf I__1963 (
            .O(N__12378),
            .I(N__12372));
    CascadeBuf I__1962 (
            .O(N__12375),
            .I(N__12369));
    CascadeMux I__1961 (
            .O(N__12372),
            .I(N__12366));
    CascadeMux I__1960 (
            .O(N__12369),
            .I(N__12363));
    CascadeBuf I__1959 (
            .O(N__12366),
            .I(N__12360));
    CascadeBuf I__1958 (
            .O(N__12363),
            .I(N__12357));
    CascadeMux I__1957 (
            .O(N__12360),
            .I(N__12354));
    CascadeMux I__1956 (
            .O(N__12357),
            .I(N__12351));
    CascadeBuf I__1955 (
            .O(N__12354),
            .I(N__12348));
    CascadeBuf I__1954 (
            .O(N__12351),
            .I(N__12345));
    CascadeMux I__1953 (
            .O(N__12348),
            .I(N__12342));
    CascadeMux I__1952 (
            .O(N__12345),
            .I(N__12339));
    CascadeBuf I__1951 (
            .O(N__12342),
            .I(N__12336));
    CascadeBuf I__1950 (
            .O(N__12339),
            .I(N__12333));
    CascadeMux I__1949 (
            .O(N__12336),
            .I(N__12330));
    CascadeMux I__1948 (
            .O(N__12333),
            .I(N__12327));
    CascadeBuf I__1947 (
            .O(N__12330),
            .I(N__12324));
    CascadeBuf I__1946 (
            .O(N__12327),
            .I(N__12321));
    CascadeMux I__1945 (
            .O(N__12324),
            .I(N__12318));
    CascadeMux I__1944 (
            .O(N__12321),
            .I(N__12315));
    CascadeBuf I__1943 (
            .O(N__12318),
            .I(N__12312));
    CascadeBuf I__1942 (
            .O(N__12315),
            .I(N__12309));
    CascadeMux I__1941 (
            .O(N__12312),
            .I(N__12306));
    CascadeMux I__1940 (
            .O(N__12309),
            .I(N__12303));
    CascadeBuf I__1939 (
            .O(N__12306),
            .I(N__12300));
    CascadeBuf I__1938 (
            .O(N__12303),
            .I(N__12297));
    CascadeMux I__1937 (
            .O(N__12300),
            .I(N__12294));
    CascadeMux I__1936 (
            .O(N__12297),
            .I(N__12291));
    CascadeBuf I__1935 (
            .O(N__12294),
            .I(N__12288));
    InMux I__1934 (
            .O(N__12291),
            .I(N__12285));
    CascadeMux I__1933 (
            .O(N__12288),
            .I(N__12282));
    LocalMux I__1932 (
            .O(N__12285),
            .I(N__12279));
    InMux I__1931 (
            .O(N__12282),
            .I(N__12276));
    Span4Mux_v I__1930 (
            .O(N__12279),
            .I(N__12273));
    LocalMux I__1929 (
            .O(N__12276),
            .I(N__12270));
    Span4Mux_v I__1928 (
            .O(N__12273),
            .I(N__12267));
    Span4Mux_v I__1927 (
            .O(N__12270),
            .I(N__12264));
    Span4Mux_v I__1926 (
            .O(N__12267),
            .I(N__12261));
    Span4Mux_v I__1925 (
            .O(N__12264),
            .I(N__12258));
    Span4Mux_h I__1924 (
            .O(N__12261),
            .I(N__12255));
    Span4Mux_v I__1923 (
            .O(N__12258),
            .I(N__12252));
    Span4Mux_h I__1922 (
            .O(N__12255),
            .I(N__12247));
    Span4Mux_h I__1921 (
            .O(N__12252),
            .I(N__12247));
    Odrv4 I__1920 (
            .O(N__12247),
            .I(n18));
    InMux I__1919 (
            .O(N__12244),
            .I(N__12241));
    LocalMux I__1918 (
            .O(N__12241),
            .I(\transmit_module.ADDR_Y_COMPONENT_0 ));
    InMux I__1917 (
            .O(N__12238),
            .I(N__12235));
    LocalMux I__1916 (
            .O(N__12235),
            .I(\line_buffer.n3722 ));
    InMux I__1915 (
            .O(N__12232),
            .I(N__12229));
    LocalMux I__1914 (
            .O(N__12229),
            .I(N__12226));
    Odrv4 I__1913 (
            .O(N__12226),
            .I(TX_DATA_6));
    IoInMux I__1912 (
            .O(N__12223),
            .I(N__12220));
    LocalMux I__1911 (
            .O(N__12220),
            .I(N__12216));
    IoInMux I__1910 (
            .O(N__12219),
            .I(N__12212));
    Span4Mux_s2_v I__1909 (
            .O(N__12216),
            .I(N__12209));
    IoInMux I__1908 (
            .O(N__12215),
            .I(N__12206));
    LocalMux I__1907 (
            .O(N__12212),
            .I(N__12203));
    Span4Mux_h I__1906 (
            .O(N__12209),
            .I(N__12200));
    LocalMux I__1905 (
            .O(N__12206),
            .I(N__12197));
    Span4Mux_s2_v I__1904 (
            .O(N__12203),
            .I(N__12194));
    Sp12to4 I__1903 (
            .O(N__12200),
            .I(N__12191));
    Span12Mux_s1_h I__1902 (
            .O(N__12197),
            .I(N__12188));
    Span4Mux_h I__1901 (
            .O(N__12194),
            .I(N__12185));
    Span12Mux_h I__1900 (
            .O(N__12191),
            .I(N__12180));
    Span12Mux_h I__1899 (
            .O(N__12188),
            .I(N__12180));
    Span4Mux_v I__1898 (
            .O(N__12185),
            .I(N__12177));
    Odrv12 I__1897 (
            .O(N__12180),
            .I(n1792));
    Odrv4 I__1896 (
            .O(N__12177),
            .I(n1792));
    IoInMux I__1895 (
            .O(N__12172),
            .I(N__12169));
    LocalMux I__1894 (
            .O(N__12169),
            .I(N__12164));
    IoInMux I__1893 (
            .O(N__12168),
            .I(N__12161));
    IoInMux I__1892 (
            .O(N__12167),
            .I(N__12158));
    Span4Mux_s1_h I__1891 (
            .O(N__12164),
            .I(N__12155));
    LocalMux I__1890 (
            .O(N__12161),
            .I(N__12152));
    LocalMux I__1889 (
            .O(N__12158),
            .I(N__12149));
    Span4Mux_h I__1888 (
            .O(N__12155),
            .I(N__12146));
    IoSpan4Mux I__1887 (
            .O(N__12152),
            .I(N__12143));
    Span12Mux_s8_v I__1886 (
            .O(N__12149),
            .I(N__12140));
    Span4Mux_h I__1885 (
            .O(N__12146),
            .I(N__12137));
    Span4Mux_s1_v I__1884 (
            .O(N__12143),
            .I(N__12134));
    Span12Mux_h I__1883 (
            .O(N__12140),
            .I(N__12131));
    Span4Mux_h I__1882 (
            .O(N__12137),
            .I(N__12126));
    Span4Mux_v I__1881 (
            .O(N__12134),
            .I(N__12126));
    Odrv12 I__1880 (
            .O(N__12131),
            .I(n1798));
    Odrv4 I__1879 (
            .O(N__12126),
            .I(n1798));
    InMux I__1878 (
            .O(N__12121),
            .I(N__12118));
    LocalMux I__1877 (
            .O(N__12118),
            .I(N__12115));
    Span4Mux_h I__1876 (
            .O(N__12115),
            .I(N__12112));
    Span4Mux_h I__1875 (
            .O(N__12112),
            .I(N__12109));
    Span4Mux_h I__1874 (
            .O(N__12109),
            .I(N__12106));
    Odrv4 I__1873 (
            .O(N__12106),
            .I(\line_buffer.n448 ));
    InMux I__1872 (
            .O(N__12103),
            .I(N__12100));
    LocalMux I__1871 (
            .O(N__12100),
            .I(N__12097));
    Span4Mux_v I__1870 (
            .O(N__12097),
            .I(N__12094));
    Span4Mux_h I__1869 (
            .O(N__12094),
            .I(N__12091));
    Odrv4 I__1868 (
            .O(N__12091),
            .I(\line_buffer.n440 ));
    InMux I__1867 (
            .O(N__12088),
            .I(N__12085));
    LocalMux I__1866 (
            .O(N__12085),
            .I(N__12082));
    Odrv12 I__1865 (
            .O(N__12082),
            .I(\line_buffer.n3679 ));
    InMux I__1864 (
            .O(N__12079),
            .I(N__12075));
    InMux I__1863 (
            .O(N__12078),
            .I(N__12072));
    LocalMux I__1862 (
            .O(N__12075),
            .I(N__12069));
    LocalMux I__1861 (
            .O(N__12072),
            .I(N__12066));
    Span4Mux_v I__1860 (
            .O(N__12069),
            .I(N__12063));
    Span4Mux_v I__1859 (
            .O(N__12066),
            .I(N__12060));
    Span4Mux_v I__1858 (
            .O(N__12063),
            .I(N__12057));
    Odrv4 I__1857 (
            .O(N__12060),
            .I(\transmit_module.n116 ));
    Odrv4 I__1856 (
            .O(N__12057),
            .I(\transmit_module.n116 ));
    InMux I__1855 (
            .O(N__12052),
            .I(N__12048));
    InMux I__1854 (
            .O(N__12051),
            .I(N__12045));
    LocalMux I__1853 (
            .O(N__12048),
            .I(N__12042));
    LocalMux I__1852 (
            .O(N__12045),
            .I(N__12039));
    Span12Mux_v I__1851 (
            .O(N__12042),
            .I(N__12036));
    Odrv4 I__1850 (
            .O(N__12039),
            .I(\transmit_module.n147 ));
    Odrv12 I__1849 (
            .O(N__12036),
            .I(\transmit_module.n147 ));
    CascadeMux I__1848 (
            .O(N__12031),
            .I(N__12028));
    CascadeBuf I__1847 (
            .O(N__12028),
            .I(N__12024));
    CascadeMux I__1846 (
            .O(N__12027),
            .I(N__12021));
    CascadeMux I__1845 (
            .O(N__12024),
            .I(N__12018));
    CascadeBuf I__1844 (
            .O(N__12021),
            .I(N__12015));
    CascadeBuf I__1843 (
            .O(N__12018),
            .I(N__12012));
    CascadeMux I__1842 (
            .O(N__12015),
            .I(N__12009));
    CascadeMux I__1841 (
            .O(N__12012),
            .I(N__12006));
    CascadeBuf I__1840 (
            .O(N__12009),
            .I(N__12003));
    CascadeBuf I__1839 (
            .O(N__12006),
            .I(N__12000));
    CascadeMux I__1838 (
            .O(N__12003),
            .I(N__11997));
    CascadeMux I__1837 (
            .O(N__12000),
            .I(N__11994));
    CascadeBuf I__1836 (
            .O(N__11997),
            .I(N__11991));
    CascadeBuf I__1835 (
            .O(N__11994),
            .I(N__11988));
    CascadeMux I__1834 (
            .O(N__11991),
            .I(N__11985));
    CascadeMux I__1833 (
            .O(N__11988),
            .I(N__11982));
    CascadeBuf I__1832 (
            .O(N__11985),
            .I(N__11979));
    CascadeBuf I__1831 (
            .O(N__11982),
            .I(N__11976));
    CascadeMux I__1830 (
            .O(N__11979),
            .I(N__11973));
    CascadeMux I__1829 (
            .O(N__11976),
            .I(N__11970));
    CascadeBuf I__1828 (
            .O(N__11973),
            .I(N__11967));
    CascadeBuf I__1827 (
            .O(N__11970),
            .I(N__11964));
    CascadeMux I__1826 (
            .O(N__11967),
            .I(N__11961));
    CascadeMux I__1825 (
            .O(N__11964),
            .I(N__11958));
    CascadeBuf I__1824 (
            .O(N__11961),
            .I(N__11955));
    CascadeBuf I__1823 (
            .O(N__11958),
            .I(N__11952));
    CascadeMux I__1822 (
            .O(N__11955),
            .I(N__11949));
    CascadeMux I__1821 (
            .O(N__11952),
            .I(N__11946));
    CascadeBuf I__1820 (
            .O(N__11949),
            .I(N__11943));
    CascadeBuf I__1819 (
            .O(N__11946),
            .I(N__11940));
    CascadeMux I__1818 (
            .O(N__11943),
            .I(N__11937));
    CascadeMux I__1817 (
            .O(N__11940),
            .I(N__11934));
    CascadeBuf I__1816 (
            .O(N__11937),
            .I(N__11931));
    CascadeBuf I__1815 (
            .O(N__11934),
            .I(N__11928));
    CascadeMux I__1814 (
            .O(N__11931),
            .I(N__11925));
    CascadeMux I__1813 (
            .O(N__11928),
            .I(N__11922));
    CascadeBuf I__1812 (
            .O(N__11925),
            .I(N__11919));
    CascadeBuf I__1811 (
            .O(N__11922),
            .I(N__11916));
    CascadeMux I__1810 (
            .O(N__11919),
            .I(N__11913));
    CascadeMux I__1809 (
            .O(N__11916),
            .I(N__11910));
    CascadeBuf I__1808 (
            .O(N__11913),
            .I(N__11907));
    CascadeBuf I__1807 (
            .O(N__11910),
            .I(N__11904));
    CascadeMux I__1806 (
            .O(N__11907),
            .I(N__11901));
    CascadeMux I__1805 (
            .O(N__11904),
            .I(N__11898));
    CascadeBuf I__1804 (
            .O(N__11901),
            .I(N__11895));
    CascadeBuf I__1803 (
            .O(N__11898),
            .I(N__11892));
    CascadeMux I__1802 (
            .O(N__11895),
            .I(N__11889));
    CascadeMux I__1801 (
            .O(N__11892),
            .I(N__11886));
    CascadeBuf I__1800 (
            .O(N__11889),
            .I(N__11883));
    CascadeBuf I__1799 (
            .O(N__11886),
            .I(N__11880));
    CascadeMux I__1798 (
            .O(N__11883),
            .I(N__11877));
    CascadeMux I__1797 (
            .O(N__11880),
            .I(N__11874));
    CascadeBuf I__1796 (
            .O(N__11877),
            .I(N__11871));
    CascadeBuf I__1795 (
            .O(N__11874),
            .I(N__11868));
    CascadeMux I__1794 (
            .O(N__11871),
            .I(N__11865));
    CascadeMux I__1793 (
            .O(N__11868),
            .I(N__11862));
    CascadeBuf I__1792 (
            .O(N__11865),
            .I(N__11859));
    CascadeBuf I__1791 (
            .O(N__11862),
            .I(N__11856));
    CascadeMux I__1790 (
            .O(N__11859),
            .I(N__11853));
    CascadeMux I__1789 (
            .O(N__11856),
            .I(N__11850));
    CascadeBuf I__1788 (
            .O(N__11853),
            .I(N__11847));
    InMux I__1787 (
            .O(N__11850),
            .I(N__11844));
    CascadeMux I__1786 (
            .O(N__11847),
            .I(N__11841));
    LocalMux I__1785 (
            .O(N__11844),
            .I(N__11838));
    InMux I__1784 (
            .O(N__11841),
            .I(N__11835));
    Span4Mux_v I__1783 (
            .O(N__11838),
            .I(N__11832));
    LocalMux I__1782 (
            .O(N__11835),
            .I(N__11829));
    Span4Mux_h I__1781 (
            .O(N__11832),
            .I(N__11826));
    Span4Mux_h I__1780 (
            .O(N__11829),
            .I(N__11823));
    Span4Mux_h I__1779 (
            .O(N__11826),
            .I(N__11820));
    Span4Mux_v I__1778 (
            .O(N__11823),
            .I(N__11817));
    Odrv4 I__1777 (
            .O(N__11820),
            .I(n28));
    Odrv4 I__1776 (
            .O(N__11817),
            .I(n28));
    InMux I__1775 (
            .O(N__11812),
            .I(N__11809));
    LocalMux I__1774 (
            .O(N__11809),
            .I(\transmit_module.n146 ));
    CascadeMux I__1773 (
            .O(N__11806),
            .I(\transmit_module.n146_cascade_ ));
    InMux I__1772 (
            .O(N__11803),
            .I(N__11799));
    InMux I__1771 (
            .O(N__11802),
            .I(N__11796));
    LocalMux I__1770 (
            .O(N__11799),
            .I(N__11793));
    LocalMux I__1769 (
            .O(N__11796),
            .I(\transmit_module.n115 ));
    Odrv4 I__1768 (
            .O(N__11793),
            .I(\transmit_module.n115 ));
    CascadeMux I__1767 (
            .O(N__11788),
            .I(N__11785));
    CascadeBuf I__1766 (
            .O(N__11785),
            .I(N__11781));
    CascadeMux I__1765 (
            .O(N__11784),
            .I(N__11778));
    CascadeMux I__1764 (
            .O(N__11781),
            .I(N__11775));
    CascadeBuf I__1763 (
            .O(N__11778),
            .I(N__11772));
    CascadeBuf I__1762 (
            .O(N__11775),
            .I(N__11769));
    CascadeMux I__1761 (
            .O(N__11772),
            .I(N__11766));
    CascadeMux I__1760 (
            .O(N__11769),
            .I(N__11763));
    CascadeBuf I__1759 (
            .O(N__11766),
            .I(N__11760));
    CascadeBuf I__1758 (
            .O(N__11763),
            .I(N__11757));
    CascadeMux I__1757 (
            .O(N__11760),
            .I(N__11754));
    CascadeMux I__1756 (
            .O(N__11757),
            .I(N__11751));
    CascadeBuf I__1755 (
            .O(N__11754),
            .I(N__11748));
    CascadeBuf I__1754 (
            .O(N__11751),
            .I(N__11745));
    CascadeMux I__1753 (
            .O(N__11748),
            .I(N__11742));
    CascadeMux I__1752 (
            .O(N__11745),
            .I(N__11739));
    CascadeBuf I__1751 (
            .O(N__11742),
            .I(N__11736));
    CascadeBuf I__1750 (
            .O(N__11739),
            .I(N__11733));
    CascadeMux I__1749 (
            .O(N__11736),
            .I(N__11730));
    CascadeMux I__1748 (
            .O(N__11733),
            .I(N__11727));
    CascadeBuf I__1747 (
            .O(N__11730),
            .I(N__11724));
    CascadeBuf I__1746 (
            .O(N__11727),
            .I(N__11721));
    CascadeMux I__1745 (
            .O(N__11724),
            .I(N__11718));
    CascadeMux I__1744 (
            .O(N__11721),
            .I(N__11715));
    CascadeBuf I__1743 (
            .O(N__11718),
            .I(N__11712));
    CascadeBuf I__1742 (
            .O(N__11715),
            .I(N__11709));
    CascadeMux I__1741 (
            .O(N__11712),
            .I(N__11706));
    CascadeMux I__1740 (
            .O(N__11709),
            .I(N__11703));
    CascadeBuf I__1739 (
            .O(N__11706),
            .I(N__11700));
    CascadeBuf I__1738 (
            .O(N__11703),
            .I(N__11697));
    CascadeMux I__1737 (
            .O(N__11700),
            .I(N__11694));
    CascadeMux I__1736 (
            .O(N__11697),
            .I(N__11691));
    CascadeBuf I__1735 (
            .O(N__11694),
            .I(N__11688));
    CascadeBuf I__1734 (
            .O(N__11691),
            .I(N__11685));
    CascadeMux I__1733 (
            .O(N__11688),
            .I(N__11682));
    CascadeMux I__1732 (
            .O(N__11685),
            .I(N__11679));
    CascadeBuf I__1731 (
            .O(N__11682),
            .I(N__11676));
    CascadeBuf I__1730 (
            .O(N__11679),
            .I(N__11673));
    CascadeMux I__1729 (
            .O(N__11676),
            .I(N__11670));
    CascadeMux I__1728 (
            .O(N__11673),
            .I(N__11667));
    CascadeBuf I__1727 (
            .O(N__11670),
            .I(N__11664));
    CascadeBuf I__1726 (
            .O(N__11667),
            .I(N__11661));
    CascadeMux I__1725 (
            .O(N__11664),
            .I(N__11658));
    CascadeMux I__1724 (
            .O(N__11661),
            .I(N__11655));
    CascadeBuf I__1723 (
            .O(N__11658),
            .I(N__11652));
    CascadeBuf I__1722 (
            .O(N__11655),
            .I(N__11649));
    CascadeMux I__1721 (
            .O(N__11652),
            .I(N__11646));
    CascadeMux I__1720 (
            .O(N__11649),
            .I(N__11643));
    CascadeBuf I__1719 (
            .O(N__11646),
            .I(N__11640));
    CascadeBuf I__1718 (
            .O(N__11643),
            .I(N__11637));
    CascadeMux I__1717 (
            .O(N__11640),
            .I(N__11634));
    CascadeMux I__1716 (
            .O(N__11637),
            .I(N__11631));
    CascadeBuf I__1715 (
            .O(N__11634),
            .I(N__11628));
    CascadeBuf I__1714 (
            .O(N__11631),
            .I(N__11625));
    CascadeMux I__1713 (
            .O(N__11628),
            .I(N__11622));
    CascadeMux I__1712 (
            .O(N__11625),
            .I(N__11619));
    CascadeBuf I__1711 (
            .O(N__11622),
            .I(N__11616));
    CascadeBuf I__1710 (
            .O(N__11619),
            .I(N__11613));
    CascadeMux I__1709 (
            .O(N__11616),
            .I(N__11610));
    CascadeMux I__1708 (
            .O(N__11613),
            .I(N__11607));
    CascadeBuf I__1707 (
            .O(N__11610),
            .I(N__11604));
    InMux I__1706 (
            .O(N__11607),
            .I(N__11601));
    CascadeMux I__1705 (
            .O(N__11604),
            .I(N__11598));
    LocalMux I__1704 (
            .O(N__11601),
            .I(N__11595));
    InMux I__1703 (
            .O(N__11598),
            .I(N__11592));
    Span4Mux_v I__1702 (
            .O(N__11595),
            .I(N__11589));
    LocalMux I__1701 (
            .O(N__11592),
            .I(N__11586));
    Span4Mux_v I__1700 (
            .O(N__11589),
            .I(N__11583));
    Span4Mux_v I__1699 (
            .O(N__11586),
            .I(N__11580));
    Span4Mux_v I__1698 (
            .O(N__11583),
            .I(N__11577));
    Span4Mux_v I__1697 (
            .O(N__11580),
            .I(N__11574));
    Span4Mux_v I__1696 (
            .O(N__11577),
            .I(N__11571));
    Span4Mux_v I__1695 (
            .O(N__11574),
            .I(N__11568));
    Span4Mux_h I__1694 (
            .O(N__11571),
            .I(N__11565));
    Span4Mux_v I__1693 (
            .O(N__11568),
            .I(N__11562));
    Span4Mux_h I__1692 (
            .O(N__11565),
            .I(N__11557));
    Span4Mux_h I__1691 (
            .O(N__11562),
            .I(N__11557));
    Odrv4 I__1690 (
            .O(N__11557),
            .I(n27));
    InMux I__1689 (
            .O(N__11554),
            .I(N__11551));
    LocalMux I__1688 (
            .O(N__11551),
            .I(N__11548));
    Odrv4 I__1687 (
            .O(N__11548),
            .I(\transmit_module.Y_DELTA_PATTERN_2 ));
    InMux I__1686 (
            .O(N__11545),
            .I(N__11542));
    LocalMux I__1685 (
            .O(N__11542),
            .I(\transmit_module.Y_DELTA_PATTERN_1 ));
    InMux I__1684 (
            .O(N__11539),
            .I(N__11536));
    LocalMux I__1683 (
            .O(N__11536),
            .I(\transmit_module.Y_DELTA_PATTERN_9 ));
    InMux I__1682 (
            .O(N__11533),
            .I(N__11530));
    LocalMux I__1681 (
            .O(N__11530),
            .I(N__11527));
    Odrv12 I__1680 (
            .O(N__11527),
            .I(\transmit_module.Y_DELTA_PATTERN_8 ));
    InMux I__1679 (
            .O(N__11524),
            .I(N__11521));
    LocalMux I__1678 (
            .O(N__11521),
            .I(\transmit_module.Y_DELTA_PATTERN_10 ));
    InMux I__1677 (
            .O(N__11518),
            .I(N__11515));
    LocalMux I__1676 (
            .O(N__11515),
            .I(N__11512));
    Span4Mux_h I__1675 (
            .O(N__11512),
            .I(N__11509));
    Span4Mux_h I__1674 (
            .O(N__11509),
            .I(N__11506));
    Span4Mux_v I__1673 (
            .O(N__11506),
            .I(N__11503));
    Span4Mux_v I__1672 (
            .O(N__11503),
            .I(N__11500));
    Odrv4 I__1671 (
            .O(N__11500),
            .I(\line_buffer.n507 ));
    CascadeMux I__1670 (
            .O(N__11497),
            .I(N__11494));
    InMux I__1669 (
            .O(N__11494),
            .I(N__11491));
    LocalMux I__1668 (
            .O(N__11491),
            .I(N__11488));
    Span4Mux_v I__1667 (
            .O(N__11488),
            .I(N__11485));
    Sp12to4 I__1666 (
            .O(N__11485),
            .I(N__11482));
    Span12Mux_h I__1665 (
            .O(N__11482),
            .I(N__11479));
    Odrv12 I__1664 (
            .O(N__11479),
            .I(\line_buffer.n499 ));
    InMux I__1663 (
            .O(N__11476),
            .I(N__11473));
    LocalMux I__1662 (
            .O(N__11473),
            .I(\line_buffer.n3752 ));
    CascadeMux I__1661 (
            .O(N__11470),
            .I(\transmit_module.n141_cascade_ ));
    CascadeMux I__1660 (
            .O(N__11467),
            .I(\transmit_module.n137_cascade_ ));
    CascadeMux I__1659 (
            .O(N__11464),
            .I(N__11461));
    InMux I__1658 (
            .O(N__11461),
            .I(N__11458));
    LocalMux I__1657 (
            .O(N__11458),
            .I(\transmit_module.ADDR_Y_COMPONENT_1 ));
    CascadeMux I__1656 (
            .O(N__11455),
            .I(N__11452));
    InMux I__1655 (
            .O(N__11452),
            .I(N__11449));
    LocalMux I__1654 (
            .O(N__11449),
            .I(\transmit_module.ADDR_Y_COMPONENT_10 ));
    InMux I__1653 (
            .O(N__11446),
            .I(N__11443));
    LocalMux I__1652 (
            .O(N__11443),
            .I(\transmit_module.video_signal_controller.n3632 ));
    InMux I__1651 (
            .O(N__11440),
            .I(N__11437));
    LocalMux I__1650 (
            .O(N__11437),
            .I(N__11434));
    Odrv4 I__1649 (
            .O(N__11434),
            .I(\transmit_module.video_signal_controller.n18_adj_616 ));
    CascadeMux I__1648 (
            .O(N__11431),
            .I(N__11428));
    InMux I__1647 (
            .O(N__11428),
            .I(N__11425));
    LocalMux I__1646 (
            .O(N__11425),
            .I(\transmit_module.video_signal_controller.n3614 ));
    InMux I__1645 (
            .O(N__11422),
            .I(N__11419));
    LocalMux I__1644 (
            .O(N__11419),
            .I(N__11416));
    Span4Mux_h I__1643 (
            .O(N__11416),
            .I(N__11411));
    InMux I__1642 (
            .O(N__11415),
            .I(N__11408));
    InMux I__1641 (
            .O(N__11414),
            .I(N__11405));
    Odrv4 I__1640 (
            .O(N__11411),
            .I(\transmit_module.video_signal_controller.VGA_Y_10 ));
    LocalMux I__1639 (
            .O(N__11408),
            .I(\transmit_module.video_signal_controller.VGA_Y_10 ));
    LocalMux I__1638 (
            .O(N__11405),
            .I(\transmit_module.video_signal_controller.VGA_Y_10 ));
    InMux I__1637 (
            .O(N__11398),
            .I(N__11395));
    LocalMux I__1636 (
            .O(N__11395),
            .I(N__11392));
    Span4Mux_h I__1635 (
            .O(N__11392),
            .I(N__11388));
    InMux I__1634 (
            .O(N__11391),
            .I(N__11385));
    Odrv4 I__1633 (
            .O(N__11388),
            .I(\transmit_module.video_signal_controller.VGA_Y_0 ));
    LocalMux I__1632 (
            .O(N__11385),
            .I(\transmit_module.video_signal_controller.VGA_Y_0 ));
    InMux I__1631 (
            .O(N__11380),
            .I(N__11374));
    InMux I__1630 (
            .O(N__11379),
            .I(N__11369));
    InMux I__1629 (
            .O(N__11378),
            .I(N__11369));
    InMux I__1628 (
            .O(N__11377),
            .I(N__11366));
    LocalMux I__1627 (
            .O(N__11374),
            .I(N__11361));
    LocalMux I__1626 (
            .O(N__11369),
            .I(N__11361));
    LocalMux I__1625 (
            .O(N__11366),
            .I(\transmit_module.video_signal_controller.VGA_Y_3 ));
    Odrv4 I__1624 (
            .O(N__11361),
            .I(\transmit_module.video_signal_controller.VGA_Y_3 ));
    CascadeMux I__1623 (
            .O(N__11356),
            .I(\transmit_module.video_signal_controller.n3626_cascade_ ));
    InMux I__1622 (
            .O(N__11353),
            .I(N__11349));
    CascadeMux I__1621 (
            .O(N__11352),
            .I(N__11345));
    LocalMux I__1620 (
            .O(N__11349),
            .I(N__11341));
    InMux I__1619 (
            .O(N__11348),
            .I(N__11338));
    InMux I__1618 (
            .O(N__11345),
            .I(N__11333));
    InMux I__1617 (
            .O(N__11344),
            .I(N__11333));
    Odrv4 I__1616 (
            .O(N__11341),
            .I(\transmit_module.video_signal_controller.VGA_Y_1 ));
    LocalMux I__1615 (
            .O(N__11338),
            .I(\transmit_module.video_signal_controller.VGA_Y_1 ));
    LocalMux I__1614 (
            .O(N__11333),
            .I(\transmit_module.video_signal_controller.VGA_Y_1 ));
    InMux I__1613 (
            .O(N__11326),
            .I(N__11323));
    LocalMux I__1612 (
            .O(N__11323),
            .I(N__11320));
    Odrv4 I__1611 (
            .O(N__11320),
            .I(\transmit_module.n111 ));
    InMux I__1610 (
            .O(N__11317),
            .I(N__11314));
    LocalMux I__1609 (
            .O(N__11314),
            .I(N__11311));
    Span4Mux_h I__1608 (
            .O(N__11311),
            .I(N__11308));
    Odrv4 I__1607 (
            .O(N__11308),
            .I(\transmit_module.n143 ));
    CascadeMux I__1606 (
            .O(N__11305),
            .I(\transmit_module.n143_cascade_ ));
    InMux I__1605 (
            .O(N__11302),
            .I(N__11299));
    LocalMux I__1604 (
            .O(N__11299),
            .I(\transmit_module.n112 ));
    InMux I__1603 (
            .O(N__11296),
            .I(N__11292));
    InMux I__1602 (
            .O(N__11295),
            .I(N__11289));
    LocalMux I__1601 (
            .O(N__11292),
            .I(\transmit_module.n142 ));
    LocalMux I__1600 (
            .O(N__11289),
            .I(\transmit_module.n142 ));
    InMux I__1599 (
            .O(N__11284),
            .I(N__11278));
    InMux I__1598 (
            .O(N__11283),
            .I(N__11271));
    InMux I__1597 (
            .O(N__11282),
            .I(N__11271));
    InMux I__1596 (
            .O(N__11281),
            .I(N__11271));
    LocalMux I__1595 (
            .O(N__11278),
            .I(\receive_module.rx_counter.Y_3 ));
    LocalMux I__1594 (
            .O(N__11271),
            .I(\receive_module.rx_counter.Y_3 ));
    InMux I__1593 (
            .O(N__11266),
            .I(N__11260));
    InMux I__1592 (
            .O(N__11265),
            .I(N__11253));
    InMux I__1591 (
            .O(N__11264),
            .I(N__11253));
    InMux I__1590 (
            .O(N__11263),
            .I(N__11253));
    LocalMux I__1589 (
            .O(N__11260),
            .I(\receive_module.rx_counter.Y_2 ));
    LocalMux I__1588 (
            .O(N__11253),
            .I(\receive_module.rx_counter.Y_2 ));
    CascadeMux I__1587 (
            .O(N__11248),
            .I(N__11242));
    InMux I__1586 (
            .O(N__11247),
            .I(N__11239));
    InMux I__1585 (
            .O(N__11246),
            .I(N__11232));
    InMux I__1584 (
            .O(N__11245),
            .I(N__11232));
    InMux I__1583 (
            .O(N__11242),
            .I(N__11232));
    LocalMux I__1582 (
            .O(N__11239),
            .I(\receive_module.rx_counter.Y_1 ));
    LocalMux I__1581 (
            .O(N__11232),
            .I(\receive_module.rx_counter.Y_1 ));
    InMux I__1580 (
            .O(N__11227),
            .I(N__11222));
    InMux I__1579 (
            .O(N__11226),
            .I(N__11217));
    InMux I__1578 (
            .O(N__11225),
            .I(N__11217));
    LocalMux I__1577 (
            .O(N__11222),
            .I(\receive_module.rx_counter.Y_5 ));
    LocalMux I__1576 (
            .O(N__11217),
            .I(\receive_module.rx_counter.Y_5 ));
    InMux I__1575 (
            .O(N__11212),
            .I(N__11207));
    InMux I__1574 (
            .O(N__11211),
            .I(N__11204));
    InMux I__1573 (
            .O(N__11210),
            .I(N__11201));
    LocalMux I__1572 (
            .O(N__11207),
            .I(\receive_module.rx_counter.Y_6 ));
    LocalMux I__1571 (
            .O(N__11204),
            .I(\receive_module.rx_counter.Y_6 ));
    LocalMux I__1570 (
            .O(N__11201),
            .I(\receive_module.rx_counter.Y_6 ));
    InMux I__1569 (
            .O(N__11194),
            .I(N__11191));
    LocalMux I__1568 (
            .O(N__11191),
            .I(\receive_module.rx_counter.n4_adj_604 ));
    CascadeMux I__1567 (
            .O(N__11188),
            .I(\receive_module.rx_counter.n5_cascade_ ));
    InMux I__1566 (
            .O(N__11185),
            .I(N__11182));
    LocalMux I__1565 (
            .O(N__11182),
            .I(\receive_module.rx_counter.n3548 ));
    InMux I__1564 (
            .O(N__11179),
            .I(N__11173));
    InMux I__1563 (
            .O(N__11178),
            .I(N__11170));
    InMux I__1562 (
            .O(N__11177),
            .I(N__11165));
    InMux I__1561 (
            .O(N__11176),
            .I(N__11165));
    LocalMux I__1560 (
            .O(N__11173),
            .I(\receive_module.rx_counter.Y_0 ));
    LocalMux I__1559 (
            .O(N__11170),
            .I(\receive_module.rx_counter.Y_0 ));
    LocalMux I__1558 (
            .O(N__11165),
            .I(\receive_module.rx_counter.Y_0 ));
    InMux I__1557 (
            .O(N__11158),
            .I(N__11155));
    LocalMux I__1556 (
            .O(N__11155),
            .I(\receive_module.rx_counter.n14_adj_611 ));
    CascadeMux I__1555 (
            .O(N__11152),
            .I(N__11149));
    InMux I__1554 (
            .O(N__11149),
            .I(N__11146));
    LocalMux I__1553 (
            .O(N__11146),
            .I(\receive_module.rx_counter.n10_adj_610 ));
    InMux I__1552 (
            .O(N__11143),
            .I(N__11140));
    LocalMux I__1551 (
            .O(N__11140),
            .I(\transmit_module.ADDR_Y_COMPONENT_7 ));
    InMux I__1550 (
            .O(N__11137),
            .I(N__11134));
    LocalMux I__1549 (
            .O(N__11134),
            .I(N__11131));
    Odrv12 I__1548 (
            .O(N__11131),
            .I(\transmit_module.X_DELTA_PATTERN_1 ));
    CEMux I__1547 (
            .O(N__11128),
            .I(N__11124));
    CEMux I__1546 (
            .O(N__11127),
            .I(N__11119));
    LocalMux I__1545 (
            .O(N__11124),
            .I(N__11116));
    CEMux I__1544 (
            .O(N__11123),
            .I(N__11113));
    CEMux I__1543 (
            .O(N__11122),
            .I(N__11110));
    LocalMux I__1542 (
            .O(N__11119),
            .I(N__11107));
    Span4Mux_h I__1541 (
            .O(N__11116),
            .I(N__11103));
    LocalMux I__1540 (
            .O(N__11113),
            .I(N__11100));
    LocalMux I__1539 (
            .O(N__11110),
            .I(N__11097));
    Span4Mux_v I__1538 (
            .O(N__11107),
            .I(N__11094));
    CEMux I__1537 (
            .O(N__11106),
            .I(N__11091));
    Span4Mux_h I__1536 (
            .O(N__11103),
            .I(N__11086));
    Span4Mux_h I__1535 (
            .O(N__11100),
            .I(N__11086));
    Span4Mux_h I__1534 (
            .O(N__11097),
            .I(N__11079));
    Span4Mux_h I__1533 (
            .O(N__11094),
            .I(N__11079));
    LocalMux I__1532 (
            .O(N__11091),
            .I(N__11079));
    Odrv4 I__1531 (
            .O(N__11086),
            .I(\transmit_module.n2093 ));
    Odrv4 I__1530 (
            .O(N__11079),
            .I(\transmit_module.n2093 ));
    CEMux I__1529 (
            .O(N__11074),
            .I(N__11070));
    CEMux I__1528 (
            .O(N__11073),
            .I(N__11066));
    LocalMux I__1527 (
            .O(N__11070),
            .I(N__11061));
    CEMux I__1526 (
            .O(N__11069),
            .I(N__11058));
    LocalMux I__1525 (
            .O(N__11066),
            .I(N__11055));
    CEMux I__1524 (
            .O(N__11065),
            .I(N__11052));
    SRMux I__1523 (
            .O(N__11064),
            .I(N__11049));
    Span4Mux_v I__1522 (
            .O(N__11061),
            .I(N__11044));
    LocalMux I__1521 (
            .O(N__11058),
            .I(N__11044));
    Span4Mux_v I__1520 (
            .O(N__11055),
            .I(N__11041));
    LocalMux I__1519 (
            .O(N__11052),
            .I(N__11038));
    LocalMux I__1518 (
            .O(N__11049),
            .I(N__11035));
    Span4Mux_v I__1517 (
            .O(N__11044),
            .I(N__11032));
    Span4Mux_h I__1516 (
            .O(N__11041),
            .I(N__11027));
    Span4Mux_v I__1515 (
            .O(N__11038),
            .I(N__11027));
    Span4Mux_v I__1514 (
            .O(N__11035),
            .I(N__11024));
    Odrv4 I__1513 (
            .O(N__11032),
            .I(\transmit_module.n2147 ));
    Odrv4 I__1512 (
            .O(N__11027),
            .I(\transmit_module.n2147 ));
    Odrv4 I__1511 (
            .O(N__11024),
            .I(\transmit_module.n2147 ));
    InMux I__1510 (
            .O(N__11017),
            .I(N__11013));
    InMux I__1509 (
            .O(N__11016),
            .I(N__11008));
    LocalMux I__1508 (
            .O(N__11013),
            .I(N__11005));
    InMux I__1507 (
            .O(N__11012),
            .I(N__11000));
    InMux I__1506 (
            .O(N__11011),
            .I(N__11000));
    LocalMux I__1505 (
            .O(N__11008),
            .I(\transmit_module.video_signal_controller.VGA_Y_4 ));
    Odrv4 I__1504 (
            .O(N__11005),
            .I(\transmit_module.video_signal_controller.VGA_Y_4 ));
    LocalMux I__1503 (
            .O(N__11000),
            .I(\transmit_module.video_signal_controller.VGA_Y_4 ));
    InMux I__1502 (
            .O(N__10993),
            .I(N__10989));
    InMux I__1501 (
            .O(N__10992),
            .I(N__10985));
    LocalMux I__1500 (
            .O(N__10989),
            .I(N__10982));
    InMux I__1499 (
            .O(N__10988),
            .I(N__10978));
    LocalMux I__1498 (
            .O(N__10985),
            .I(N__10973));
    Span4Mux_v I__1497 (
            .O(N__10982),
            .I(N__10973));
    InMux I__1496 (
            .O(N__10981),
            .I(N__10970));
    LocalMux I__1495 (
            .O(N__10978),
            .I(\transmit_module.video_signal_controller.VGA_Y_8 ));
    Odrv4 I__1494 (
            .O(N__10973),
            .I(\transmit_module.video_signal_controller.VGA_Y_8 ));
    LocalMux I__1493 (
            .O(N__10970),
            .I(\transmit_module.video_signal_controller.VGA_Y_8 ));
    InMux I__1492 (
            .O(N__10963),
            .I(N__10960));
    LocalMux I__1491 (
            .O(N__10960),
            .I(\transmit_module.ADDR_Y_COMPONENT_4 ));
    InMux I__1490 (
            .O(N__10957),
            .I(N__10954));
    LocalMux I__1489 (
            .O(N__10954),
            .I(\transmit_module.ADDR_Y_COMPONENT_5 ));
    InMux I__1488 (
            .O(N__10951),
            .I(N__10948));
    LocalMux I__1487 (
            .O(N__10948),
            .I(N__10945));
    Span4Mux_v I__1486 (
            .O(N__10945),
            .I(N__10942));
    Span4Mux_h I__1485 (
            .O(N__10942),
            .I(N__10939));
    Odrv4 I__1484 (
            .O(N__10939),
            .I(\line_buffer.n571 ));
    InMux I__1483 (
            .O(N__10936),
            .I(N__10933));
    LocalMux I__1482 (
            .O(N__10933),
            .I(N__10930));
    Span12Mux_v I__1481 (
            .O(N__10930),
            .I(N__10927));
    Span12Mux_h I__1480 (
            .O(N__10927),
            .I(N__10924));
    Odrv12 I__1479 (
            .O(N__10924),
            .I(\line_buffer.n563 ));
    InMux I__1478 (
            .O(N__10921),
            .I(N__10918));
    LocalMux I__1477 (
            .O(N__10918),
            .I(N__10915));
    Span4Mux_v I__1476 (
            .O(N__10915),
            .I(N__10912));
    Span4Mux_h I__1475 (
            .O(N__10912),
            .I(N__10909));
    Odrv4 I__1474 (
            .O(N__10909),
            .I(\line_buffer.n514 ));
    CascadeMux I__1473 (
            .O(N__10906),
            .I(N__10903));
    InMux I__1472 (
            .O(N__10903),
            .I(N__10900));
    LocalMux I__1471 (
            .O(N__10900),
            .I(N__10897));
    Span12Mux_v I__1470 (
            .O(N__10897),
            .I(N__10894));
    Span12Mux_v I__1469 (
            .O(N__10894),
            .I(N__10891));
    Span12Mux_h I__1468 (
            .O(N__10891),
            .I(N__10888));
    Odrv12 I__1467 (
            .O(N__10888),
            .I(\line_buffer.n506 ));
    InMux I__1466 (
            .O(N__10885),
            .I(N__10882));
    LocalMux I__1465 (
            .O(N__10882),
            .I(\line_buffer.n3764 ));
    InMux I__1464 (
            .O(N__10879),
            .I(N__10876));
    LocalMux I__1463 (
            .O(N__10876),
            .I(N__10873));
    Span4Mux_h I__1462 (
            .O(N__10873),
            .I(N__10870));
    Span4Mux_h I__1461 (
            .O(N__10870),
            .I(N__10867));
    Odrv4 I__1460 (
            .O(N__10867),
            .I(\line_buffer.n513 ));
    InMux I__1459 (
            .O(N__10864),
            .I(N__10861));
    LocalMux I__1458 (
            .O(N__10861),
            .I(N__10858));
    Span12Mux_v I__1457 (
            .O(N__10858),
            .I(N__10855));
    Span12Mux_v I__1456 (
            .O(N__10855),
            .I(N__10852));
    Span12Mux_h I__1455 (
            .O(N__10852),
            .I(N__10849));
    Odrv12 I__1454 (
            .O(N__10849),
            .I(\line_buffer.n505 ));
    CascadeMux I__1453 (
            .O(N__10846),
            .I(\line_buffer.n3646_cascade_ ));
    InMux I__1452 (
            .O(N__10843),
            .I(N__10840));
    LocalMux I__1451 (
            .O(N__10840),
            .I(\line_buffer.n3647 ));
    CascadeMux I__1450 (
            .O(N__10837),
            .I(\transmit_module.n112_cascade_ ));
    CascadeMux I__1449 (
            .O(N__10834),
            .I(N__10831));
    CascadeBuf I__1448 (
            .O(N__10831),
            .I(N__10828));
    CascadeMux I__1447 (
            .O(N__10828),
            .I(N__10824));
    CascadeMux I__1446 (
            .O(N__10827),
            .I(N__10821));
    CascadeBuf I__1445 (
            .O(N__10824),
            .I(N__10818));
    CascadeBuf I__1444 (
            .O(N__10821),
            .I(N__10815));
    CascadeMux I__1443 (
            .O(N__10818),
            .I(N__10812));
    CascadeMux I__1442 (
            .O(N__10815),
            .I(N__10809));
    CascadeBuf I__1441 (
            .O(N__10812),
            .I(N__10806));
    CascadeBuf I__1440 (
            .O(N__10809),
            .I(N__10803));
    CascadeMux I__1439 (
            .O(N__10806),
            .I(N__10800));
    CascadeMux I__1438 (
            .O(N__10803),
            .I(N__10797));
    CascadeBuf I__1437 (
            .O(N__10800),
            .I(N__10794));
    CascadeBuf I__1436 (
            .O(N__10797),
            .I(N__10791));
    CascadeMux I__1435 (
            .O(N__10794),
            .I(N__10788));
    CascadeMux I__1434 (
            .O(N__10791),
            .I(N__10785));
    CascadeBuf I__1433 (
            .O(N__10788),
            .I(N__10782));
    CascadeBuf I__1432 (
            .O(N__10785),
            .I(N__10779));
    CascadeMux I__1431 (
            .O(N__10782),
            .I(N__10776));
    CascadeMux I__1430 (
            .O(N__10779),
            .I(N__10773));
    CascadeBuf I__1429 (
            .O(N__10776),
            .I(N__10770));
    CascadeBuf I__1428 (
            .O(N__10773),
            .I(N__10767));
    CascadeMux I__1427 (
            .O(N__10770),
            .I(N__10764));
    CascadeMux I__1426 (
            .O(N__10767),
            .I(N__10761));
    CascadeBuf I__1425 (
            .O(N__10764),
            .I(N__10758));
    CascadeBuf I__1424 (
            .O(N__10761),
            .I(N__10755));
    CascadeMux I__1423 (
            .O(N__10758),
            .I(N__10752));
    CascadeMux I__1422 (
            .O(N__10755),
            .I(N__10749));
    CascadeBuf I__1421 (
            .O(N__10752),
            .I(N__10746));
    CascadeBuf I__1420 (
            .O(N__10749),
            .I(N__10743));
    CascadeMux I__1419 (
            .O(N__10746),
            .I(N__10740));
    CascadeMux I__1418 (
            .O(N__10743),
            .I(N__10737));
    CascadeBuf I__1417 (
            .O(N__10740),
            .I(N__10734));
    CascadeBuf I__1416 (
            .O(N__10737),
            .I(N__10731));
    CascadeMux I__1415 (
            .O(N__10734),
            .I(N__10728));
    CascadeMux I__1414 (
            .O(N__10731),
            .I(N__10725));
    CascadeBuf I__1413 (
            .O(N__10728),
            .I(N__10722));
    CascadeBuf I__1412 (
            .O(N__10725),
            .I(N__10719));
    CascadeMux I__1411 (
            .O(N__10722),
            .I(N__10716));
    CascadeMux I__1410 (
            .O(N__10719),
            .I(N__10713));
    CascadeBuf I__1409 (
            .O(N__10716),
            .I(N__10710));
    CascadeBuf I__1408 (
            .O(N__10713),
            .I(N__10707));
    CascadeMux I__1407 (
            .O(N__10710),
            .I(N__10704));
    CascadeMux I__1406 (
            .O(N__10707),
            .I(N__10701));
    CascadeBuf I__1405 (
            .O(N__10704),
            .I(N__10698));
    CascadeBuf I__1404 (
            .O(N__10701),
            .I(N__10695));
    CascadeMux I__1403 (
            .O(N__10698),
            .I(N__10692));
    CascadeMux I__1402 (
            .O(N__10695),
            .I(N__10689));
    CascadeBuf I__1401 (
            .O(N__10692),
            .I(N__10686));
    CascadeBuf I__1400 (
            .O(N__10689),
            .I(N__10683));
    CascadeMux I__1399 (
            .O(N__10686),
            .I(N__10680));
    CascadeMux I__1398 (
            .O(N__10683),
            .I(N__10677));
    CascadeBuf I__1397 (
            .O(N__10680),
            .I(N__10674));
    CascadeBuf I__1396 (
            .O(N__10677),
            .I(N__10671));
    CascadeMux I__1395 (
            .O(N__10674),
            .I(N__10668));
    CascadeMux I__1394 (
            .O(N__10671),
            .I(N__10665));
    CascadeBuf I__1393 (
            .O(N__10668),
            .I(N__10662));
    CascadeBuf I__1392 (
            .O(N__10665),
            .I(N__10659));
    CascadeMux I__1391 (
            .O(N__10662),
            .I(N__10656));
    CascadeMux I__1390 (
            .O(N__10659),
            .I(N__10653));
    InMux I__1389 (
            .O(N__10656),
            .I(N__10650));
    CascadeBuf I__1388 (
            .O(N__10653),
            .I(N__10647));
    LocalMux I__1387 (
            .O(N__10650),
            .I(N__10644));
    CascadeMux I__1386 (
            .O(N__10647),
            .I(N__10641));
    Span4Mux_s3_v I__1385 (
            .O(N__10644),
            .I(N__10638));
    InMux I__1384 (
            .O(N__10641),
            .I(N__10635));
    Span4Mux_h I__1383 (
            .O(N__10638),
            .I(N__10632));
    LocalMux I__1382 (
            .O(N__10635),
            .I(N__10629));
    Span4Mux_v I__1381 (
            .O(N__10632),
            .I(N__10626));
    Span12Mux_s7_v I__1380 (
            .O(N__10629),
            .I(N__10623));
    Sp12to4 I__1379 (
            .O(N__10626),
            .I(N__10618));
    Span12Mux_h I__1378 (
            .O(N__10623),
            .I(N__10618));
    Odrv12 I__1377 (
            .O(N__10618),
            .I(n24));
    CascadeMux I__1376 (
            .O(N__10615),
            .I(N__10610));
    InMux I__1375 (
            .O(N__10614),
            .I(N__10604));
    InMux I__1374 (
            .O(N__10613),
            .I(N__10604));
    InMux I__1373 (
            .O(N__10610),
            .I(N__10599));
    InMux I__1372 (
            .O(N__10609),
            .I(N__10599));
    LocalMux I__1371 (
            .O(N__10604),
            .I(\transmit_module.old_VGA_HS ));
    LocalMux I__1370 (
            .O(N__10599),
            .I(\transmit_module.old_VGA_HS ));
    CascadeMux I__1369 (
            .O(N__10594),
            .I(N__10591));
    InMux I__1368 (
            .O(N__10591),
            .I(N__10585));
    InMux I__1367 (
            .O(N__10590),
            .I(N__10585));
    LocalMux I__1366 (
            .O(N__10585),
            .I(N__10580));
    InMux I__1365 (
            .O(N__10584),
            .I(N__10575));
    InMux I__1364 (
            .O(N__10583),
            .I(N__10575));
    Odrv4 I__1363 (
            .O(N__10580),
            .I(\transmit_module.VGA_VISIBLE_Y ));
    LocalMux I__1362 (
            .O(N__10575),
            .I(\transmit_module.VGA_VISIBLE_Y ));
    IoInMux I__1361 (
            .O(N__10570),
            .I(N__10567));
    LocalMux I__1360 (
            .O(N__10567),
            .I(N__10564));
    IoSpan4Mux I__1359 (
            .O(N__10564),
            .I(N__10561));
    Span4Mux_s2_h I__1358 (
            .O(N__10561),
            .I(N__10558));
    Span4Mux_h I__1357 (
            .O(N__10558),
            .I(N__10553));
    InMux I__1356 (
            .O(N__10557),
            .I(N__10548));
    InMux I__1355 (
            .O(N__10556),
            .I(N__10548));
    Span4Mux_h I__1354 (
            .O(N__10553),
            .I(N__10542));
    LocalMux I__1353 (
            .O(N__10548),
            .I(N__10539));
    InMux I__1352 (
            .O(N__10547),
            .I(N__10532));
    InMux I__1351 (
            .O(N__10546),
            .I(N__10532));
    InMux I__1350 (
            .O(N__10545),
            .I(N__10532));
    Odrv4 I__1349 (
            .O(N__10542),
            .I(ADV_HSYNC_c));
    Odrv4 I__1348 (
            .O(N__10539),
            .I(ADV_HSYNC_c));
    LocalMux I__1347 (
            .O(N__10532),
            .I(ADV_HSYNC_c));
    InMux I__1346 (
            .O(N__10525),
            .I(N__10522));
    LocalMux I__1345 (
            .O(N__10522),
            .I(N__10518));
    InMux I__1344 (
            .O(N__10521),
            .I(N__10515));
    Odrv4 I__1343 (
            .O(N__10518),
            .I(\transmit_module.video_signal_controller.n3486 ));
    LocalMux I__1342 (
            .O(N__10515),
            .I(\transmit_module.video_signal_controller.n3486 ));
    InMux I__1341 (
            .O(N__10510),
            .I(N__10507));
    LocalMux I__1340 (
            .O(N__10507),
            .I(N__10504));
    Span4Mux_h I__1339 (
            .O(N__10504),
            .I(N__10501));
    Odrv4 I__1338 (
            .O(N__10501),
            .I(\transmit_module.video_signal_controller.n7 ));
    CascadeMux I__1337 (
            .O(N__10498),
            .I(N__10495));
    InMux I__1336 (
            .O(N__10495),
            .I(N__10492));
    LocalMux I__1335 (
            .O(N__10492),
            .I(N__10486));
    InMux I__1334 (
            .O(N__10491),
            .I(N__10480));
    InMux I__1333 (
            .O(N__10490),
            .I(N__10480));
    InMux I__1332 (
            .O(N__10489),
            .I(N__10477));
    Span4Mux_h I__1331 (
            .O(N__10486),
            .I(N__10474));
    InMux I__1330 (
            .O(N__10485),
            .I(N__10471));
    LocalMux I__1329 (
            .O(N__10480),
            .I(N__10468));
    LocalMux I__1328 (
            .O(N__10477),
            .I(\transmit_module.video_signal_controller.VGA_X_11 ));
    Odrv4 I__1327 (
            .O(N__10474),
            .I(\transmit_module.video_signal_controller.VGA_X_11 ));
    LocalMux I__1326 (
            .O(N__10471),
            .I(\transmit_module.video_signal_controller.VGA_X_11 ));
    Odrv4 I__1325 (
            .O(N__10468),
            .I(\transmit_module.video_signal_controller.VGA_X_11 ));
    InMux I__1324 (
            .O(N__10459),
            .I(N__10456));
    LocalMux I__1323 (
            .O(N__10456),
            .I(N__10452));
    InMux I__1322 (
            .O(N__10455),
            .I(N__10449));
    Odrv4 I__1321 (
            .O(N__10452),
            .I(\transmit_module.video_signal_controller.VGA_VISIBLE_N_578 ));
    LocalMux I__1320 (
            .O(N__10449),
            .I(\transmit_module.video_signal_controller.VGA_VISIBLE_N_578 ));
    CascadeMux I__1319 (
            .O(N__10444),
            .I(\transmit_module.n111_cascade_ ));
    CascadeMux I__1318 (
            .O(N__10441),
            .I(N__10438));
    CascadeBuf I__1317 (
            .O(N__10438),
            .I(N__10435));
    CascadeMux I__1316 (
            .O(N__10435),
            .I(N__10432));
    CascadeBuf I__1315 (
            .O(N__10432),
            .I(N__10428));
    CascadeMux I__1314 (
            .O(N__10431),
            .I(N__10425));
    CascadeMux I__1313 (
            .O(N__10428),
            .I(N__10422));
    CascadeBuf I__1312 (
            .O(N__10425),
            .I(N__10419));
    CascadeBuf I__1311 (
            .O(N__10422),
            .I(N__10416));
    CascadeMux I__1310 (
            .O(N__10419),
            .I(N__10413));
    CascadeMux I__1309 (
            .O(N__10416),
            .I(N__10410));
    CascadeBuf I__1308 (
            .O(N__10413),
            .I(N__10407));
    CascadeBuf I__1307 (
            .O(N__10410),
            .I(N__10404));
    CascadeMux I__1306 (
            .O(N__10407),
            .I(N__10401));
    CascadeMux I__1305 (
            .O(N__10404),
            .I(N__10398));
    CascadeBuf I__1304 (
            .O(N__10401),
            .I(N__10395));
    CascadeBuf I__1303 (
            .O(N__10398),
            .I(N__10392));
    CascadeMux I__1302 (
            .O(N__10395),
            .I(N__10389));
    CascadeMux I__1301 (
            .O(N__10392),
            .I(N__10386));
    CascadeBuf I__1300 (
            .O(N__10389),
            .I(N__10383));
    CascadeBuf I__1299 (
            .O(N__10386),
            .I(N__10380));
    CascadeMux I__1298 (
            .O(N__10383),
            .I(N__10377));
    CascadeMux I__1297 (
            .O(N__10380),
            .I(N__10374));
    CascadeBuf I__1296 (
            .O(N__10377),
            .I(N__10371));
    CascadeBuf I__1295 (
            .O(N__10374),
            .I(N__10368));
    CascadeMux I__1294 (
            .O(N__10371),
            .I(N__10365));
    CascadeMux I__1293 (
            .O(N__10368),
            .I(N__10362));
    CascadeBuf I__1292 (
            .O(N__10365),
            .I(N__10359));
    CascadeBuf I__1291 (
            .O(N__10362),
            .I(N__10356));
    CascadeMux I__1290 (
            .O(N__10359),
            .I(N__10353));
    CascadeMux I__1289 (
            .O(N__10356),
            .I(N__10350));
    CascadeBuf I__1288 (
            .O(N__10353),
            .I(N__10347));
    CascadeBuf I__1287 (
            .O(N__10350),
            .I(N__10344));
    CascadeMux I__1286 (
            .O(N__10347),
            .I(N__10341));
    CascadeMux I__1285 (
            .O(N__10344),
            .I(N__10338));
    CascadeBuf I__1284 (
            .O(N__10341),
            .I(N__10335));
    CascadeBuf I__1283 (
            .O(N__10338),
            .I(N__10332));
    CascadeMux I__1282 (
            .O(N__10335),
            .I(N__10329));
    CascadeMux I__1281 (
            .O(N__10332),
            .I(N__10326));
    CascadeBuf I__1280 (
            .O(N__10329),
            .I(N__10323));
    CascadeBuf I__1279 (
            .O(N__10326),
            .I(N__10320));
    CascadeMux I__1278 (
            .O(N__10323),
            .I(N__10317));
    CascadeMux I__1277 (
            .O(N__10320),
            .I(N__10314));
    CascadeBuf I__1276 (
            .O(N__10317),
            .I(N__10311));
    CascadeBuf I__1275 (
            .O(N__10314),
            .I(N__10308));
    CascadeMux I__1274 (
            .O(N__10311),
            .I(N__10305));
    CascadeMux I__1273 (
            .O(N__10308),
            .I(N__10302));
    CascadeBuf I__1272 (
            .O(N__10305),
            .I(N__10299));
    CascadeBuf I__1271 (
            .O(N__10302),
            .I(N__10296));
    CascadeMux I__1270 (
            .O(N__10299),
            .I(N__10293));
    CascadeMux I__1269 (
            .O(N__10296),
            .I(N__10290));
    CascadeBuf I__1268 (
            .O(N__10293),
            .I(N__10287));
    CascadeBuf I__1267 (
            .O(N__10290),
            .I(N__10284));
    CascadeMux I__1266 (
            .O(N__10287),
            .I(N__10281));
    CascadeMux I__1265 (
            .O(N__10284),
            .I(N__10278));
    CascadeBuf I__1264 (
            .O(N__10281),
            .I(N__10275));
    CascadeBuf I__1263 (
            .O(N__10278),
            .I(N__10272));
    CascadeMux I__1262 (
            .O(N__10275),
            .I(N__10269));
    CascadeMux I__1261 (
            .O(N__10272),
            .I(N__10266));
    CascadeBuf I__1260 (
            .O(N__10269),
            .I(N__10263));
    InMux I__1259 (
            .O(N__10266),
            .I(N__10260));
    CascadeMux I__1258 (
            .O(N__10263),
            .I(N__10257));
    LocalMux I__1257 (
            .O(N__10260),
            .I(N__10254));
    CascadeBuf I__1256 (
            .O(N__10257),
            .I(N__10251));
    Span4Mux_v I__1255 (
            .O(N__10254),
            .I(N__10248));
    CascadeMux I__1254 (
            .O(N__10251),
            .I(N__10245));
    Span4Mux_v I__1253 (
            .O(N__10248),
            .I(N__10242));
    InMux I__1252 (
            .O(N__10245),
            .I(N__10239));
    Span4Mux_v I__1251 (
            .O(N__10242),
            .I(N__10236));
    LocalMux I__1250 (
            .O(N__10239),
            .I(N__10233));
    Span4Mux_h I__1249 (
            .O(N__10236),
            .I(N__10230));
    Span4Mux_v I__1248 (
            .O(N__10233),
            .I(N__10227));
    Span4Mux_h I__1247 (
            .O(N__10230),
            .I(N__10224));
    Span4Mux_v I__1246 (
            .O(N__10227),
            .I(N__10221));
    Span4Mux_h I__1245 (
            .O(N__10224),
            .I(N__10216));
    Span4Mux_h I__1244 (
            .O(N__10221),
            .I(N__10216));
    Sp12to4 I__1243 (
            .O(N__10216),
            .I(N__10213));
    Odrv12 I__1242 (
            .O(N__10213),
            .I(n23));
    InMux I__1241 (
            .O(N__10210),
            .I(N__10207));
    LocalMux I__1240 (
            .O(N__10207),
            .I(\transmit_module.video_signal_controller.n8 ));
    CascadeMux I__1239 (
            .O(N__10204),
            .I(\transmit_module.video_signal_controller.n7_adj_615_cascade_ ));
    CascadeMux I__1238 (
            .O(N__10201),
            .I(\transmit_module.video_signal_controller.n2_cascade_ ));
    InMux I__1237 (
            .O(N__10198),
            .I(N__10195));
    LocalMux I__1236 (
            .O(N__10195),
            .I(\transmit_module.video_signal_controller.n3785 ));
    CascadeMux I__1235 (
            .O(N__10192),
            .I(\transmit_module.video_signal_controller.n3577_cascade_ ));
    InMux I__1234 (
            .O(N__10189),
            .I(N__10183));
    InMux I__1233 (
            .O(N__10188),
            .I(N__10183));
    LocalMux I__1232 (
            .O(N__10183),
            .I(\transmit_module.video_signal_controller.n3485 ));
    InMux I__1231 (
            .O(N__10180),
            .I(N__10172));
    InMux I__1230 (
            .O(N__10179),
            .I(N__10172));
    InMux I__1229 (
            .O(N__10178),
            .I(N__10169));
    InMux I__1228 (
            .O(N__10177),
            .I(N__10166));
    LocalMux I__1227 (
            .O(N__10172),
            .I(N__10163));
    LocalMux I__1226 (
            .O(N__10169),
            .I(\transmit_module.video_signal_controller.VGA_Y_9 ));
    LocalMux I__1225 (
            .O(N__10166),
            .I(\transmit_module.video_signal_controller.VGA_Y_9 ));
    Odrv4 I__1224 (
            .O(N__10163),
            .I(\transmit_module.video_signal_controller.VGA_Y_9 ));
    InMux I__1223 (
            .O(N__10156),
            .I(N__10150));
    InMux I__1222 (
            .O(N__10155),
            .I(N__10147));
    InMux I__1221 (
            .O(N__10154),
            .I(N__10142));
    InMux I__1220 (
            .O(N__10153),
            .I(N__10142));
    LocalMux I__1219 (
            .O(N__10150),
            .I(\transmit_module.video_signal_controller.VGA_Y_6 ));
    LocalMux I__1218 (
            .O(N__10147),
            .I(\transmit_module.video_signal_controller.VGA_Y_6 ));
    LocalMux I__1217 (
            .O(N__10142),
            .I(\transmit_module.video_signal_controller.VGA_Y_6 ));
    InMux I__1216 (
            .O(N__10135),
            .I(N__10130));
    InMux I__1215 (
            .O(N__10134),
            .I(N__10125));
    InMux I__1214 (
            .O(N__10133),
            .I(N__10125));
    LocalMux I__1213 (
            .O(N__10130),
            .I(\transmit_module.video_signal_controller.VGA_Y_11 ));
    LocalMux I__1212 (
            .O(N__10125),
            .I(\transmit_module.video_signal_controller.VGA_Y_11 ));
    InMux I__1211 (
            .O(N__10120),
            .I(N__10114));
    InMux I__1210 (
            .O(N__10119),
            .I(N__10111));
    InMux I__1209 (
            .O(N__10118),
            .I(N__10106));
    InMux I__1208 (
            .O(N__10117),
            .I(N__10106));
    LocalMux I__1207 (
            .O(N__10114),
            .I(\transmit_module.video_signal_controller.VGA_Y_7 ));
    LocalMux I__1206 (
            .O(N__10111),
            .I(\transmit_module.video_signal_controller.VGA_Y_7 ));
    LocalMux I__1205 (
            .O(N__10106),
            .I(\transmit_module.video_signal_controller.VGA_Y_7 ));
    CascadeMux I__1204 (
            .O(N__10099),
            .I(N__10096));
    InMux I__1203 (
            .O(N__10096),
            .I(N__10090));
    InMux I__1202 (
            .O(N__10095),
            .I(N__10087));
    InMux I__1201 (
            .O(N__10094),
            .I(N__10082));
    InMux I__1200 (
            .O(N__10093),
            .I(N__10082));
    LocalMux I__1199 (
            .O(N__10090),
            .I(\transmit_module.video_signal_controller.VGA_Y_5 ));
    LocalMux I__1198 (
            .O(N__10087),
            .I(\transmit_module.video_signal_controller.VGA_Y_5 ));
    LocalMux I__1197 (
            .O(N__10082),
            .I(\transmit_module.video_signal_controller.VGA_Y_5 ));
    InMux I__1196 (
            .O(N__10075),
            .I(N__10069));
    InMux I__1195 (
            .O(N__10074),
            .I(N__10066));
    InMux I__1194 (
            .O(N__10073),
            .I(N__10061));
    InMux I__1193 (
            .O(N__10072),
            .I(N__10061));
    LocalMux I__1192 (
            .O(N__10069),
            .I(\transmit_module.video_signal_controller.VGA_Y_2 ));
    LocalMux I__1191 (
            .O(N__10066),
            .I(\transmit_module.video_signal_controller.VGA_Y_2 ));
    LocalMux I__1190 (
            .O(N__10061),
            .I(\transmit_module.video_signal_controller.VGA_Y_2 ));
    CEMux I__1189 (
            .O(N__10054),
            .I(N__10046));
    CEMux I__1188 (
            .O(N__10053),
            .I(N__10043));
    CEMux I__1187 (
            .O(N__10052),
            .I(N__10040));
    CEMux I__1186 (
            .O(N__10051),
            .I(N__10036));
    CEMux I__1185 (
            .O(N__10050),
            .I(N__10032));
    CEMux I__1184 (
            .O(N__10049),
            .I(N__10029));
    LocalMux I__1183 (
            .O(N__10046),
            .I(N__10025));
    LocalMux I__1182 (
            .O(N__10043),
            .I(N__10021));
    LocalMux I__1181 (
            .O(N__10040),
            .I(N__10018));
    CEMux I__1180 (
            .O(N__10039),
            .I(N__10015));
    LocalMux I__1179 (
            .O(N__10036),
            .I(N__10012));
    CEMux I__1178 (
            .O(N__10035),
            .I(N__10009));
    LocalMux I__1177 (
            .O(N__10032),
            .I(N__10006));
    LocalMux I__1176 (
            .O(N__10029),
            .I(N__10003));
    CEMux I__1175 (
            .O(N__10028),
            .I(N__10000));
    Span4Mux_h I__1174 (
            .O(N__10025),
            .I(N__9997));
    CEMux I__1173 (
            .O(N__10024),
            .I(N__9994));
    Span4Mux_v I__1172 (
            .O(N__10021),
            .I(N__9989));
    Span4Mux_v I__1171 (
            .O(N__10018),
            .I(N__9989));
    LocalMux I__1170 (
            .O(N__10015),
            .I(N__9986));
    Span4Mux_v I__1169 (
            .O(N__10012),
            .I(N__9981));
    LocalMux I__1168 (
            .O(N__10009),
            .I(N__9981));
    Span4Mux_v I__1167 (
            .O(N__10006),
            .I(N__9976));
    Span4Mux_h I__1166 (
            .O(N__10003),
            .I(N__9976));
    LocalMux I__1165 (
            .O(N__10000),
            .I(N__9973));
    Span4Mux_h I__1164 (
            .O(N__9997),
            .I(N__9968));
    LocalMux I__1163 (
            .O(N__9994),
            .I(N__9968));
    Span4Mux_v I__1162 (
            .O(N__9989),
            .I(N__9965));
    Span12Mux_h I__1161 (
            .O(N__9986),
            .I(N__9962));
    Span4Mux_h I__1160 (
            .O(N__9981),
            .I(N__9959));
    Span4Mux_h I__1159 (
            .O(N__9976),
            .I(N__9954));
    Span4Mux_h I__1158 (
            .O(N__9973),
            .I(N__9954));
    Span4Mux_h I__1157 (
            .O(N__9968),
            .I(N__9951));
    Odrv4 I__1156 (
            .O(N__9965),
            .I(\transmit_module.n3798 ));
    Odrv12 I__1155 (
            .O(N__9962),
            .I(\transmit_module.n3798 ));
    Odrv4 I__1154 (
            .O(N__9959),
            .I(\transmit_module.n3798 ));
    Odrv4 I__1153 (
            .O(N__9954),
            .I(\transmit_module.n3798 ));
    Odrv4 I__1152 (
            .O(N__9951),
            .I(\transmit_module.n3798 ));
    InMux I__1151 (
            .O(N__9940),
            .I(\receive_module.rx_counter.n3275 ));
    InMux I__1150 (
            .O(N__9937),
            .I(\receive_module.rx_counter.n3276 ));
    InMux I__1149 (
            .O(N__9934),
            .I(\receive_module.rx_counter.n3277 ));
    InMux I__1148 (
            .O(N__9931),
            .I(bfn_13_11_0_));
    CascadeMux I__1147 (
            .O(N__9928),
            .I(\transmit_module.video_signal_controller.n3786_cascade_ ));
    InMux I__1146 (
            .O(N__9925),
            .I(N__9922));
    LocalMux I__1145 (
            .O(N__9922),
            .I(\transmit_module.Y_DELTA_PATTERN_4 ));
    InMux I__1144 (
            .O(N__9919),
            .I(N__9916));
    LocalMux I__1143 (
            .O(N__9916),
            .I(\transmit_module.Y_DELTA_PATTERN_3 ));
    InMux I__1142 (
            .O(N__9913),
            .I(N__9910));
    LocalMux I__1141 (
            .O(N__9910),
            .I(N__9907));
    Span12Mux_v I__1140 (
            .O(N__9907),
            .I(N__9904));
    Odrv12 I__1139 (
            .O(N__9904),
            .I(\line_buffer.n578 ));
    InMux I__1138 (
            .O(N__9901),
            .I(N__9898));
    LocalMux I__1137 (
            .O(N__9898),
            .I(N__9895));
    Span4Mux_h I__1136 (
            .O(N__9895),
            .I(N__9892));
    Odrv4 I__1135 (
            .O(N__9892),
            .I(\line_buffer.n570 ));
    InMux I__1134 (
            .O(N__9889),
            .I(N__9886));
    LocalMux I__1133 (
            .O(N__9886),
            .I(N__9883));
    Span12Mux_v I__1132 (
            .O(N__9883),
            .I(N__9880));
    Odrv12 I__1131 (
            .O(N__9880),
            .I(\line_buffer.n577 ));
    InMux I__1130 (
            .O(N__9877),
            .I(N__9874));
    LocalMux I__1129 (
            .O(N__9874),
            .I(N__9871));
    Span12Mux_v I__1128 (
            .O(N__9871),
            .I(N__9868));
    Odrv12 I__1127 (
            .O(N__9868),
            .I(\line_buffer.n569 ));
    InMux I__1126 (
            .O(N__9865),
            .I(bfn_13_10_0_));
    InMux I__1125 (
            .O(N__9862),
            .I(\receive_module.rx_counter.n3271 ));
    InMux I__1124 (
            .O(N__9859),
            .I(\receive_module.rx_counter.n3272 ));
    InMux I__1123 (
            .O(N__9856),
            .I(\receive_module.rx_counter.n3273 ));
    InMux I__1122 (
            .O(N__9853),
            .I(\receive_module.rx_counter.n3274 ));
    SRMux I__1121 (
            .O(N__9850),
            .I(N__9846));
    SRMux I__1120 (
            .O(N__9849),
            .I(N__9843));
    LocalMux I__1119 (
            .O(N__9846),
            .I(\transmit_module.video_signal_controller.n2361 ));
    LocalMux I__1118 (
            .O(N__9843),
            .I(\transmit_module.video_signal_controller.n2361 ));
    CascadeMux I__1117 (
            .O(N__9838),
            .I(\transmit_module.n3787_cascade_ ));
    InMux I__1116 (
            .O(N__9835),
            .I(N__9832));
    LocalMux I__1115 (
            .O(N__9832),
            .I(\transmit_module.Y_DELTA_PATTERN_7 ));
    InMux I__1114 (
            .O(N__9829),
            .I(N__9826));
    LocalMux I__1113 (
            .O(N__9826),
            .I(\transmit_module.Y_DELTA_PATTERN_6 ));
    InMux I__1112 (
            .O(N__9823),
            .I(N__9820));
    LocalMux I__1111 (
            .O(N__9820),
            .I(\transmit_module.Y_DELTA_PATTERN_5 ));
    InMux I__1110 (
            .O(N__9817),
            .I(\transmit_module.video_signal_controller.n3292 ));
    InMux I__1109 (
            .O(N__9814),
            .I(\transmit_module.video_signal_controller.n3293 ));
    InMux I__1108 (
            .O(N__9811),
            .I(\transmit_module.video_signal_controller.n3294 ));
    InMux I__1107 (
            .O(N__9808),
            .I(\transmit_module.video_signal_controller.n3295 ));
    InMux I__1106 (
            .O(N__9805),
            .I(\transmit_module.video_signal_controller.n3296 ));
    InMux I__1105 (
            .O(N__9802),
            .I(bfn_12_14_0_));
    InMux I__1104 (
            .O(N__9799),
            .I(\transmit_module.video_signal_controller.n3298 ));
    InMux I__1103 (
            .O(N__9796),
            .I(\transmit_module.video_signal_controller.n3299 ));
    InMux I__1102 (
            .O(N__9793),
            .I(\transmit_module.video_signal_controller.n3300 ));
    SRMux I__1101 (
            .O(N__9790),
            .I(N__9787));
    LocalMux I__1100 (
            .O(N__9787),
            .I(N__9783));
    SRMux I__1099 (
            .O(N__9786),
            .I(N__9779));
    Span4Mux_v I__1098 (
            .O(N__9783),
            .I(N__9775));
    CEMux I__1097 (
            .O(N__9782),
            .I(N__9772));
    LocalMux I__1096 (
            .O(N__9779),
            .I(N__9769));
    CEMux I__1095 (
            .O(N__9778),
            .I(N__9766));
    Span4Mux_h I__1094 (
            .O(N__9775),
            .I(N__9759));
    LocalMux I__1093 (
            .O(N__9772),
            .I(N__9759));
    Span4Mux_v I__1092 (
            .O(N__9769),
            .I(N__9759));
    LocalMux I__1091 (
            .O(N__9766),
            .I(\transmit_module.video_signal_controller.n2010 ));
    Odrv4 I__1090 (
            .O(N__9759),
            .I(\transmit_module.video_signal_controller.n2010 ));
    InMux I__1089 (
            .O(N__9754),
            .I(N__9751));
    LocalMux I__1088 (
            .O(N__9751),
            .I(\transmit_module.Y_DELTA_PATTERN_60 ));
    InMux I__1087 (
            .O(N__9748),
            .I(N__9745));
    LocalMux I__1086 (
            .O(N__9745),
            .I(\transmit_module.Y_DELTA_PATTERN_59 ));
    InMux I__1085 (
            .O(N__9742),
            .I(N__9739));
    LocalMux I__1084 (
            .O(N__9739),
            .I(\transmit_module.Y_DELTA_PATTERN_98 ));
    InMux I__1083 (
            .O(N__9736),
            .I(N__9733));
    LocalMux I__1082 (
            .O(N__9733),
            .I(N__9730));
    Odrv4 I__1081 (
            .O(N__9730),
            .I(\transmit_module.Y_DELTA_PATTERN_86 ));
    InMux I__1080 (
            .O(N__9727),
            .I(N__9724));
    LocalMux I__1079 (
            .O(N__9724),
            .I(\transmit_module.Y_DELTA_PATTERN_85 ));
    InMux I__1078 (
            .O(N__9721),
            .I(N__9718));
    LocalMux I__1077 (
            .O(N__9718),
            .I(\transmit_module.Y_DELTA_PATTERN_84 ));
    InMux I__1076 (
            .O(N__9715),
            .I(N__9712));
    LocalMux I__1075 (
            .O(N__9712),
            .I(\transmit_module.Y_DELTA_PATTERN_83 ));
    InMux I__1074 (
            .O(N__9709),
            .I(N__9706));
    LocalMux I__1073 (
            .O(N__9706),
            .I(\transmit_module.Y_DELTA_PATTERN_99 ));
    InMux I__1072 (
            .O(N__9703),
            .I(bfn_12_13_0_));
    InMux I__1071 (
            .O(N__9700),
            .I(\transmit_module.video_signal_controller.n3290 ));
    InMux I__1070 (
            .O(N__9697),
            .I(\transmit_module.video_signal_controller.n3291 ));
    CascadeMux I__1069 (
            .O(N__9694),
            .I(N__9691));
    InMux I__1068 (
            .O(N__9691),
            .I(N__9683));
    InMux I__1067 (
            .O(N__9690),
            .I(N__9683));
    InMux I__1066 (
            .O(N__9689),
            .I(N__9680));
    InMux I__1065 (
            .O(N__9688),
            .I(N__9677));
    LocalMux I__1064 (
            .O(N__9683),
            .I(N__9674));
    LocalMux I__1063 (
            .O(N__9680),
            .I(\transmit_module.video_signal_controller.VGA_X_8 ));
    LocalMux I__1062 (
            .O(N__9677),
            .I(\transmit_module.video_signal_controller.VGA_X_8 ));
    Odrv4 I__1061 (
            .O(N__9674),
            .I(\transmit_module.video_signal_controller.VGA_X_8 ));
    CascadeMux I__1060 (
            .O(N__9667),
            .I(\transmit_module.video_signal_controller.n4_adj_617_cascade_ ));
    InMux I__1059 (
            .O(N__9664),
            .I(N__9658));
    InMux I__1058 (
            .O(N__9663),
            .I(N__9655));
    InMux I__1057 (
            .O(N__9662),
            .I(N__9652));
    InMux I__1056 (
            .O(N__9661),
            .I(N__9649));
    LocalMux I__1055 (
            .O(N__9658),
            .I(\transmit_module.video_signal_controller.VGA_X_6 ));
    LocalMux I__1054 (
            .O(N__9655),
            .I(\transmit_module.video_signal_controller.VGA_X_6 ));
    LocalMux I__1053 (
            .O(N__9652),
            .I(\transmit_module.video_signal_controller.VGA_X_6 ));
    LocalMux I__1052 (
            .O(N__9649),
            .I(\transmit_module.video_signal_controller.VGA_X_6 ));
    CascadeMux I__1051 (
            .O(N__9640),
            .I(N__9636));
    InMux I__1050 (
            .O(N__9639),
            .I(N__9630));
    InMux I__1049 (
            .O(N__9636),
            .I(N__9630));
    InMux I__1048 (
            .O(N__9635),
            .I(N__9626));
    LocalMux I__1047 (
            .O(N__9630),
            .I(N__9623));
    InMux I__1046 (
            .O(N__9629),
            .I(N__9620));
    LocalMux I__1045 (
            .O(N__9626),
            .I(\transmit_module.video_signal_controller.VGA_X_9 ));
    Odrv4 I__1044 (
            .O(N__9623),
            .I(\transmit_module.video_signal_controller.VGA_X_9 ));
    LocalMux I__1043 (
            .O(N__9620),
            .I(\transmit_module.video_signal_controller.VGA_X_9 ));
    InMux I__1042 (
            .O(N__9613),
            .I(N__9607));
    InMux I__1041 (
            .O(N__9612),
            .I(N__9607));
    LocalMux I__1040 (
            .O(N__9607),
            .I(N__9603));
    InMux I__1039 (
            .O(N__9606),
            .I(N__9599));
    Span4Mux_v I__1038 (
            .O(N__9603),
            .I(N__9596));
    InMux I__1037 (
            .O(N__9602),
            .I(N__9593));
    LocalMux I__1036 (
            .O(N__9599),
            .I(\transmit_module.video_signal_controller.VGA_X_10 ));
    Odrv4 I__1035 (
            .O(N__9596),
            .I(\transmit_module.video_signal_controller.VGA_X_10 ));
    LocalMux I__1034 (
            .O(N__9593),
            .I(\transmit_module.video_signal_controller.VGA_X_10 ));
    InMux I__1033 (
            .O(N__9586),
            .I(N__9583));
    LocalMux I__1032 (
            .O(N__9583),
            .I(\transmit_module.video_signal_controller.n4 ));
    CascadeMux I__1031 (
            .O(N__9580),
            .I(N__9577));
    InMux I__1030 (
            .O(N__9577),
            .I(N__9569));
    InMux I__1029 (
            .O(N__9576),
            .I(N__9569));
    InMux I__1028 (
            .O(N__9575),
            .I(N__9566));
    InMux I__1027 (
            .O(N__9574),
            .I(N__9563));
    LocalMux I__1026 (
            .O(N__9569),
            .I(\transmit_module.video_signal_controller.VGA_X_7 ));
    LocalMux I__1025 (
            .O(N__9566),
            .I(\transmit_module.video_signal_controller.VGA_X_7 ));
    LocalMux I__1024 (
            .O(N__9563),
            .I(\transmit_module.video_signal_controller.VGA_X_7 ));
    CascadeMux I__1023 (
            .O(N__9556),
            .I(\transmit_module.video_signal_controller.n3794_cascade_ ));
    InMux I__1022 (
            .O(N__9553),
            .I(N__9545));
    InMux I__1021 (
            .O(N__9552),
            .I(N__9545));
    InMux I__1020 (
            .O(N__9551),
            .I(N__9542));
    InMux I__1019 (
            .O(N__9550),
            .I(N__9539));
    LocalMux I__1018 (
            .O(N__9545),
            .I(\transmit_module.video_signal_controller.VGA_X_4 ));
    LocalMux I__1017 (
            .O(N__9542),
            .I(\transmit_module.video_signal_controller.VGA_X_4 ));
    LocalMux I__1016 (
            .O(N__9539),
            .I(\transmit_module.video_signal_controller.VGA_X_4 ));
    InMux I__1015 (
            .O(N__9532),
            .I(N__9529));
    LocalMux I__1014 (
            .O(N__9529),
            .I(\transmit_module.video_signal_controller.n3618 ));
    InMux I__1013 (
            .O(N__9526),
            .I(N__9523));
    LocalMux I__1012 (
            .O(N__9523),
            .I(\transmit_module.Y_DELTA_PATTERN_61 ));
    InMux I__1011 (
            .O(N__9520),
            .I(N__9517));
    LocalMux I__1010 (
            .O(N__9517),
            .I(\transmit_module.Y_DELTA_PATTERN_37 ));
    InMux I__1009 (
            .O(N__9514),
            .I(N__9511));
    LocalMux I__1008 (
            .O(N__9511),
            .I(\transmit_module.Y_DELTA_PATTERN_39 ));
    InMux I__1007 (
            .O(N__9508),
            .I(N__9505));
    LocalMux I__1006 (
            .O(N__9505),
            .I(\transmit_module.Y_DELTA_PATTERN_38 ));
    InMux I__1005 (
            .O(N__9502),
            .I(N__9499));
    LocalMux I__1004 (
            .O(N__9499),
            .I(\transmit_module.Y_DELTA_PATTERN_58 ));
    InMux I__1003 (
            .O(N__9496),
            .I(N__9493));
    LocalMux I__1002 (
            .O(N__9493),
            .I(\transmit_module.Y_DELTA_PATTERN_57 ));
    InMux I__1001 (
            .O(N__9490),
            .I(N__9487));
    LocalMux I__1000 (
            .O(N__9487),
            .I(\transmit_module.Y_DELTA_PATTERN_71 ));
    InMux I__999 (
            .O(N__9484),
            .I(N__9481));
    LocalMux I__998 (
            .O(N__9481),
            .I(\transmit_module.Y_DELTA_PATTERN_70 ));
    InMux I__997 (
            .O(N__9478),
            .I(N__9475));
    LocalMux I__996 (
            .O(N__9475),
            .I(\transmit_module.Y_DELTA_PATTERN_68 ));
    InMux I__995 (
            .O(N__9472),
            .I(N__9469));
    LocalMux I__994 (
            .O(N__9469),
            .I(N__9466));
    Odrv4 I__993 (
            .O(N__9466),
            .I(\transmit_module.Y_DELTA_PATTERN_67 ));
    InMux I__992 (
            .O(N__9463),
            .I(N__9460));
    LocalMux I__991 (
            .O(N__9460),
            .I(\transmit_module.video_signal_controller.n2886 ));
    CascadeMux I__990 (
            .O(N__9457),
            .I(\transmit_module.video_signal_controller.n1983_cascade_ ));
    InMux I__989 (
            .O(N__9454),
            .I(N__9451));
    LocalMux I__988 (
            .O(N__9451),
            .I(\transmit_module.video_signal_controller.n2926 ));
    CascadeMux I__987 (
            .O(N__9448),
            .I(\transmit_module.video_signal_controller.n2010_cascade_ ));
    InMux I__986 (
            .O(N__9445),
            .I(N__9442));
    LocalMux I__985 (
            .O(N__9442),
            .I(\transmit_module.video_signal_controller.n1983 ));
    InMux I__984 (
            .O(N__9439),
            .I(N__9436));
    LocalMux I__983 (
            .O(N__9436),
            .I(\transmit_module.video_signal_controller.n3789 ));
    InMux I__982 (
            .O(N__9433),
            .I(N__9427));
    InMux I__981 (
            .O(N__9432),
            .I(N__9427));
    LocalMux I__980 (
            .O(N__9427),
            .I(\transmit_module.video_signal_controller.n3467 ));
    CascadeMux I__979 (
            .O(N__9424),
            .I(\transmit_module.video_signal_controller.n18_cascade_ ));
    InMux I__978 (
            .O(N__9421),
            .I(N__9416));
    InMux I__977 (
            .O(N__9420),
            .I(N__9412));
    InMux I__976 (
            .O(N__9419),
            .I(N__9409));
    LocalMux I__975 (
            .O(N__9416),
            .I(N__9406));
    InMux I__974 (
            .O(N__9415),
            .I(N__9403));
    LocalMux I__973 (
            .O(N__9412),
            .I(\transmit_module.video_signal_controller.VGA_X_3 ));
    LocalMux I__972 (
            .O(N__9409),
            .I(\transmit_module.video_signal_controller.VGA_X_3 ));
    Odrv4 I__971 (
            .O(N__9406),
            .I(\transmit_module.video_signal_controller.VGA_X_3 ));
    LocalMux I__970 (
            .O(N__9403),
            .I(\transmit_module.video_signal_controller.VGA_X_3 ));
    InMux I__969 (
            .O(N__9394),
            .I(N__9388));
    InMux I__968 (
            .O(N__9393),
            .I(N__9385));
    InMux I__967 (
            .O(N__9392),
            .I(N__9382));
    InMux I__966 (
            .O(N__9391),
            .I(N__9379));
    LocalMux I__965 (
            .O(N__9388),
            .I(\transmit_module.video_signal_controller.VGA_X_5 ));
    LocalMux I__964 (
            .O(N__9385),
            .I(\transmit_module.video_signal_controller.VGA_X_5 ));
    LocalMux I__963 (
            .O(N__9382),
            .I(\transmit_module.video_signal_controller.VGA_X_5 ));
    LocalMux I__962 (
            .O(N__9379),
            .I(\transmit_module.video_signal_controller.VGA_X_5 ));
    InMux I__961 (
            .O(N__9370),
            .I(N__9367));
    LocalMux I__960 (
            .O(N__9367),
            .I(\transmit_module.Y_DELTA_PATTERN_81 ));
    InMux I__959 (
            .O(N__9364),
            .I(N__9361));
    LocalMux I__958 (
            .O(N__9361),
            .I(\transmit_module.Y_DELTA_PATTERN_50 ));
    InMux I__957 (
            .O(N__9358),
            .I(N__9355));
    LocalMux I__956 (
            .O(N__9355),
            .I(\transmit_module.Y_DELTA_PATTERN_49 ));
    InMux I__955 (
            .O(N__9352),
            .I(N__9349));
    LocalMux I__954 (
            .O(N__9349),
            .I(N__9346));
    Odrv4 I__953 (
            .O(N__9346),
            .I(\transmit_module.Y_DELTA_PATTERN_35 ));
    InMux I__952 (
            .O(N__9343),
            .I(N__9340));
    LocalMux I__951 (
            .O(N__9340),
            .I(\transmit_module.Y_DELTA_PATTERN_34 ));
    InMux I__950 (
            .O(N__9337),
            .I(N__9334));
    LocalMux I__949 (
            .O(N__9334),
            .I(\transmit_module.Y_DELTA_PATTERN_72 ));
    InMux I__948 (
            .O(N__9331),
            .I(N__9328));
    LocalMux I__947 (
            .O(N__9328),
            .I(\transmit_module.Y_DELTA_PATTERN_82 ));
    InMux I__946 (
            .O(N__9325),
            .I(N__9322));
    LocalMux I__945 (
            .O(N__9322),
            .I(\transmit_module.Y_DELTA_PATTERN_69 ));
    InMux I__944 (
            .O(N__9319),
            .I(N__9316));
    LocalMux I__943 (
            .O(N__9316),
            .I(N__9313));
    Span4Mux_h I__942 (
            .O(N__9313),
            .I(N__9310));
    Odrv4 I__941 (
            .O(N__9310),
            .I(\transmit_module.Y_DELTA_PATTERN_78 ));
    InMux I__940 (
            .O(N__9307),
            .I(N__9304));
    LocalMux I__939 (
            .O(N__9304),
            .I(\transmit_module.Y_DELTA_PATTERN_80 ));
    InMux I__938 (
            .O(N__9301),
            .I(N__9298));
    LocalMux I__937 (
            .O(N__9298),
            .I(\transmit_module.Y_DELTA_PATTERN_79 ));
    InMux I__936 (
            .O(N__9295),
            .I(N__9292));
    LocalMux I__935 (
            .O(N__9292),
            .I(\transmit_module.Y_DELTA_PATTERN_36 ));
    InMux I__934 (
            .O(N__9289),
            .I(N__9286));
    LocalMux I__933 (
            .O(N__9286),
            .I(\transmit_module.Y_DELTA_PATTERN_62 ));
    InMux I__932 (
            .O(N__9283),
            .I(N__9280));
    LocalMux I__931 (
            .O(N__9280),
            .I(\transmit_module.Y_DELTA_PATTERN_66 ));
    InMux I__930 (
            .O(N__9277),
            .I(N__9274));
    LocalMux I__929 (
            .O(N__9274),
            .I(N__9271));
    Odrv12 I__928 (
            .O(N__9271),
            .I(\transmit_module.Y_DELTA_PATTERN_53 ));
    InMux I__927 (
            .O(N__9268),
            .I(N__9265));
    LocalMux I__926 (
            .O(N__9265),
            .I(\transmit_module.Y_DELTA_PATTERN_52 ));
    InMux I__925 (
            .O(N__9262),
            .I(N__9259));
    LocalMux I__924 (
            .O(N__9259),
            .I(\transmit_module.Y_DELTA_PATTERN_51 ));
    InMux I__923 (
            .O(N__9256),
            .I(bfn_10_16_0_));
    InMux I__922 (
            .O(N__9253),
            .I(\transmit_module.video_signal_controller.n3287 ));
    InMux I__921 (
            .O(N__9250),
            .I(\transmit_module.video_signal_controller.n3288 ));
    InMux I__920 (
            .O(N__9247),
            .I(\transmit_module.video_signal_controller.n3289 ));
    InMux I__919 (
            .O(N__9244),
            .I(N__9241));
    LocalMux I__918 (
            .O(N__9241),
            .I(\transmit_module.Y_DELTA_PATTERN_55 ));
    InMux I__917 (
            .O(N__9238),
            .I(N__9235));
    LocalMux I__916 (
            .O(N__9235),
            .I(\transmit_module.Y_DELTA_PATTERN_54 ));
    InMux I__915 (
            .O(N__9232),
            .I(N__9229));
    LocalMux I__914 (
            .O(N__9229),
            .I(\transmit_module.Y_DELTA_PATTERN_40 ));
    InMux I__913 (
            .O(N__9226),
            .I(N__9223));
    LocalMux I__912 (
            .O(N__9223),
            .I(\transmit_module.Y_DELTA_PATTERN_56 ));
    InMux I__911 (
            .O(N__9220),
            .I(N__9217));
    LocalMux I__910 (
            .O(N__9217),
            .I(N__9214));
    Span4Mux_h I__909 (
            .O(N__9214),
            .I(N__9211));
    Odrv4 I__908 (
            .O(N__9211),
            .I(\transmit_module.Y_DELTA_PATTERN_97 ));
    InMux I__907 (
            .O(N__9208),
            .I(N__9203));
    InMux I__906 (
            .O(N__9207),
            .I(N__9198));
    InMux I__905 (
            .O(N__9206),
            .I(N__9198));
    LocalMux I__904 (
            .O(N__9203),
            .I(\transmit_module.video_signal_controller.VGA_X_0 ));
    LocalMux I__903 (
            .O(N__9198),
            .I(\transmit_module.video_signal_controller.VGA_X_0 ));
    InMux I__902 (
            .O(N__9193),
            .I(bfn_10_15_0_));
    CascadeMux I__901 (
            .O(N__9190),
            .I(N__9184));
    InMux I__900 (
            .O(N__9189),
            .I(N__9181));
    InMux I__899 (
            .O(N__9188),
            .I(N__9174));
    InMux I__898 (
            .O(N__9187),
            .I(N__9174));
    InMux I__897 (
            .O(N__9184),
            .I(N__9174));
    LocalMux I__896 (
            .O(N__9181),
            .I(\transmit_module.video_signal_controller.VGA_X_1 ));
    LocalMux I__895 (
            .O(N__9174),
            .I(\transmit_module.video_signal_controller.VGA_X_1 ));
    InMux I__894 (
            .O(N__9169),
            .I(\transmit_module.video_signal_controller.n3279 ));
    InMux I__893 (
            .O(N__9166),
            .I(N__9160));
    InMux I__892 (
            .O(N__9165),
            .I(N__9153));
    InMux I__891 (
            .O(N__9164),
            .I(N__9153));
    InMux I__890 (
            .O(N__9163),
            .I(N__9153));
    LocalMux I__889 (
            .O(N__9160),
            .I(\transmit_module.video_signal_controller.VGA_X_2 ));
    LocalMux I__888 (
            .O(N__9153),
            .I(\transmit_module.video_signal_controller.VGA_X_2 ));
    InMux I__887 (
            .O(N__9148),
            .I(\transmit_module.video_signal_controller.n3280 ));
    InMux I__886 (
            .O(N__9145),
            .I(\transmit_module.video_signal_controller.n3281 ));
    InMux I__885 (
            .O(N__9142),
            .I(\transmit_module.video_signal_controller.n3282 ));
    InMux I__884 (
            .O(N__9139),
            .I(\transmit_module.video_signal_controller.n3283 ));
    InMux I__883 (
            .O(N__9136),
            .I(\transmit_module.video_signal_controller.n3284 ));
    InMux I__882 (
            .O(N__9133),
            .I(\transmit_module.video_signal_controller.n3285 ));
    InMux I__881 (
            .O(N__9130),
            .I(N__9127));
    LocalMux I__880 (
            .O(N__9127),
            .I(N__9124));
    Odrv4 I__879 (
            .O(N__9124),
            .I(\transmit_module.Y_DELTA_PATTERN_42 ));
    InMux I__878 (
            .O(N__9121),
            .I(N__9118));
    LocalMux I__877 (
            .O(N__9118),
            .I(\transmit_module.Y_DELTA_PATTERN_96 ));
    InMux I__876 (
            .O(N__9115),
            .I(N__9112));
    LocalMux I__875 (
            .O(N__9112),
            .I(\transmit_module.Y_DELTA_PATTERN_45 ));
    InMux I__874 (
            .O(N__9109),
            .I(N__9106));
    LocalMux I__873 (
            .O(N__9106),
            .I(\transmit_module.Y_DELTA_PATTERN_44 ));
    InMux I__872 (
            .O(N__9103),
            .I(N__9100));
    LocalMux I__871 (
            .O(N__9100),
            .I(\transmit_module.Y_DELTA_PATTERN_43 ));
    CascadeMux I__870 (
            .O(N__9097),
            .I(\transmit_module.video_signal_controller.n3788_cascade_ ));
    InMux I__869 (
            .O(N__9094),
            .I(N__9091));
    LocalMux I__868 (
            .O(N__9091),
            .I(\transmit_module.video_signal_controller.n2876 ));
    InMux I__867 (
            .O(N__9088),
            .I(N__9085));
    LocalMux I__866 (
            .O(N__9085),
            .I(\transmit_module.Y_DELTA_PATTERN_63 ));
    InMux I__865 (
            .O(N__9082),
            .I(N__9079));
    LocalMux I__864 (
            .O(N__9079),
            .I(\transmit_module.Y_DELTA_PATTERN_74 ));
    InMux I__863 (
            .O(N__9076),
            .I(N__9073));
    LocalMux I__862 (
            .O(N__9073),
            .I(\transmit_module.Y_DELTA_PATTERN_76 ));
    InMux I__861 (
            .O(N__9070),
            .I(N__9067));
    LocalMux I__860 (
            .O(N__9067),
            .I(\transmit_module.Y_DELTA_PATTERN_75 ));
    InMux I__859 (
            .O(N__9064),
            .I(N__9061));
    LocalMux I__858 (
            .O(N__9061),
            .I(\transmit_module.Y_DELTA_PATTERN_73 ));
    InMux I__857 (
            .O(N__9058),
            .I(N__9055));
    LocalMux I__856 (
            .O(N__9055),
            .I(\transmit_module.Y_DELTA_PATTERN_48 ));
    InMux I__855 (
            .O(N__9052),
            .I(N__9049));
    LocalMux I__854 (
            .O(N__9049),
            .I(\transmit_module.Y_DELTA_PATTERN_47 ));
    InMux I__853 (
            .O(N__9046),
            .I(N__9043));
    LocalMux I__852 (
            .O(N__9043),
            .I(\transmit_module.Y_DELTA_PATTERN_46 ));
    InMux I__851 (
            .O(N__9040),
            .I(N__9037));
    LocalMux I__850 (
            .O(N__9037),
            .I(\transmit_module.X_DELTA_PATTERN_15 ));
    InMux I__849 (
            .O(N__9034),
            .I(N__9031));
    LocalMux I__848 (
            .O(N__9031),
            .I(\transmit_module.X_DELTA_PATTERN_12 ));
    InMux I__847 (
            .O(N__9028),
            .I(N__9025));
    LocalMux I__846 (
            .O(N__9025),
            .I(\transmit_module.X_DELTA_PATTERN_11 ));
    InMux I__845 (
            .O(N__9022),
            .I(N__9019));
    LocalMux I__844 (
            .O(N__9019),
            .I(\transmit_module.X_DELTA_PATTERN_14 ));
    InMux I__843 (
            .O(N__9016),
            .I(N__9013));
    LocalMux I__842 (
            .O(N__9013),
            .I(\transmit_module.X_DELTA_PATTERN_13 ));
    InMux I__841 (
            .O(N__9010),
            .I(N__9007));
    LocalMux I__840 (
            .O(N__9007),
            .I(\transmit_module.Y_DELTA_PATTERN_64 ));
    InMux I__839 (
            .O(N__9004),
            .I(N__9001));
    LocalMux I__838 (
            .O(N__9001),
            .I(\transmit_module.Y_DELTA_PATTERN_65 ));
    InMux I__837 (
            .O(N__8998),
            .I(N__8995));
    LocalMux I__836 (
            .O(N__8995),
            .I(\transmit_module.Y_DELTA_PATTERN_41 ));
    InMux I__835 (
            .O(N__8992),
            .I(N__8989));
    LocalMux I__834 (
            .O(N__8989),
            .I(\transmit_module.Y_DELTA_PATTERN_92 ));
    InMux I__833 (
            .O(N__8986),
            .I(N__8983));
    LocalMux I__832 (
            .O(N__8983),
            .I(\transmit_module.Y_DELTA_PATTERN_93 ));
    InMux I__831 (
            .O(N__8980),
            .I(N__8977));
    LocalMux I__830 (
            .O(N__8977),
            .I(\transmit_module.Y_DELTA_PATTERN_95 ));
    InMux I__829 (
            .O(N__8974),
            .I(N__8971));
    LocalMux I__828 (
            .O(N__8971),
            .I(\transmit_module.Y_DELTA_PATTERN_94 ));
    InMux I__827 (
            .O(N__8968),
            .I(N__8965));
    LocalMux I__826 (
            .O(N__8965),
            .I(N__8962));
    Odrv4 I__825 (
            .O(N__8962),
            .I(\transmit_module.X_DELTA_PATTERN_8 ));
    InMux I__824 (
            .O(N__8959),
            .I(N__8956));
    LocalMux I__823 (
            .O(N__8956),
            .I(\transmit_module.X_DELTA_PATTERN_7 ));
    InMux I__822 (
            .O(N__8953),
            .I(N__8950));
    LocalMux I__821 (
            .O(N__8950),
            .I(N__8947));
    Odrv4 I__820 (
            .O(N__8947),
            .I(\transmit_module.X_DELTA_PATTERN_10 ));
    InMux I__819 (
            .O(N__8944),
            .I(N__8941));
    LocalMux I__818 (
            .O(N__8941),
            .I(\transmit_module.X_DELTA_PATTERN_6 ));
    InMux I__817 (
            .O(N__8938),
            .I(N__8935));
    LocalMux I__816 (
            .O(N__8935),
            .I(N__8932));
    Odrv12 I__815 (
            .O(N__8932),
            .I(\transmit_module.X_DELTA_PATTERN_5 ));
    InMux I__814 (
            .O(N__8929),
            .I(N__8926));
    LocalMux I__813 (
            .O(N__8926),
            .I(\transmit_module.X_DELTA_PATTERN_4 ));
    InMux I__812 (
            .O(N__8923),
            .I(N__8920));
    LocalMux I__811 (
            .O(N__8920),
            .I(\transmit_module.X_DELTA_PATTERN_9 ));
    InMux I__810 (
            .O(N__8917),
            .I(N__8914));
    LocalMux I__809 (
            .O(N__8914),
            .I(\transmit_module.Y_DELTA_PATTERN_87 ));
    InMux I__808 (
            .O(N__8911),
            .I(N__8908));
    LocalMux I__807 (
            .O(N__8908),
            .I(\transmit_module.Y_DELTA_PATTERN_89 ));
    InMux I__806 (
            .O(N__8905),
            .I(N__8902));
    LocalMux I__805 (
            .O(N__8902),
            .I(\transmit_module.Y_DELTA_PATTERN_88 ));
    InMux I__804 (
            .O(N__8899),
            .I(N__8896));
    LocalMux I__803 (
            .O(N__8896),
            .I(\transmit_module.Y_DELTA_PATTERN_90 ));
    InMux I__802 (
            .O(N__8893),
            .I(N__8890));
    LocalMux I__801 (
            .O(N__8890),
            .I(\transmit_module.Y_DELTA_PATTERN_91 ));
    InMux I__800 (
            .O(N__8887),
            .I(N__8884));
    LocalMux I__799 (
            .O(N__8884),
            .I(\transmit_module.Y_DELTA_PATTERN_77 ));
    InMux I__798 (
            .O(N__8881),
            .I(N__8878));
    LocalMux I__797 (
            .O(N__8878),
            .I(N__8875));
    Span4Mux_s2_v I__796 (
            .O(N__8875),
            .I(N__8871));
    InMux I__795 (
            .O(N__8874),
            .I(N__8868));
    Span4Mux_v I__794 (
            .O(N__8871),
            .I(N__8863));
    LocalMux I__793 (
            .O(N__8868),
            .I(N__8863));
    Span4Mux_v I__792 (
            .O(N__8863),
            .I(N__8859));
    InMux I__791 (
            .O(N__8862),
            .I(N__8856));
    Span4Mux_v I__790 (
            .O(N__8859),
            .I(N__8850));
    LocalMux I__789 (
            .O(N__8856),
            .I(N__8850));
    InMux I__788 (
            .O(N__8855),
            .I(N__8847));
    Span4Mux_v I__787 (
            .O(N__8850),
            .I(N__8842));
    LocalMux I__786 (
            .O(N__8847),
            .I(N__8842));
    Span4Mux_v I__785 (
            .O(N__8842),
            .I(N__8837));
    InMux I__784 (
            .O(N__8841),
            .I(N__8834));
    InMux I__783 (
            .O(N__8840),
            .I(N__8831));
    Span4Mux_v I__782 (
            .O(N__8837),
            .I(N__8826));
    LocalMux I__781 (
            .O(N__8834),
            .I(N__8826));
    LocalMux I__780 (
            .O(N__8831),
            .I(N__8823));
    Span4Mux_h I__779 (
            .O(N__8826),
            .I(N__8819));
    Span4Mux_h I__778 (
            .O(N__8823),
            .I(N__8816));
    InMux I__777 (
            .O(N__8822),
            .I(N__8813));
    Span4Mux_h I__776 (
            .O(N__8819),
            .I(N__8810));
    Span4Mux_v I__775 (
            .O(N__8816),
            .I(N__8806));
    LocalMux I__774 (
            .O(N__8813),
            .I(N__8803));
    Span4Mux_h I__773 (
            .O(N__8810),
            .I(N__8800));
    InMux I__772 (
            .O(N__8809),
            .I(N__8797));
    Span4Mux_v I__771 (
            .O(N__8806),
            .I(N__8792));
    Span4Mux_h I__770 (
            .O(N__8803),
            .I(N__8792));
    Span4Mux_h I__769 (
            .O(N__8800),
            .I(N__8787));
    LocalMux I__768 (
            .O(N__8797),
            .I(N__8787));
    Span4Mux_v I__767 (
            .O(N__8792),
            .I(N__8784));
    Span4Mux_h I__766 (
            .O(N__8787),
            .I(N__8781));
    Span4Mux_v I__765 (
            .O(N__8784),
            .I(N__8778));
    Span4Mux_v I__764 (
            .O(N__8781),
            .I(N__8775));
    Odrv4 I__763 (
            .O(N__8778),
            .I(TVP_VIDEO_c_2));
    Odrv4 I__762 (
            .O(N__8775),
            .I(TVP_VIDEO_c_2));
    InMux I__761 (
            .O(N__8770),
            .I(N__8767));
    LocalMux I__760 (
            .O(N__8767),
            .I(\transmit_module.X_DELTA_PATTERN_3 ));
    InMux I__759 (
            .O(N__8764),
            .I(N__8761));
    LocalMux I__758 (
            .O(N__8761),
            .I(N__8758));
    Odrv4 I__757 (
            .O(N__8758),
            .I(\transmit_module.X_DELTA_PATTERN_2 ));
    InMux I__756 (
            .O(N__8755),
            .I(N__8750));
    InMux I__755 (
            .O(N__8754),
            .I(N__8747));
    InMux I__754 (
            .O(N__8753),
            .I(N__8744));
    LocalMux I__753 (
            .O(N__8750),
            .I(N__8741));
    LocalMux I__752 (
            .O(N__8747),
            .I(N__8734));
    LocalMux I__751 (
            .O(N__8744),
            .I(N__8734));
    Span4Mux_v I__750 (
            .O(N__8741),
            .I(N__8731));
    InMux I__749 (
            .O(N__8740),
            .I(N__8728));
    InMux I__748 (
            .O(N__8739),
            .I(N__8724));
    Span4Mux_v I__747 (
            .O(N__8734),
            .I(N__8721));
    Span4Mux_v I__746 (
            .O(N__8731),
            .I(N__8716));
    LocalMux I__745 (
            .O(N__8728),
            .I(N__8716));
    InMux I__744 (
            .O(N__8727),
            .I(N__8713));
    LocalMux I__743 (
            .O(N__8724),
            .I(N__8708));
    Span4Mux_v I__742 (
            .O(N__8721),
            .I(N__8701));
    Span4Mux_v I__741 (
            .O(N__8716),
            .I(N__8701));
    LocalMux I__740 (
            .O(N__8713),
            .I(N__8701));
    InMux I__739 (
            .O(N__8712),
            .I(N__8698));
    InMux I__738 (
            .O(N__8711),
            .I(N__8695));
    Span4Mux_v I__737 (
            .O(N__8708),
            .I(N__8692));
    Span4Mux_v I__736 (
            .O(N__8701),
            .I(N__8689));
    LocalMux I__735 (
            .O(N__8698),
            .I(N__8686));
    LocalMux I__734 (
            .O(N__8695),
            .I(N__8683));
    Sp12to4 I__733 (
            .O(N__8692),
            .I(N__8680));
    Span4Mux_v I__732 (
            .O(N__8689),
            .I(N__8677));
    Span4Mux_h I__731 (
            .O(N__8686),
            .I(N__8674));
    Span4Mux_h I__730 (
            .O(N__8683),
            .I(N__8671));
    Span12Mux_h I__729 (
            .O(N__8680),
            .I(N__8668));
    Sp12to4 I__728 (
            .O(N__8677),
            .I(N__8665));
    IoSpan4Mux I__727 (
            .O(N__8674),
            .I(N__8662));
    Span4Mux_h I__726 (
            .O(N__8671),
            .I(N__8659));
    Span12Mux_v I__725 (
            .O(N__8668),
            .I(N__8654));
    Span12Mux_h I__724 (
            .O(N__8665),
            .I(N__8654));
    IoSpan4Mux I__723 (
            .O(N__8662),
            .I(N__8649));
    IoSpan4Mux I__722 (
            .O(N__8659),
            .I(N__8649));
    Odrv12 I__721 (
            .O(N__8654),
            .I(TVP_VIDEO_c_8));
    Odrv4 I__720 (
            .O(N__8649),
            .I(TVP_VIDEO_c_8));
    InMux I__719 (
            .O(N__8644),
            .I(N__8641));
    LocalMux I__718 (
            .O(N__8641),
            .I(N__8636));
    InMux I__717 (
            .O(N__8640),
            .I(N__8633));
    InMux I__716 (
            .O(N__8639),
            .I(N__8630));
    Span4Mux_v I__715 (
            .O(N__8636),
            .I(N__8621));
    LocalMux I__714 (
            .O(N__8633),
            .I(N__8621));
    LocalMux I__713 (
            .O(N__8630),
            .I(N__8621));
    InMux I__712 (
            .O(N__8629),
            .I(N__8618));
    InMux I__711 (
            .O(N__8628),
            .I(N__8615));
    Span4Mux_v I__710 (
            .O(N__8621),
            .I(N__8609));
    LocalMux I__709 (
            .O(N__8618),
            .I(N__8609));
    LocalMux I__708 (
            .O(N__8615),
            .I(N__8606));
    InMux I__707 (
            .O(N__8614),
            .I(N__8603));
    Span4Mux_h I__706 (
            .O(N__8609),
            .I(N__8600));
    Span4Mux_h I__705 (
            .O(N__8606),
            .I(N__8597));
    LocalMux I__704 (
            .O(N__8603),
            .I(N__8594));
    Sp12to4 I__703 (
            .O(N__8600),
            .I(N__8588));
    Sp12to4 I__702 (
            .O(N__8597),
            .I(N__8588));
    Span12Mux_s8_h I__701 (
            .O(N__8594),
            .I(N__8585));
    InMux I__700 (
            .O(N__8593),
            .I(N__8582));
    Span12Mux_v I__699 (
            .O(N__8588),
            .I(N__8579));
    Span12Mux_v I__698 (
            .O(N__8585),
            .I(N__8576));
    LocalMux I__697 (
            .O(N__8582),
            .I(N__8573));
    Span12Mux_h I__696 (
            .O(N__8579),
            .I(N__8569));
    Span12Mux_v I__695 (
            .O(N__8576),
            .I(N__8566));
    Span4Mux_h I__694 (
            .O(N__8573),
            .I(N__8563));
    InMux I__693 (
            .O(N__8572),
            .I(N__8560));
    Odrv12 I__692 (
            .O(N__8569),
            .I(TVP_VIDEO_c_9));
    Odrv12 I__691 (
            .O(N__8566),
            .I(TVP_VIDEO_c_9));
    Odrv4 I__690 (
            .O(N__8563),
            .I(TVP_VIDEO_c_9));
    LocalMux I__689 (
            .O(N__8560),
            .I(TVP_VIDEO_c_9));
    InMux I__688 (
            .O(N__8551),
            .I(N__8548));
    LocalMux I__687 (
            .O(N__8548),
            .I(N__8545));
    Span4Mux_v I__686 (
            .O(N__8545),
            .I(N__8541));
    InMux I__685 (
            .O(N__8544),
            .I(N__8538));
    Span4Mux_v I__684 (
            .O(N__8541),
            .I(N__8534));
    LocalMux I__683 (
            .O(N__8538),
            .I(N__8529));
    InMux I__682 (
            .O(N__8537),
            .I(N__8526));
    Span4Mux_v I__681 (
            .O(N__8534),
            .I(N__8523));
    InMux I__680 (
            .O(N__8533),
            .I(N__8520));
    InMux I__679 (
            .O(N__8532),
            .I(N__8517));
    Span12Mux_h I__678 (
            .O(N__8529),
            .I(N__8513));
    LocalMux I__677 (
            .O(N__8526),
            .I(N__8510));
    Span4Mux_v I__676 (
            .O(N__8523),
            .I(N__8505));
    LocalMux I__675 (
            .O(N__8520),
            .I(N__8505));
    LocalMux I__674 (
            .O(N__8517),
            .I(N__8502));
    InMux I__673 (
            .O(N__8516),
            .I(N__8497));
    Span12Mux_v I__672 (
            .O(N__8513),
            .I(N__8494));
    Span4Mux_v I__671 (
            .O(N__8510),
            .I(N__8491));
    Span4Mux_v I__670 (
            .O(N__8505),
            .I(N__8488));
    Span12Mux_h I__669 (
            .O(N__8502),
            .I(N__8485));
    InMux I__668 (
            .O(N__8501),
            .I(N__8482));
    InMux I__667 (
            .O(N__8500),
            .I(N__8479));
    LocalMux I__666 (
            .O(N__8497),
            .I(N__8476));
    Span12Mux_v I__665 (
            .O(N__8494),
            .I(N__8473));
    Sp12to4 I__664 (
            .O(N__8491),
            .I(N__8470));
    Sp12to4 I__663 (
            .O(N__8488),
            .I(N__8467));
    Span12Mux_v I__662 (
            .O(N__8485),
            .I(N__8462));
    LocalMux I__661 (
            .O(N__8482),
            .I(N__8462));
    LocalMux I__660 (
            .O(N__8479),
            .I(N__8459));
    Span4Mux_h I__659 (
            .O(N__8476),
            .I(N__8456));
    Span12Mux_h I__658 (
            .O(N__8473),
            .I(N__8453));
    Span12Mux_h I__657 (
            .O(N__8470),
            .I(N__8448));
    Span12Mux_h I__656 (
            .O(N__8467),
            .I(N__8448));
    Span12Mux_h I__655 (
            .O(N__8462),
            .I(N__8443));
    Span12Mux_h I__654 (
            .O(N__8459),
            .I(N__8443));
    Span4Mux_h I__653 (
            .O(N__8456),
            .I(N__8440));
    Odrv12 I__652 (
            .O(N__8453),
            .I(TVP_VIDEO_c_7));
    Odrv12 I__651 (
            .O(N__8448),
            .I(TVP_VIDEO_c_7));
    Odrv12 I__650 (
            .O(N__8443),
            .I(TVP_VIDEO_c_7));
    Odrv4 I__649 (
            .O(N__8440),
            .I(TVP_VIDEO_c_7));
    InMux I__648 (
            .O(N__8431),
            .I(N__8427));
    InMux I__647 (
            .O(N__8430),
            .I(N__8424));
    LocalMux I__646 (
            .O(N__8427),
            .I(N__8421));
    LocalMux I__645 (
            .O(N__8424),
            .I(N__8417));
    Span4Mux_v I__644 (
            .O(N__8421),
            .I(N__8414));
    InMux I__643 (
            .O(N__8420),
            .I(N__8411));
    Span4Mux_v I__642 (
            .O(N__8417),
            .I(N__8407));
    Span4Mux_v I__641 (
            .O(N__8414),
            .I(N__8402));
    LocalMux I__640 (
            .O(N__8411),
            .I(N__8402));
    InMux I__639 (
            .O(N__8410),
            .I(N__8399));
    Span4Mux_v I__638 (
            .O(N__8407),
            .I(N__8396));
    Span4Mux_v I__637 (
            .O(N__8402),
            .I(N__8390));
    LocalMux I__636 (
            .O(N__8399),
            .I(N__8390));
    Span4Mux_v I__635 (
            .O(N__8396),
            .I(N__8386));
    InMux I__634 (
            .O(N__8395),
            .I(N__8383));
    Span4Mux_v I__633 (
            .O(N__8390),
            .I(N__8379));
    InMux I__632 (
            .O(N__8389),
            .I(N__8376));
    Span4Mux_v I__631 (
            .O(N__8386),
            .I(N__8371));
    LocalMux I__630 (
            .O(N__8383),
            .I(N__8371));
    InMux I__629 (
            .O(N__8382),
            .I(N__8368));
    Span4Mux_v I__628 (
            .O(N__8379),
            .I(N__8363));
    LocalMux I__627 (
            .O(N__8376),
            .I(N__8363));
    Span4Mux_v I__626 (
            .O(N__8371),
            .I(N__8358));
    LocalMux I__625 (
            .O(N__8368),
            .I(N__8358));
    Span4Mux_v I__624 (
            .O(N__8363),
            .I(N__8354));
    Span4Mux_v I__623 (
            .O(N__8358),
            .I(N__8351));
    InMux I__622 (
            .O(N__8357),
            .I(N__8348));
    Sp12to4 I__621 (
            .O(N__8354),
            .I(N__8345));
    Span4Mux_v I__620 (
            .O(N__8351),
            .I(N__8340));
    LocalMux I__619 (
            .O(N__8348),
            .I(N__8340));
    Span12Mux_h I__618 (
            .O(N__8345),
            .I(N__8337));
    Span4Mux_h I__617 (
            .O(N__8340),
            .I(N__8334));
    Odrv12 I__616 (
            .O(N__8337),
            .I(TVP_VIDEO_c_6));
    Odrv4 I__615 (
            .O(N__8334),
            .I(TVP_VIDEO_c_6));
    InMux I__614 (
            .O(N__8329),
            .I(N__8326));
    LocalMux I__613 (
            .O(N__8326),
            .I(N__8322));
    InMux I__612 (
            .O(N__8325),
            .I(N__8318));
    Span4Mux_v I__611 (
            .O(N__8322),
            .I(N__8315));
    InMux I__610 (
            .O(N__8321),
            .I(N__8311));
    LocalMux I__609 (
            .O(N__8318),
            .I(N__8308));
    Span4Mux_v I__608 (
            .O(N__8315),
            .I(N__8304));
    InMux I__607 (
            .O(N__8314),
            .I(N__8301));
    LocalMux I__606 (
            .O(N__8311),
            .I(N__8298));
    Span4Mux_v I__605 (
            .O(N__8308),
            .I(N__8295));
    InMux I__604 (
            .O(N__8307),
            .I(N__8292));
    Span4Mux_v I__603 (
            .O(N__8304),
            .I(N__8286));
    LocalMux I__602 (
            .O(N__8301),
            .I(N__8286));
    Span4Mux_h I__601 (
            .O(N__8298),
            .I(N__8282));
    Span4Mux_v I__600 (
            .O(N__8295),
            .I(N__8277));
    LocalMux I__599 (
            .O(N__8292),
            .I(N__8277));
    InMux I__598 (
            .O(N__8291),
            .I(N__8274));
    Span4Mux_v I__597 (
            .O(N__8286),
            .I(N__8271));
    InMux I__596 (
            .O(N__8285),
            .I(N__8268));
    Sp12to4 I__595 (
            .O(N__8282),
            .I(N__8265));
    Span4Mux_v I__594 (
            .O(N__8277),
            .I(N__8260));
    LocalMux I__593 (
            .O(N__8274),
            .I(N__8260));
    Span4Mux_v I__592 (
            .O(N__8271),
            .I(N__8255));
    LocalMux I__591 (
            .O(N__8268),
            .I(N__8255));
    Span12Mux_v I__590 (
            .O(N__8265),
            .I(N__8251));
    Span4Mux_v I__589 (
            .O(N__8260),
            .I(N__8248));
    Span4Mux_v I__588 (
            .O(N__8255),
            .I(N__8245));
    InMux I__587 (
            .O(N__8254),
            .I(N__8242));
    Span12Mux_v I__586 (
            .O(N__8251),
            .I(N__8237));
    Sp12to4 I__585 (
            .O(N__8248),
            .I(N__8237));
    Span4Mux_v I__584 (
            .O(N__8245),
            .I(N__8232));
    LocalMux I__583 (
            .O(N__8242),
            .I(N__8232));
    Span12Mux_h I__582 (
            .O(N__8237),
            .I(N__8229));
    Span4Mux_h I__581 (
            .O(N__8232),
            .I(N__8226));
    Odrv12 I__580 (
            .O(N__8229),
            .I(TVP_VIDEO_c_5));
    Odrv4 I__579 (
            .O(N__8226),
            .I(TVP_VIDEO_c_5));
    InMux I__578 (
            .O(N__8221),
            .I(N__8218));
    LocalMux I__577 (
            .O(N__8218),
            .I(N__8215));
    Span4Mux_v I__576 (
            .O(N__8215),
            .I(N__8209));
    InMux I__575 (
            .O(N__8214),
            .I(N__8206));
    InMux I__574 (
            .O(N__8213),
            .I(N__8202));
    InMux I__573 (
            .O(N__8212),
            .I(N__8198));
    Span4Mux_v I__572 (
            .O(N__8209),
            .I(N__8193));
    LocalMux I__571 (
            .O(N__8206),
            .I(N__8193));
    InMux I__570 (
            .O(N__8205),
            .I(N__8190));
    LocalMux I__569 (
            .O(N__8202),
            .I(N__8187));
    InMux I__568 (
            .O(N__8201),
            .I(N__8184));
    LocalMux I__567 (
            .O(N__8198),
            .I(N__8181));
    Span4Mux_v I__566 (
            .O(N__8193),
            .I(N__8176));
    LocalMux I__565 (
            .O(N__8190),
            .I(N__8176));
    Span4Mux_h I__564 (
            .O(N__8187),
            .I(N__8173));
    LocalMux I__563 (
            .O(N__8184),
            .I(N__8170));
    Span4Mux_s1_v I__562 (
            .O(N__8181),
            .I(N__8166));
    Span4Mux_v I__561 (
            .O(N__8176),
            .I(N__8163));
    Span4Mux_h I__560 (
            .O(N__8173),
            .I(N__8160));
    Span4Mux_h I__559 (
            .O(N__8170),
            .I(N__8157));
    InMux I__558 (
            .O(N__8169),
            .I(N__8154));
    Sp12to4 I__557 (
            .O(N__8166),
            .I(N__8151));
    Span4Mux_h I__556 (
            .O(N__8163),
            .I(N__8148));
    Span4Mux_h I__555 (
            .O(N__8160),
            .I(N__8145));
    Span4Mux_v I__554 (
            .O(N__8157),
            .I(N__8142));
    LocalMux I__553 (
            .O(N__8154),
            .I(N__8139));
    Span12Mux_s10_h I__552 (
            .O(N__8151),
            .I(N__8135));
    Sp12to4 I__551 (
            .O(N__8148),
            .I(N__8132));
    Span4Mux_h I__550 (
            .O(N__8145),
            .I(N__8125));
    Span4Mux_v I__549 (
            .O(N__8142),
            .I(N__8125));
    Span4Mux_h I__548 (
            .O(N__8139),
            .I(N__8125));
    InMux I__547 (
            .O(N__8138),
            .I(N__8122));
    Span12Mux_v I__546 (
            .O(N__8135),
            .I(N__8119));
    Span12Mux_h I__545 (
            .O(N__8132),
            .I(N__8116));
    Span4Mux_v I__544 (
            .O(N__8125),
            .I(N__8113));
    LocalMux I__543 (
            .O(N__8122),
            .I(N__8110));
    Span12Mux_v I__542 (
            .O(N__8119),
            .I(N__8107));
    Span12Mux_v I__541 (
            .O(N__8116),
            .I(N__8104));
    Span4Mux_v I__540 (
            .O(N__8113),
            .I(N__8101));
    Span4Mux_h I__539 (
            .O(N__8110),
            .I(N__8098));
    Odrv12 I__538 (
            .O(N__8107),
            .I(TVP_VIDEO_c_4));
    Odrv12 I__537 (
            .O(N__8104),
            .I(TVP_VIDEO_c_4));
    Odrv4 I__536 (
            .O(N__8101),
            .I(TVP_VIDEO_c_4));
    Odrv4 I__535 (
            .O(N__8098),
            .I(TVP_VIDEO_c_4));
    InMux I__534 (
            .O(N__8089),
            .I(N__8085));
    InMux I__533 (
            .O(N__8088),
            .I(N__8082));
    LocalMux I__532 (
            .O(N__8085),
            .I(N__8078));
    LocalMux I__531 (
            .O(N__8082),
            .I(N__8075));
    InMux I__530 (
            .O(N__8081),
            .I(N__8072));
    Sp12to4 I__529 (
            .O(N__8078),
            .I(N__8068));
    Span4Mux_h I__528 (
            .O(N__8075),
            .I(N__8065));
    LocalMux I__527 (
            .O(N__8072),
            .I(N__8062));
    InMux I__526 (
            .O(N__8071),
            .I(N__8058));
    Span12Mux_h I__525 (
            .O(N__8068),
            .I(N__8053));
    Span4Mux_h I__524 (
            .O(N__8065),
            .I(N__8050));
    Span4Mux_v I__523 (
            .O(N__8062),
            .I(N__8047));
    InMux I__522 (
            .O(N__8061),
            .I(N__8044));
    LocalMux I__521 (
            .O(N__8058),
            .I(N__8041));
    InMux I__520 (
            .O(N__8057),
            .I(N__8038));
    InMux I__519 (
            .O(N__8056),
            .I(N__8034));
    Span12Mux_v I__518 (
            .O(N__8053),
            .I(N__8029));
    Sp12to4 I__517 (
            .O(N__8050),
            .I(N__8029));
    Sp12to4 I__516 (
            .O(N__8047),
            .I(N__8026));
    LocalMux I__515 (
            .O(N__8044),
            .I(N__8023));
    Span12Mux_h I__514 (
            .O(N__8041),
            .I(N__8020));
    LocalMux I__513 (
            .O(N__8038),
            .I(N__8017));
    InMux I__512 (
            .O(N__8037),
            .I(N__8014));
    LocalMux I__511 (
            .O(N__8034),
            .I(N__8011));
    Span12Mux_v I__510 (
            .O(N__8029),
            .I(N__8006));
    Span12Mux_h I__509 (
            .O(N__8026),
            .I(N__8006));
    Span12Mux_h I__508 (
            .O(N__8023),
            .I(N__8003));
    Span12Mux_v I__507 (
            .O(N__8020),
            .I(N__7996));
    Span12Mux_h I__506 (
            .O(N__8017),
            .I(N__7996));
    LocalMux I__505 (
            .O(N__8014),
            .I(N__7996));
    Span4Mux_h I__504 (
            .O(N__8011),
            .I(N__7993));
    Span12Mux_h I__503 (
            .O(N__8006),
            .I(N__7988));
    Span12Mux_v I__502 (
            .O(N__8003),
            .I(N__7988));
    Span12Mux_h I__501 (
            .O(N__7996),
            .I(N__7985));
    Span4Mux_v I__500 (
            .O(N__7993),
            .I(N__7982));
    Odrv12 I__499 (
            .O(N__7988),
            .I(TVP_VIDEO_c_3));
    Odrv12 I__498 (
            .O(N__7985),
            .I(TVP_VIDEO_c_3));
    Odrv4 I__497 (
            .O(N__7982),
            .I(TVP_VIDEO_c_3));
    INV \INVsync_buffer.WIRE_OUT_8C  (
            .O(\INVsync_buffer.WIRE_OUT_8C_net ),
            .I(N__22997));
    defparam IN_MUX_bfv_12_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_13_0_));
    defparam IN_MUX_bfv_12_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_14_0_ (
            .carryinitin(\transmit_module.video_signal_controller.n3297 ),
            .carryinitout(bfn_12_14_0_));
    defparam IN_MUX_bfv_10_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_15_0_));
    defparam IN_MUX_bfv_10_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_16_0_ (
            .carryinitin(\transmit_module.video_signal_controller.n3286 ),
            .carryinitout(bfn_10_16_0_));
    defparam IN_MUX_bfv_15_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_13_0_));
    defparam IN_MUX_bfv_15_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_14_0_ (
            .carryinitin(\transmit_module.n3265 ),
            .carryinitout(bfn_15_14_0_));
    defparam IN_MUX_bfv_13_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_10_0_));
    defparam IN_MUX_bfv_13_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_11_0_ (
            .carryinitin(\receive_module.rx_counter.n3278 ),
            .carryinitout(bfn_13_11_0_));
    defparam IN_MUX_bfv_17_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_10_0_));
    defparam IN_MUX_bfv_17_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_11_0_ (
            .carryinitin(\receive_module.rx_counter.n3308 ),
            .carryinitout(bfn_17_11_0_));
    defparam IN_MUX_bfv_16_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_5_0_));
    defparam IN_MUX_bfv_15_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_11_0_));
    defparam IN_MUX_bfv_15_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_12_0_ (
            .carryinitin(\receive_module.n3252 ),
            .carryinitout(bfn_15_12_0_));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \transmit_module.X_DELTA_PATTERN_i1_LC_7_12_5 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i1_LC_7_12_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.X_DELTA_PATTERN_i1_LC_7_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i1_LC_7_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8764),
            .lcout(\transmit_module.X_DELTA_PATTERN_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23190),
            .ce(N__11128),
            .sr(N__21488));
    defparam \transmit_module.X_DELTA_PATTERN_i3_LC_7_15_0 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i3_LC_7_15_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.X_DELTA_PATTERN_i3_LC_7_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i3_LC_7_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8929),
            .lcout(\transmit_module.X_DELTA_PATTERN_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23224),
            .ce(N__11122),
            .sr(N__21458));
    defparam \transmit_module.X_DELTA_PATTERN_i2_LC_7_15_2 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i2_LC_7_15_2 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i2_LC_7_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i2_LC_7_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8770),
            .lcout(\transmit_module.X_DELTA_PATTERN_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23224),
            .ce(N__11122),
            .sr(N__21458));
    defparam \transmit_module.X_DELTA_PATTERN_i8_LC_7_15_3 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i8_LC_7_15_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.X_DELTA_PATTERN_i8_LC_7_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i8_LC_7_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8923),
            .lcout(\transmit_module.X_DELTA_PATTERN_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23224),
            .ce(N__11122),
            .sr(N__21458));
    defparam \transmit_module.X_DELTA_PATTERN_i4_LC_7_15_4 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i4_LC_7_15_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i4_LC_7_15_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i4_LC_7_15_4  (
            .in0(N__8938),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.X_DELTA_PATTERN_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23224),
            .ce(N__11122),
            .sr(N__21458));
    defparam \transmit_module.X_DELTA_PATTERN_i9_LC_7_15_6 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i9_LC_7_15_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i9_LC_7_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i9_LC_7_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8953),
            .lcout(\transmit_module.X_DELTA_PATTERN_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23224),
            .ce(N__11122),
            .sr(N__21458));
    defparam \transmit_module.Y_DELTA_PATTERN_i89_LC_9_11_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i89_LC_9_11_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i89_LC_9_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i89_LC_9_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8899),
            .lcout(\transmit_module.Y_DELTA_PATTERN_89 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23268),
            .ce(N__11074),
            .sr(N__21320));
    defparam \transmit_module.Y_DELTA_PATTERN_i86_LC_9_11_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i86_LC_9_11_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i86_LC_9_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i86_LC_9_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8917),
            .lcout(\transmit_module.Y_DELTA_PATTERN_86 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23268),
            .ce(N__11074),
            .sr(N__21320));
    defparam \transmit_module.Y_DELTA_PATTERN_i87_LC_9_11_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i87_LC_9_11_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i87_LC_9_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i87_LC_9_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8905),
            .lcout(\transmit_module.Y_DELTA_PATTERN_87 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23268),
            .ce(N__11074),
            .sr(N__21320));
    defparam \transmit_module.Y_DELTA_PATTERN_i88_LC_9_11_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i88_LC_9_11_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i88_LC_9_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i88_LC_9_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8911),
            .lcout(\transmit_module.Y_DELTA_PATTERN_88 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23268),
            .ce(N__11074),
            .sr(N__21320));
    defparam \transmit_module.Y_DELTA_PATTERN_i76_LC_9_12_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i76_LC_9_12_2 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i76_LC_9_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i76_LC_9_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8887),
            .lcout(\transmit_module.Y_DELTA_PATTERN_76 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23225),
            .ce(N__11073),
            .sr(N__21348));
    defparam \transmit_module.Y_DELTA_PATTERN_i90_LC_9_12_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i90_LC_9_12_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i90_LC_9_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i90_LC_9_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8893),
            .lcout(\transmit_module.Y_DELTA_PATTERN_90 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23225),
            .ce(N__11073),
            .sr(N__21348));
    defparam \transmit_module.Y_DELTA_PATTERN_i91_LC_9_12_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i91_LC_9_12_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i91_LC_9_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i91_LC_9_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8992),
            .lcout(\transmit_module.Y_DELTA_PATTERN_91 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23225),
            .ce(N__11073),
            .sr(N__21348));
    defparam \transmit_module.Y_DELTA_PATTERN_i77_LC_9_12_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i77_LC_9_12_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i77_LC_9_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i77_LC_9_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9319),
            .lcout(\transmit_module.Y_DELTA_PATTERN_77 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23225),
            .ce(N__11073),
            .sr(N__21348));
    defparam \transmit_module.Y_DELTA_PATTERN_i92_LC_9_12_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i92_LC_9_12_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i92_LC_9_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i92_LC_9_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8986),
            .lcout(\transmit_module.Y_DELTA_PATTERN_92 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23225),
            .ce(N__11073),
            .sr(N__21348));
    defparam \transmit_module.Y_DELTA_PATTERN_i93_LC_9_13_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i93_LC_9_13_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i93_LC_9_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i93_LC_9_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8974),
            .lcout(\transmit_module.Y_DELTA_PATTERN_93 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23160),
            .ce(N__11069),
            .sr(N__21351));
    defparam \transmit_module.Y_DELTA_PATTERN_i95_LC_9_13_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i95_LC_9_13_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i95_LC_9_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i95_LC_9_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9121),
            .lcout(\transmit_module.Y_DELTA_PATTERN_95 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23160),
            .ce(N__11069),
            .sr(N__21351));
    defparam \transmit_module.Y_DELTA_PATTERN_i94_LC_9_14_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i94_LC_9_14_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i94_LC_9_14_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i94_LC_9_14_5  (
            .in0(N__8980),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.Y_DELTA_PATTERN_94 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23080),
            .ce(N__21460),
            .sr(N__21304));
    defparam \transmit_module.X_DELTA_PATTERN_i7_LC_9_15_0 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i7_LC_9_15_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i7_LC_9_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i7_LC_9_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8968),
            .lcout(\transmit_module.X_DELTA_PATTERN_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23175),
            .ce(N__11106),
            .sr(N__21457));
    defparam \transmit_module.X_DELTA_PATTERN_i6_LC_9_15_1 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i6_LC_9_15_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i6_LC_9_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i6_LC_9_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8959),
            .lcout(\transmit_module.X_DELTA_PATTERN_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23175),
            .ce(N__11106),
            .sr(N__21457));
    defparam \transmit_module.X_DELTA_PATTERN_i15_LC_9_15_2 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i15_LC_9_15_2 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i15_LC_9_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i15_LC_9_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13426),
            .lcout(\transmit_module.X_DELTA_PATTERN_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23175),
            .ce(N__11106),
            .sr(N__21457));
    defparam \transmit_module.X_DELTA_PATTERN_i10_LC_9_15_4 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i10_LC_9_15_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.X_DELTA_PATTERN_i10_LC_9_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i10_LC_9_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9028),
            .lcout(\transmit_module.X_DELTA_PATTERN_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23175),
            .ce(N__11106),
            .sr(N__21457));
    defparam \transmit_module.X_DELTA_PATTERN_i5_LC_9_15_6 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i5_LC_9_15_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.X_DELTA_PATTERN_i5_LC_9_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i5_LC_9_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8944),
            .lcout(\transmit_module.X_DELTA_PATTERN_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23175),
            .ce(N__11106),
            .sr(N__21457));
    defparam \transmit_module.X_DELTA_PATTERN_i14_LC_9_15_7 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i14_LC_9_15_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.X_DELTA_PATTERN_i14_LC_9_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i14_LC_9_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9040),
            .lcout(\transmit_module.X_DELTA_PATTERN_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23175),
            .ce(N__11106),
            .sr(N__21457));
    defparam \transmit_module.X_DELTA_PATTERN_i12_LC_9_16_0 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i12_LC_9_16_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.X_DELTA_PATTERN_i12_LC_9_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i12_LC_9_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9016),
            .lcout(\transmit_module.X_DELTA_PATTERN_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23055),
            .ce(N__11127),
            .sr(N__21474));
    defparam \transmit_module.X_DELTA_PATTERN_i11_LC_9_16_3 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i11_LC_9_16_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i11_LC_9_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i11_LC_9_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9034),
            .lcout(\transmit_module.X_DELTA_PATTERN_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23055),
            .ce(N__11127),
            .sr(N__21474));
    defparam \transmit_module.X_DELTA_PATTERN_i13_LC_9_16_6 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i13_LC_9_16_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i13_LC_9_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i13_LC_9_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9022),
            .lcout(\transmit_module.X_DELTA_PATTERN_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23055),
            .ce(N__11127),
            .sr(N__21474));
    defparam \transmit_module.Y_DELTA_PATTERN_i40_LC_10_10_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i40_LC_10_10_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i40_LC_10_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i40_LC_10_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8998),
            .lcout(\transmit_module.Y_DELTA_PATTERN_40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23151),
            .ce(N__10051),
            .sr(N__21350));
    defparam \transmit_module.Y_DELTA_PATTERN_i64_LC_10_11_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i64_LC_10_11_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i64_LC_10_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i64_LC_10_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9004),
            .lcout(\transmit_module.Y_DELTA_PATTERN_64 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23292),
            .ce(N__10039),
            .sr(N__21325));
    defparam \transmit_module.Y_DELTA_PATTERN_i63_LC_10_11_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i63_LC_10_11_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i63_LC_10_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i63_LC_10_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9010),
            .lcout(\transmit_module.Y_DELTA_PATTERN_63 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23292),
            .ce(N__10039),
            .sr(N__21325));
    defparam \transmit_module.Y_DELTA_PATTERN_i65_LC_10_11_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i65_LC_10_11_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i65_LC_10_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i65_LC_10_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9283),
            .lcout(\transmit_module.Y_DELTA_PATTERN_65 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23292),
            .ce(N__10039),
            .sr(N__21325));
    defparam \transmit_module.Y_DELTA_PATTERN_i41_LC_10_11_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i41_LC_10_11_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i41_LC_10_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i41_LC_10_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9130),
            .lcout(\transmit_module.Y_DELTA_PATTERN_41 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23292),
            .ce(N__10039),
            .sr(N__21325));
    defparam \transmit_module.Y_DELTA_PATTERN_i62_LC_10_11_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i62_LC_10_11_7 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i62_LC_10_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i62_LC_10_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9088),
            .lcout(\transmit_module.Y_DELTA_PATTERN_62 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23292),
            .ce(N__10039),
            .sr(N__21325));
    defparam \transmit_module.Y_DELTA_PATTERN_i73_LC_10_12_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i73_LC_10_12_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i73_LC_10_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i73_LC_10_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9082),
            .lcout(\transmit_module.Y_DELTA_PATTERN_73 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23134),
            .ce(N__10049),
            .sr(N__21349));
    defparam \transmit_module.Y_DELTA_PATTERN_i74_LC_10_12_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i74_LC_10_12_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i74_LC_10_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i74_LC_10_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9070),
            .lcout(\transmit_module.Y_DELTA_PATTERN_74 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23134),
            .ce(N__10049),
            .sr(N__21349));
    defparam \transmit_module.Y_DELTA_PATTERN_i75_LC_10_12_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i75_LC_10_12_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i75_LC_10_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i75_LC_10_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9076),
            .lcout(\transmit_module.Y_DELTA_PATTERN_75 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23134),
            .ce(N__10049),
            .sr(N__21349));
    defparam \transmit_module.Y_DELTA_PATTERN_i72_LC_10_12_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i72_LC_10_12_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i72_LC_10_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i72_LC_10_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9064),
            .lcout(\transmit_module.Y_DELTA_PATTERN_72 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23134),
            .ce(N__10049),
            .sr(N__21349));
    defparam \transmit_module.Y_DELTA_PATTERN_i48_LC_10_12_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i48_LC_10_12_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i48_LC_10_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i48_LC_10_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9358),
            .lcout(\transmit_module.Y_DELTA_PATTERN_48 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23134),
            .ce(N__10049),
            .sr(N__21349));
    defparam \transmit_module.Y_DELTA_PATTERN_i46_LC_10_12_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i46_LC_10_12_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i46_LC_10_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i46_LC_10_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9052),
            .lcout(\transmit_module.Y_DELTA_PATTERN_46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23134),
            .ce(N__10049),
            .sr(N__21349));
    defparam \transmit_module.Y_DELTA_PATTERN_i47_LC_10_12_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i47_LC_10_12_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i47_LC_10_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i47_LC_10_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9058),
            .lcout(\transmit_module.Y_DELTA_PATTERN_47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23134),
            .ce(N__10049),
            .sr(N__21349));
    defparam \transmit_module.Y_DELTA_PATTERN_i45_LC_10_12_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i45_LC_10_12_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i45_LC_10_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i45_LC_10_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9046),
            .lcout(\transmit_module.Y_DELTA_PATTERN_45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23134),
            .ce(N__10049),
            .sr(N__21349));
    defparam \transmit_module.Y_DELTA_PATTERN_i42_LC_10_13_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i42_LC_10_13_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i42_LC_10_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i42_LC_10_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9103),
            .lcout(\transmit_module.Y_DELTA_PATTERN_42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23201),
            .ce(N__10054),
            .sr(N__21347));
    defparam \transmit_module.Y_DELTA_PATTERN_i96_LC_10_13_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i96_LC_10_13_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i96_LC_10_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i96_LC_10_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9220),
            .lcout(\transmit_module.Y_DELTA_PATTERN_96 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23201),
            .ce(N__10054),
            .sr(N__21347));
    defparam \transmit_module.Y_DELTA_PATTERN_i44_LC_10_13_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i44_LC_10_13_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i44_LC_10_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i44_LC_10_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9115),
            .lcout(\transmit_module.Y_DELTA_PATTERN_44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23201),
            .ce(N__10054),
            .sr(N__21347));
    defparam \transmit_module.Y_DELTA_PATTERN_i43_LC_10_13_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i43_LC_10_13_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i43_LC_10_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i43_LC_10_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9109),
            .lcout(\transmit_module.Y_DELTA_PATTERN_43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23201),
            .ce(N__10054),
            .sr(N__21347));
    defparam \transmit_module.video_signal_controller.i1653_2_lut_3_lut_LC_10_14_0 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1653_2_lut_3_lut_LC_10_14_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1653_2_lut_3_lut_LC_10_14_0 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \transmit_module.video_signal_controller.i1653_2_lut_3_lut_LC_10_14_0  (
            .in0(_gnd_net_),
            .in1(N__9163),
            .in2(N__9190),
            .in3(N__9206),
            .lcout(\transmit_module.video_signal_controller.n2886 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_2_lut_adj_23_LC_10_14_2 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_2_lut_adj_23_LC_10_14_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_2_lut_adj_23_LC_10_14_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \transmit_module.video_signal_controller.i1_2_lut_adj_23_LC_10_14_2  (
            .in0(_gnd_net_),
            .in1(N__9550),
            .in2(_gnd_net_),
            .in3(N__9415),
            .lcout(\transmit_module.video_signal_controller.n3467 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1643_2_lut_LC_10_14_3 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1643_2_lut_LC_10_14_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1643_2_lut_LC_10_14_3 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \transmit_module.video_signal_controller.i1643_2_lut_LC_10_14_3  (
            .in0(N__9207),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9188),
            .lcout(\transmit_module.video_signal_controller.n2876 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_21_LC_10_14_4 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_21_LC_10_14_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_21_LC_10_14_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \transmit_module.video_signal_controller.i1_2_lut_rep_21_LC_10_14_4  (
            .in0(_gnd_net_),
            .in1(N__9662),
            .in2(_gnd_net_),
            .in3(N__9392),
            .lcout(),
            .ltout(\transmit_module.video_signal_controller.n3788_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_4_lut_adj_25_LC_10_14_5 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_4_lut_adj_25_LC_10_14_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_4_lut_adj_25_LC_10_14_5 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \transmit_module.video_signal_controller.i1_4_lut_adj_25_LC_10_14_5  (
            .in0(N__9165),
            .in1(N__9421),
            .in2(N__9097),
            .in3(N__9094),
            .lcout(\transmit_module.video_signal_controller.n4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i495_2_lut_rep_22_LC_10_14_6 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i495_2_lut_rep_22_LC_10_14_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i495_2_lut_rep_22_LC_10_14_6 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \transmit_module.video_signal_controller.i495_2_lut_rep_22_LC_10_14_6  (
            .in0(N__9187),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9164),
            .lcout(\transmit_module.video_signal_controller.n3789 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.VGA_X_i0_LC_10_15_0 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i0_LC_10_15_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i0_LC_10_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i0_LC_10_15_0  (
            .in0(_gnd_net_),
            .in1(N__9208),
            .in2(_gnd_net_),
            .in3(N__9193),
            .lcout(\transmit_module.video_signal_controller.VGA_X_0 ),
            .ltout(),
            .carryin(bfn_10_15_0_),
            .carryout(\transmit_module.video_signal_controller.n3279 ),
            .clk(N__23174),
            .ce(),
            .sr(N__9790));
    defparam \transmit_module.video_signal_controller.VGA_X_i1_LC_10_15_1 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i1_LC_10_15_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i1_LC_10_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i1_LC_10_15_1  (
            .in0(_gnd_net_),
            .in1(N__9189),
            .in2(_gnd_net_),
            .in3(N__9169),
            .lcout(\transmit_module.video_signal_controller.VGA_X_1 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3279 ),
            .carryout(\transmit_module.video_signal_controller.n3280 ),
            .clk(N__23174),
            .ce(),
            .sr(N__9790));
    defparam \transmit_module.video_signal_controller.VGA_X_i2_LC_10_15_2 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i2_LC_10_15_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i2_LC_10_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i2_LC_10_15_2  (
            .in0(_gnd_net_),
            .in1(N__9166),
            .in2(_gnd_net_),
            .in3(N__9148),
            .lcout(\transmit_module.video_signal_controller.VGA_X_2 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3280 ),
            .carryout(\transmit_module.video_signal_controller.n3281 ),
            .clk(N__23174),
            .ce(),
            .sr(N__9790));
    defparam \transmit_module.video_signal_controller.VGA_X_i3_LC_10_15_3 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i3_LC_10_15_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i3_LC_10_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i3_LC_10_15_3  (
            .in0(_gnd_net_),
            .in1(N__9419),
            .in2(_gnd_net_),
            .in3(N__9145),
            .lcout(\transmit_module.video_signal_controller.VGA_X_3 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3281 ),
            .carryout(\transmit_module.video_signal_controller.n3282 ),
            .clk(N__23174),
            .ce(),
            .sr(N__9790));
    defparam \transmit_module.video_signal_controller.VGA_X_i4_LC_10_15_4 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i4_LC_10_15_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i4_LC_10_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i4_LC_10_15_4  (
            .in0(_gnd_net_),
            .in1(N__9551),
            .in2(_gnd_net_),
            .in3(N__9142),
            .lcout(\transmit_module.video_signal_controller.VGA_X_4 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3282 ),
            .carryout(\transmit_module.video_signal_controller.n3283 ),
            .clk(N__23174),
            .ce(),
            .sr(N__9790));
    defparam \transmit_module.video_signal_controller.VGA_X_i5_LC_10_15_5 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i5_LC_10_15_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i5_LC_10_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i5_LC_10_15_5  (
            .in0(_gnd_net_),
            .in1(N__9393),
            .in2(_gnd_net_),
            .in3(N__9139),
            .lcout(\transmit_module.video_signal_controller.VGA_X_5 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3283 ),
            .carryout(\transmit_module.video_signal_controller.n3284 ),
            .clk(N__23174),
            .ce(),
            .sr(N__9790));
    defparam \transmit_module.video_signal_controller.VGA_X_i6_LC_10_15_6 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i6_LC_10_15_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i6_LC_10_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i6_LC_10_15_6  (
            .in0(_gnd_net_),
            .in1(N__9663),
            .in2(_gnd_net_),
            .in3(N__9136),
            .lcout(\transmit_module.video_signal_controller.VGA_X_6 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3284 ),
            .carryout(\transmit_module.video_signal_controller.n3285 ),
            .clk(N__23174),
            .ce(),
            .sr(N__9790));
    defparam \transmit_module.video_signal_controller.VGA_X_i7_LC_10_15_7 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i7_LC_10_15_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i7_LC_10_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i7_LC_10_15_7  (
            .in0(_gnd_net_),
            .in1(N__9575),
            .in2(_gnd_net_),
            .in3(N__9133),
            .lcout(\transmit_module.video_signal_controller.VGA_X_7 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3285 ),
            .carryout(\transmit_module.video_signal_controller.n3286 ),
            .clk(N__23174),
            .ce(),
            .sr(N__9790));
    defparam \transmit_module.video_signal_controller.VGA_X_i8_LC_10_16_0 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i8_LC_10_16_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i8_LC_10_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i8_LC_10_16_0  (
            .in0(_gnd_net_),
            .in1(N__9688),
            .in2(_gnd_net_),
            .in3(N__9256),
            .lcout(\transmit_module.video_signal_controller.VGA_X_8 ),
            .ltout(),
            .carryin(bfn_10_16_0_),
            .carryout(\transmit_module.video_signal_controller.n3287 ),
            .clk(N__23189),
            .ce(),
            .sr(N__9786));
    defparam \transmit_module.video_signal_controller.VGA_X_i9_LC_10_16_1 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i9_LC_10_16_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i9_LC_10_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i9_LC_10_16_1  (
            .in0(_gnd_net_),
            .in1(N__9635),
            .in2(_gnd_net_),
            .in3(N__9253),
            .lcout(\transmit_module.video_signal_controller.VGA_X_9 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3287 ),
            .carryout(\transmit_module.video_signal_controller.n3288 ),
            .clk(N__23189),
            .ce(),
            .sr(N__9786));
    defparam \transmit_module.video_signal_controller.VGA_X_i10_LC_10_16_2 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i10_LC_10_16_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i10_LC_10_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i10_LC_10_16_2  (
            .in0(_gnd_net_),
            .in1(N__9606),
            .in2(_gnd_net_),
            .in3(N__9250),
            .lcout(\transmit_module.video_signal_controller.VGA_X_10 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3288 ),
            .carryout(\transmit_module.video_signal_controller.n3289 ),
            .clk(N__23189),
            .ce(),
            .sr(N__9786));
    defparam \transmit_module.video_signal_controller.VGA_X_i11_LC_10_16_3 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.VGA_X_i11_LC_10_16_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i11_LC_10_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i11_LC_10_16_3  (
            .in0(_gnd_net_),
            .in1(N__10489),
            .in2(_gnd_net_),
            .in3(N__9247),
            .lcout(\transmit_module.video_signal_controller.VGA_X_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23189),
            .ce(),
            .sr(N__9786));
    defparam \transmit_module.Y_DELTA_PATTERN_i53_LC_11_9_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i53_LC_11_9_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i53_LC_11_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i53_LC_11_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9238),
            .lcout(\transmit_module.Y_DELTA_PATTERN_53 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23079),
            .ce(N__10053),
            .sr(N__21324));
    defparam \transmit_module.Y_DELTA_PATTERN_i55_LC_11_9_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i55_LC_11_9_2 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i55_LC_11_9_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i55_LC_11_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9226),
            .lcout(\transmit_module.Y_DELTA_PATTERN_55 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23079),
            .ce(N__10053),
            .sr(N__21324));
    defparam \transmit_module.Y_DELTA_PATTERN_i54_LC_11_9_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i54_LC_11_9_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i54_LC_11_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i54_LC_11_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9244),
            .lcout(\transmit_module.Y_DELTA_PATTERN_54 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23079),
            .ce(N__10053),
            .sr(N__21324));
    defparam \transmit_module.Y_DELTA_PATTERN_i39_LC_11_10_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i39_LC_11_10_2 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i39_LC_11_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i39_LC_11_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9232),
            .lcout(\transmit_module.Y_DELTA_PATTERN_39 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23199),
            .ce(N__10052),
            .sr(N__21330));
    defparam \transmit_module.Y_DELTA_PATTERN_i56_LC_11_10_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i56_LC_11_10_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i56_LC_11_10_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i56_LC_11_10_3  (
            .in0(N__9496),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.Y_DELTA_PATTERN_56 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23199),
            .ce(N__10052),
            .sr(N__21330));
    defparam \transmit_module.Y_DELTA_PATTERN_i97_LC_11_10_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i97_LC_11_10_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i97_LC_11_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i97_LC_11_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9742),
            .lcout(\transmit_module.Y_DELTA_PATTERN_97 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23199),
            .ce(N__10052),
            .sr(N__21330));
    defparam \transmit_module.Y_DELTA_PATTERN_i35_LC_11_10_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i35_LC_11_10_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i35_LC_11_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i35_LC_11_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9295),
            .lcout(\transmit_module.Y_DELTA_PATTERN_35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23199),
            .ce(N__10052),
            .sr(N__21330));
    defparam \transmit_module.Y_DELTA_PATTERN_i36_LC_11_10_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i36_LC_11_10_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i36_LC_11_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i36_LC_11_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9520),
            .lcout(\transmit_module.Y_DELTA_PATTERN_36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23199),
            .ce(N__10052),
            .sr(N__21330));
    defparam \transmit_module.Y_DELTA_PATTERN_i61_LC_11_11_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i61_LC_11_11_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i61_LC_11_11_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i61_LC_11_11_1  (
            .in0(N__9289),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.Y_DELTA_PATTERN_61 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23081),
            .ce(N__10035),
            .sr(N__21329));
    defparam \transmit_module.Y_DELTA_PATTERN_i66_LC_11_11_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i66_LC_11_11_2 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i66_LC_11_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i66_LC_11_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9472),
            .lcout(\transmit_module.Y_DELTA_PATTERN_66 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23081),
            .ce(N__10035),
            .sr(N__21329));
    defparam \transmit_module.Y_DELTA_PATTERN_i52_LC_11_11_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i52_LC_11_11_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i52_LC_11_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i52_LC_11_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9277),
            .lcout(\transmit_module.Y_DELTA_PATTERN_52 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23081),
            .ce(N__10035),
            .sr(N__21329));
    defparam \transmit_module.Y_DELTA_PATTERN_i50_LC_11_11_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i50_LC_11_11_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i50_LC_11_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i50_LC_11_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9262),
            .lcout(\transmit_module.Y_DELTA_PATTERN_50 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23081),
            .ce(N__10035),
            .sr(N__21329));
    defparam \transmit_module.Y_DELTA_PATTERN_i51_LC_11_11_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i51_LC_11_11_7 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i51_LC_11_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i51_LC_11_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9268),
            .lcout(\transmit_module.Y_DELTA_PATTERN_51 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23081),
            .ce(N__10035),
            .sr(N__21329));
    defparam \transmit_module.Y_DELTA_PATTERN_i33_LC_11_12_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i33_LC_11_12_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i33_LC_11_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i33_LC_11_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9343),
            .lcout(\transmit_module.Y_DELTA_PATTERN_33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23086),
            .ce(N__10028),
            .sr(N__21276));
    defparam \transmit_module.Y_DELTA_PATTERN_i81_LC_11_12_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i81_LC_11_12_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i81_LC_11_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i81_LC_11_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9331),
            .lcout(\transmit_module.Y_DELTA_PATTERN_81 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23086),
            .ce(N__10028),
            .sr(N__21276));
    defparam \transmit_module.Y_DELTA_PATTERN_i80_LC_11_12_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i80_LC_11_12_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i80_LC_11_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i80_LC_11_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9370),
            .lcout(\transmit_module.Y_DELTA_PATTERN_80 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23086),
            .ce(N__10028),
            .sr(N__21276));
    defparam \transmit_module.Y_DELTA_PATTERN_i49_LC_11_12_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i49_LC_11_12_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i49_LC_11_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i49_LC_11_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9364),
            .lcout(\transmit_module.Y_DELTA_PATTERN_49 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23086),
            .ce(N__10028),
            .sr(N__21276));
    defparam \transmit_module.Y_DELTA_PATTERN_i34_LC_11_12_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i34_LC_11_12_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i34_LC_11_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i34_LC_11_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9352),
            .lcout(\transmit_module.Y_DELTA_PATTERN_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23086),
            .ce(N__10028),
            .sr(N__21276));
    defparam \transmit_module.Y_DELTA_PATTERN_i71_LC_11_12_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i71_LC_11_12_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i71_LC_11_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i71_LC_11_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9337),
            .lcout(\transmit_module.Y_DELTA_PATTERN_71 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23086),
            .ce(N__10028),
            .sr(N__21276));
    defparam \transmit_module.Y_DELTA_PATTERN_i82_LC_11_12_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i82_LC_11_12_7 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i82_LC_11_12_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i82_LC_11_12_7  (
            .in0(N__9715),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.Y_DELTA_PATTERN_82 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23086),
            .ce(N__10028),
            .sr(N__21276));
    defparam \transmit_module.Y_DELTA_PATTERN_i69_LC_11_13_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i69_LC_11_13_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i69_LC_11_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i69_LC_11_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9484),
            .lcout(\transmit_module.Y_DELTA_PATTERN_69 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23077),
            .ce(N__10024),
            .sr(N__21331));
    defparam \transmit_module.Y_DELTA_PATTERN_i68_LC_11_13_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i68_LC_11_13_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i68_LC_11_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i68_LC_11_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9325),
            .lcout(\transmit_module.Y_DELTA_PATTERN_68 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23077),
            .ce(N__10024),
            .sr(N__21331));
    defparam \transmit_module.Y_DELTA_PATTERN_i78_LC_11_13_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i78_LC_11_13_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i78_LC_11_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i78_LC_11_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9301),
            .lcout(\transmit_module.Y_DELTA_PATTERN_78 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23077),
            .ce(N__10024),
            .sr(N__21331));
    defparam \transmit_module.Y_DELTA_PATTERN_i79_LC_11_13_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i79_LC_11_13_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i79_LC_11_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i79_LC_11_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9307),
            .lcout(\transmit_module.Y_DELTA_PATTERN_79 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23077),
            .ce(N__10024),
            .sr(N__21331));
    defparam \transmit_module.Y_DELTA_PATTERN_i70_LC_11_13_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i70_LC_11_13_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i70_LC_11_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i70_LC_11_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9490),
            .lcout(\transmit_module.Y_DELTA_PATTERN_70 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23077),
            .ce(N__10024),
            .sr(N__21331));
    defparam \transmit_module.Y_DELTA_PATTERN_i67_LC_11_13_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i67_LC_11_13_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i67_LC_11_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i67_LC_11_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9478),
            .lcout(\transmit_module.Y_DELTA_PATTERN_67 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23077),
            .ce(N__10024),
            .sr(N__21331));
    defparam \transmit_module.video_signal_controller.i1_2_lut_3_lut_LC_11_14_0 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_2_lut_3_lut_LC_11_14_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_2_lut_3_lut_LC_11_14_0 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \transmit_module.video_signal_controller.i1_2_lut_3_lut_LC_11_14_0  (
            .in0(N__9661),
            .in1(N__9391),
            .in2(_gnd_net_),
            .in3(N__9574),
            .lcout(\transmit_module.video_signal_controller.n1983 ),
            .ltout(\transmit_module.video_signal_controller.n1983_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1693_4_lut_LC_11_14_1 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1693_4_lut_LC_11_14_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1693_4_lut_LC_11_14_1 .LUT_INIT=16'b1010100010100000;
    LogicCell40 \transmit_module.video_signal_controller.i1693_4_lut_LC_11_14_1  (
            .in0(N__9690),
            .in1(N__9463),
            .in2(N__9457),
            .in3(N__9432),
            .lcout(\transmit_module.video_signal_controller.n2926 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1699_4_lut_LC_11_14_3 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1699_4_lut_LC_11_14_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1699_4_lut_LC_11_14_3 .LUT_INIT=16'b1110111011101100;
    LogicCell40 \transmit_module.video_signal_controller.i1699_4_lut_LC_11_14_3  (
            .in0(N__9612),
            .in1(N__10490),
            .in2(N__9640),
            .in3(N__9454),
            .lcout(\transmit_module.video_signal_controller.n2010 ),
            .ltout(\transmit_module.video_signal_controller.n2010_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1136_2_lut_LC_11_14_4 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1136_2_lut_LC_11_14_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1136_2_lut_LC_11_14_4 .LUT_INIT=16'b1100000011000000;
    LogicCell40 \transmit_module.video_signal_controller.i1136_2_lut_LC_11_14_4  (
            .in0(_gnd_net_),
            .in1(N__17401),
            .in2(N__9448),
            .in3(_gnd_net_),
            .lcout(\transmit_module.video_signal_controller.n2361 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i483_4_lut_LC_11_14_5 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i483_4_lut_LC_11_14_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i483_4_lut_LC_11_14_5 .LUT_INIT=16'b1110000010100000;
    LogicCell40 \transmit_module.video_signal_controller.i483_4_lut_LC_11_14_5  (
            .in0(N__9445),
            .in1(N__9439),
            .in2(N__9694),
            .in3(N__9433),
            .lcout(),
            .ltout(\transmit_module.video_signal_controller.n18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i2_4_lut_4_lut_LC_11_14_6 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i2_4_lut_4_lut_LC_11_14_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i2_4_lut_4_lut_LC_11_14_6 .LUT_INIT=16'b0000001111111110;
    LogicCell40 \transmit_module.video_signal_controller.i2_4_lut_4_lut_LC_11_14_6  (
            .in0(N__10491),
            .in1(N__9639),
            .in2(N__9424),
            .in3(N__9613),
            .lcout(\transmit_module.video_signal_controller.n7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_4_lut_adj_26_LC_11_15_1 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_4_lut_adj_26_LC_11_15_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_4_lut_adj_26_LC_11_15_1 .LUT_INIT=16'b1111111011110000;
    LogicCell40 \transmit_module.video_signal_controller.i1_4_lut_adj_26_LC_11_15_1  (
            .in0(N__9553),
            .in1(N__9420),
            .in2(N__9580),
            .in3(N__9394),
            .lcout(),
            .ltout(\transmit_module.video_signal_controller.n4_adj_617_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.VGA_HS_66_LC_11_15_2 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.VGA_HS_66_LC_11_15_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_HS_66_LC_11_15_2 .LUT_INIT=16'b1110111011101111;
    LogicCell40 \transmit_module.video_signal_controller.VGA_HS_66_LC_11_15_2  (
            .in0(N__9689),
            .in1(N__9532),
            .in2(N__9667),
            .in3(N__9664),
            .lcout(ADV_HSYNC_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22972),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i2_3_lut_rep_27_LC_11_15_5 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i2_3_lut_rep_27_LC_11_15_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i2_3_lut_rep_27_LC_11_15_5 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \transmit_module.video_signal_controller.i2_3_lut_rep_27_LC_11_15_5  (
            .in0(N__9629),
            .in1(N__9602),
            .in2(_gnd_net_),
            .in3(N__10485),
            .lcout(),
            .ltout(\transmit_module.video_signal_controller.n3794_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i2292_4_lut_LC_11_15_6 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i2292_4_lut_LC_11_15_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i2292_4_lut_LC_11_15_6 .LUT_INIT=16'b1111110011111000;
    LogicCell40 \transmit_module.video_signal_controller.i2292_4_lut_LC_11_15_6  (
            .in0(N__9586),
            .in1(N__9576),
            .in2(N__9556),
            .in3(N__9552),
            .lcout(\transmit_module.video_signal_controller.n3618 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.Y_DELTA_PATTERN_i60_LC_12_10_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i60_LC_12_10_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i60_LC_12_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i60_LC_12_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9526),
            .lcout(\transmit_module.Y_DELTA_PATTERN_60 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23082),
            .ce(N__10050),
            .sr(N__21319));
    defparam \transmit_module.Y_DELTA_PATTERN_i37_LC_12_10_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i37_LC_12_10_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i37_LC_12_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i37_LC_12_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9508),
            .lcout(\transmit_module.Y_DELTA_PATTERN_37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23082),
            .ce(N__10050),
            .sr(N__21319));
    defparam \transmit_module.Y_DELTA_PATTERN_i38_LC_12_10_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i38_LC_12_10_2 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i38_LC_12_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i38_LC_12_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9514),
            .lcout(\transmit_module.Y_DELTA_PATTERN_38 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23082),
            .ce(N__10050),
            .sr(N__21319));
    defparam \transmit_module.Y_DELTA_PATTERN_i58_LC_12_10_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i58_LC_12_10_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i58_LC_12_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i58_LC_12_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9748),
            .lcout(\transmit_module.Y_DELTA_PATTERN_58 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23082),
            .ce(N__10050),
            .sr(N__21319));
    defparam \transmit_module.Y_DELTA_PATTERN_i57_LC_12_10_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i57_LC_12_10_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i57_LC_12_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i57_LC_12_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9502),
            .lcout(\transmit_module.Y_DELTA_PATTERN_57 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23082),
            .ce(N__10050),
            .sr(N__21319));
    defparam \transmit_module.Y_DELTA_PATTERN_i59_LC_12_10_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i59_LC_12_10_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i59_LC_12_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i59_LC_12_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9754),
            .lcout(\transmit_module.Y_DELTA_PATTERN_59 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23082),
            .ce(N__10050),
            .sr(N__21319));
    defparam \transmit_module.Y_DELTA_PATTERN_i98_LC_12_11_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i98_LC_12_11_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i98_LC_12_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i98_LC_12_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9709),
            .lcout(\transmit_module.Y_DELTA_PATTERN_98 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22968),
            .ce(N__11065),
            .sr(N__21284));
    defparam \transmit_module.Y_DELTA_PATTERN_i85_LC_12_11_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i85_LC_12_11_2 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i85_LC_12_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i85_LC_12_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9736),
            .lcout(\transmit_module.Y_DELTA_PATTERN_85 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22968),
            .ce(N__11065),
            .sr(N__21284));
    defparam \transmit_module.Y_DELTA_PATTERN_i84_LC_12_11_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i84_LC_12_11_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i84_LC_12_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i84_LC_12_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9727),
            .lcout(\transmit_module.Y_DELTA_PATTERN_84 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22968),
            .ce(N__11065),
            .sr(N__21284));
    defparam \transmit_module.Y_DELTA_PATTERN_i83_LC_12_11_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i83_LC_12_11_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i83_LC_12_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i83_LC_12_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9721),
            .lcout(\transmit_module.Y_DELTA_PATTERN_83 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22968),
            .ce(N__11065),
            .sr(N__21284));
    defparam \transmit_module.Y_DELTA_PATTERN_i99_LC_12_12_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i99_LC_12_12_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i99_LC_12_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i99_LC_12_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17938),
            .lcout(\transmit_module.Y_DELTA_PATTERN_99 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23144),
            .ce(N__21478),
            .sr(N__21275));
    defparam \transmit_module.video_signal_controller.VGA_Y_i0_LC_12_13_0 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i0_LC_12_13_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i0_LC_12_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i0_LC_12_13_0  (
            .in0(_gnd_net_),
            .in1(N__11391),
            .in2(_gnd_net_),
            .in3(N__9703),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_0 ),
            .ltout(),
            .carryin(bfn_12_13_0_),
            .carryout(\transmit_module.video_signal_controller.n3290 ),
            .clk(N__23101),
            .ce(N__9778),
            .sr(N__9850));
    defparam \transmit_module.video_signal_controller.VGA_Y_i1_LC_12_13_1 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i1_LC_12_13_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i1_LC_12_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i1_LC_12_13_1  (
            .in0(_gnd_net_),
            .in1(N__11348),
            .in2(_gnd_net_),
            .in3(N__9700),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_1 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3290 ),
            .carryout(\transmit_module.video_signal_controller.n3291 ),
            .clk(N__23101),
            .ce(N__9778),
            .sr(N__9850));
    defparam \transmit_module.video_signal_controller.VGA_Y_i2_LC_12_13_2 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i2_LC_12_13_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i2_LC_12_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i2_LC_12_13_2  (
            .in0(_gnd_net_),
            .in1(N__10074),
            .in2(_gnd_net_),
            .in3(N__9697),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_2 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3291 ),
            .carryout(\transmit_module.video_signal_controller.n3292 ),
            .clk(N__23101),
            .ce(N__9778),
            .sr(N__9850));
    defparam \transmit_module.video_signal_controller.VGA_Y_i3_LC_12_13_3 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i3_LC_12_13_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i3_LC_12_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i3_LC_12_13_3  (
            .in0(_gnd_net_),
            .in1(N__11377),
            .in2(_gnd_net_),
            .in3(N__9817),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_3 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3292 ),
            .carryout(\transmit_module.video_signal_controller.n3293 ),
            .clk(N__23101),
            .ce(N__9778),
            .sr(N__9850));
    defparam \transmit_module.video_signal_controller.VGA_Y_i4_LC_12_13_4 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i4_LC_12_13_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i4_LC_12_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i4_LC_12_13_4  (
            .in0(_gnd_net_),
            .in1(N__11016),
            .in2(_gnd_net_),
            .in3(N__9814),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_4 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3293 ),
            .carryout(\transmit_module.video_signal_controller.n3294 ),
            .clk(N__23101),
            .ce(N__9778),
            .sr(N__9850));
    defparam \transmit_module.video_signal_controller.VGA_Y_i5_LC_12_13_5 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i5_LC_12_13_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i5_LC_12_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i5_LC_12_13_5  (
            .in0(_gnd_net_),
            .in1(N__10095),
            .in2(_gnd_net_),
            .in3(N__9811),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_5 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3294 ),
            .carryout(\transmit_module.video_signal_controller.n3295 ),
            .clk(N__23101),
            .ce(N__9778),
            .sr(N__9850));
    defparam \transmit_module.video_signal_controller.VGA_Y_i6_LC_12_13_6 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i6_LC_12_13_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i6_LC_12_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i6_LC_12_13_6  (
            .in0(_gnd_net_),
            .in1(N__10155),
            .in2(_gnd_net_),
            .in3(N__9808),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_6 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3295 ),
            .carryout(\transmit_module.video_signal_controller.n3296 ),
            .clk(N__23101),
            .ce(N__9778),
            .sr(N__9850));
    defparam \transmit_module.video_signal_controller.VGA_Y_i7_LC_12_13_7 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i7_LC_12_13_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i7_LC_12_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i7_LC_12_13_7  (
            .in0(_gnd_net_),
            .in1(N__10119),
            .in2(_gnd_net_),
            .in3(N__9805),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_7 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3296 ),
            .carryout(\transmit_module.video_signal_controller.n3297 ),
            .clk(N__23101),
            .ce(N__9778),
            .sr(N__9850));
    defparam \transmit_module.video_signal_controller.VGA_Y_i8_LC_12_14_0 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i8_LC_12_14_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i8_LC_12_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i8_LC_12_14_0  (
            .in0(_gnd_net_),
            .in1(N__10992),
            .in2(_gnd_net_),
            .in3(N__9802),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_8 ),
            .ltout(),
            .carryin(bfn_12_14_0_),
            .carryout(\transmit_module.video_signal_controller.n3298 ),
            .clk(N__22990),
            .ce(N__9782),
            .sr(N__9849));
    defparam \transmit_module.video_signal_controller.VGA_Y_i9_LC_12_14_1 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i9_LC_12_14_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i9_LC_12_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i9_LC_12_14_1  (
            .in0(_gnd_net_),
            .in1(N__10178),
            .in2(_gnd_net_),
            .in3(N__9799),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_9 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3298 ),
            .carryout(\transmit_module.video_signal_controller.n3299 ),
            .clk(N__22990),
            .ce(N__9782),
            .sr(N__9849));
    defparam \transmit_module.video_signal_controller.VGA_Y_i10_LC_12_14_2 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i10_LC_12_14_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i10_LC_12_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i10_LC_12_14_2  (
            .in0(_gnd_net_),
            .in1(N__11415),
            .in2(_gnd_net_),
            .in3(N__9796),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_10 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3299 ),
            .carryout(\transmit_module.video_signal_controller.n3300 ),
            .clk(N__22990),
            .ce(N__9782),
            .sr(N__9849));
    defparam \transmit_module.video_signal_controller.VGA_Y_i11_LC_12_14_3 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.VGA_Y_i11_LC_12_14_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i11_LC_12_14_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i11_LC_12_14_3  (
            .in0(N__10135),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9793),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22990),
            .ce(N__9782),
            .sr(N__9849));
    defparam \transmit_module.i2_3_lut_rep_20_LC_12_15_2 .C_ON=1'b0;
    defparam \transmit_module.i2_3_lut_rep_20_LC_12_15_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i2_3_lut_rep_20_LC_12_15_2 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \transmit_module.i2_3_lut_rep_20_LC_12_15_2  (
            .in0(N__10583),
            .in1(N__10609),
            .in2(_gnd_net_),
            .in3(N__10545),
            .lcout(\transmit_module.n3787 ),
            .ltout(\transmit_module.n3787_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i2_3_lut_LC_12_15_3 .C_ON=1'b0;
    defparam \transmit_module.i2_3_lut_LC_12_15_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i2_3_lut_LC_12_15_3 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \transmit_module.i2_3_lut_LC_12_15_3  (
            .in0(_gnd_net_),
            .in1(N__21120),
            .in2(N__9838),
            .in3(N__18298),
            .lcout(\transmit_module.n2093 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.old_VGA_HS_40_LC_12_15_4 .C_ON=1'b0;
    defparam \transmit_module.old_VGA_HS_40_LC_12_15_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.old_VGA_HS_40_LC_12_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.old_VGA_HS_40_LC_12_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10547),
            .lcout(\transmit_module.old_VGA_HS ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22961),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1_3_lut_LC_12_15_5 .C_ON=1'b0;
    defparam \transmit_module.i1_3_lut_LC_12_15_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1_3_lut_LC_12_15_5 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \transmit_module.i1_3_lut_LC_12_15_5  (
            .in0(N__21118),
            .in1(N__17933),
            .in2(_gnd_net_),
            .in3(N__18989),
            .lcout(\transmit_module.n2061 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i246_2_lut_4_lut_rep_30_LC_12_15_7 .C_ON=1'b0;
    defparam \transmit_module.i246_2_lut_4_lut_rep_30_LC_12_15_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i246_2_lut_4_lut_rep_30_LC_12_15_7 .LUT_INIT=16'b1101110011001100;
    LogicCell40 \transmit_module.i246_2_lut_4_lut_rep_30_LC_12_15_7  (
            .in0(N__10546),
            .in1(N__21119),
            .in2(N__10615),
            .in3(N__10584),
            .lcout(\transmit_module.n3797 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.Y_DELTA_PATTERN_i7_LC_12_16_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i7_LC_12_16_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i7_LC_12_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i7_LC_12_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11533),
            .lcout(\transmit_module.Y_DELTA_PATTERN_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22938),
            .ce(N__21449),
            .sr(N__21195));
    defparam \transmit_module.Y_DELTA_PATTERN_i5_LC_12_16_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i5_LC_12_16_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i5_LC_12_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i5_LC_12_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9829),
            .lcout(\transmit_module.Y_DELTA_PATTERN_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22938),
            .ce(N__21449),
            .sr(N__21195));
    defparam \transmit_module.Y_DELTA_PATTERN_i6_LC_12_16_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i6_LC_12_16_2 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i6_LC_12_16_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i6_LC_12_16_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9835),
            .lcout(\transmit_module.Y_DELTA_PATTERN_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22938),
            .ce(N__21449),
            .sr(N__21195));
    defparam \transmit_module.Y_DELTA_PATTERN_i4_LC_12_16_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i4_LC_12_16_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i4_LC_12_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i4_LC_12_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9823),
            .lcout(\transmit_module.Y_DELTA_PATTERN_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22938),
            .ce(N__21449),
            .sr(N__21195));
    defparam \transmit_module.Y_DELTA_PATTERN_i2_LC_12_16_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i2_LC_12_16_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i2_LC_12_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i2_LC_12_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9919),
            .lcout(\transmit_module.Y_DELTA_PATTERN_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22938),
            .ce(N__21449),
            .sr(N__21195));
    defparam \transmit_module.Y_DELTA_PATTERN_i3_LC_12_16_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i3_LC_12_16_7 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i3_LC_12_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i3_LC_12_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9925),
            .lcout(\transmit_module.Y_DELTA_PATTERN_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22938),
            .ce(N__21449),
            .sr(N__21195));
    defparam \transmit_module.ADDR_Y_COMPONENT__i11_LC_12_17_0 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i11_LC_12_17_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i11_LC_12_17_0 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i11_LC_12_17_0  (
            .in0(_gnd_net_),
            .in1(N__23601),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23087),
            .ce(N__17743),
            .sr(N__21300));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_LC_12_18_6 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_LC_12_18_6 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_LC_12_18_6 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_LC_12_18_6  (
            .in0(N__23630),
            .in1(N__9913),
            .in2(N__22233),
            .in3(N__9901),
            .lcout(\line_buffer.n3764 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2321_3_lut_LC_12_21_6 .C_ON=1'b0;
    defparam \line_buffer.i2321_3_lut_LC_12_21_6 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2321_3_lut_LC_12_21_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \line_buffer.i2321_3_lut_LC_12_21_6  (
            .in0(N__23639),
            .in1(N__9889),
            .in2(_gnd_net_),
            .in3(N__9877),
            .lcout(\line_buffer.n3647 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.Y__i0_LC_13_10_0 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i0_LC_13_10_0 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i0_LC_13_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i0_LC_13_10_0  (
            .in0(_gnd_net_),
            .in1(N__11178),
            .in2(_gnd_net_),
            .in3(N__9865),
            .lcout(\receive_module.rx_counter.Y_0 ),
            .ltout(),
            .carryin(bfn_13_10_0_),
            .carryout(\receive_module.rx_counter.n3271 ),
            .clk(N__20141),
            .ce(N__13092),
            .sr(N__21947));
    defparam \receive_module.rx_counter.Y__i1_LC_13_10_1 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i1_LC_13_10_1 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i1_LC_13_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i1_LC_13_10_1  (
            .in0(_gnd_net_),
            .in1(N__11247),
            .in2(_gnd_net_),
            .in3(N__9862),
            .lcout(\receive_module.rx_counter.Y_1 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3271 ),
            .carryout(\receive_module.rx_counter.n3272 ),
            .clk(N__20141),
            .ce(N__13092),
            .sr(N__21947));
    defparam \receive_module.rx_counter.Y__i2_LC_13_10_2 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i2_LC_13_10_2 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i2_LC_13_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i2_LC_13_10_2  (
            .in0(_gnd_net_),
            .in1(N__11266),
            .in2(_gnd_net_),
            .in3(N__9859),
            .lcout(\receive_module.rx_counter.Y_2 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3272 ),
            .carryout(\receive_module.rx_counter.n3273 ),
            .clk(N__20141),
            .ce(N__13092),
            .sr(N__21947));
    defparam \receive_module.rx_counter.Y__i3_LC_13_10_3 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i3_LC_13_10_3 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i3_LC_13_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i3_LC_13_10_3  (
            .in0(_gnd_net_),
            .in1(N__11284),
            .in2(_gnd_net_),
            .in3(N__9856),
            .lcout(\receive_module.rx_counter.Y_3 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3273 ),
            .carryout(\receive_module.rx_counter.n3274 ),
            .clk(N__20141),
            .ce(N__13092),
            .sr(N__21947));
    defparam \receive_module.rx_counter.Y__i4_LC_13_10_4 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i4_LC_13_10_4 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i4_LC_13_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i4_LC_13_10_4  (
            .in0(_gnd_net_),
            .in1(N__13122),
            .in2(_gnd_net_),
            .in3(N__9853),
            .lcout(\receive_module.rx_counter.Y_4 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3274 ),
            .carryout(\receive_module.rx_counter.n3275 ),
            .clk(N__20141),
            .ce(N__13092),
            .sr(N__21947));
    defparam \receive_module.rx_counter.Y__i5_LC_13_10_5 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i5_LC_13_10_5 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i5_LC_13_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i5_LC_13_10_5  (
            .in0(_gnd_net_),
            .in1(N__11227),
            .in2(_gnd_net_),
            .in3(N__9940),
            .lcout(\receive_module.rx_counter.Y_5 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3275 ),
            .carryout(\receive_module.rx_counter.n3276 ),
            .clk(N__20141),
            .ce(N__13092),
            .sr(N__21947));
    defparam \receive_module.rx_counter.Y__i6_LC_13_10_6 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i6_LC_13_10_6 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i6_LC_13_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i6_LC_13_10_6  (
            .in0(_gnd_net_),
            .in1(N__11212),
            .in2(_gnd_net_),
            .in3(N__9937),
            .lcout(\receive_module.rx_counter.Y_6 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3276 ),
            .carryout(\receive_module.rx_counter.n3277 ),
            .clk(N__20141),
            .ce(N__13092),
            .sr(N__21947));
    defparam \receive_module.rx_counter.Y__i7_LC_13_10_7 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i7_LC_13_10_7 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i7_LC_13_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i7_LC_13_10_7  (
            .in0(_gnd_net_),
            .in1(N__13164),
            .in2(_gnd_net_),
            .in3(N__9934),
            .lcout(\receive_module.rx_counter.Y_7 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3277 ),
            .carryout(\receive_module.rx_counter.n3278 ),
            .clk(N__20141),
            .ce(N__13092),
            .sr(N__21947));
    defparam \receive_module.rx_counter.Y__i8_LC_13_11_0 .C_ON=1'b0;
    defparam \receive_module.rx_counter.Y__i8_LC_13_11_0 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i8_LC_13_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i8_LC_13_11_0  (
            .in0(_gnd_net_),
            .in1(N__16862),
            .in2(_gnd_net_),
            .in3(N__9931),
            .lcout(\receive_module.rx_counter.Y_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20145),
            .ce(N__13096),
            .sr(N__21956));
    defparam \transmit_module.ADDR_Y_COMPONENT__i7_LC_13_12_1 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i7_LC_13_12_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i7_LC_13_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i7_LC_13_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13543),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23274),
            .ce(N__17774),
            .sr(N__21261));
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_18_LC_13_13_0 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_18_LC_13_13_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_18_LC_13_13_0 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \transmit_module.video_signal_controller.i1_2_lut_rep_18_LC_13_13_0  (
            .in0(N__10118),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10988),
            .lcout(\transmit_module.video_signal_controller.n3785 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i2_2_lut_3_lut_LC_13_13_1 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i2_2_lut_3_lut_LC_13_13_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i2_2_lut_3_lut_LC_13_13_1 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \transmit_module.video_signal_controller.i2_2_lut_3_lut_LC_13_13_1  (
            .in0(N__10179),
            .in1(N__10981),
            .in2(_gnd_net_),
            .in3(N__10117),
            .lcout(\transmit_module.video_signal_controller.n8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_19_LC_13_13_2 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_19_LC_13_13_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_19_LC_13_13_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \transmit_module.video_signal_controller.i1_2_lut_rep_19_LC_13_13_2  (
            .in0(_gnd_net_),
            .in1(N__11344),
            .in2(_gnd_net_),
            .in3(N__10072),
            .lcout(),
            .ltout(\transmit_module.video_signal_controller.n3786_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_4_lut_adj_24_LC_13_13_3 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_4_lut_adj_24_LC_13_13_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_4_lut_adj_24_LC_13_13_3 .LUT_INIT=16'b1111111110101000;
    LogicCell40 \transmit_module.video_signal_controller.i1_4_lut_adj_24_LC_13_13_3  (
            .in0(N__11011),
            .in1(N__11379),
            .in2(N__9928),
            .in3(N__10188),
            .lcout(),
            .ltout(\transmit_module.video_signal_controller.n7_adj_615_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i5_4_lut_LC_13_13_4 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i5_4_lut_LC_13_13_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i5_4_lut_LC_13_13_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \transmit_module.video_signal_controller.i5_4_lut_LC_13_13_4  (
            .in0(N__10094),
            .in1(N__10210),
            .in2(N__10204),
            .in3(N__10154),
            .lcout(\transmit_module.video_signal_controller.VGA_VISIBLE_N_578 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_2_lut_3_lut_adj_27_LC_13_13_5 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_2_lut_3_lut_adj_27_LC_13_13_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_2_lut_3_lut_adj_27_LC_13_13_5 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \transmit_module.video_signal_controller.i1_2_lut_3_lut_adj_27_LC_13_13_5  (
            .in0(N__10073),
            .in1(_gnd_net_),
            .in2(N__11352),
            .in3(N__11378),
            .lcout(),
            .ltout(\transmit_module.video_signal_controller.n2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i2_4_lut_LC_13_13_6 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i2_4_lut_LC_13_13_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i2_4_lut_LC_13_13_6 .LUT_INIT=16'b1000100010000000;
    LogicCell40 \transmit_module.video_signal_controller.i2_4_lut_LC_13_13_6  (
            .in0(N__10093),
            .in1(N__10153),
            .in2(N__10201),
            .in3(N__11012),
            .lcout(),
            .ltout(\transmit_module.video_signal_controller.n3577_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_4_lut_LC_13_13_7 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_4_lut_LC_13_13_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_4_lut_LC_13_13_7 .LUT_INIT=16'b1111111110101000;
    LogicCell40 \transmit_module.video_signal_controller.i1_4_lut_LC_13_13_7  (
            .in0(N__10180),
            .in1(N__10198),
            .in2(N__10192),
            .in3(N__10189),
            .lcout(\transmit_module.video_signal_controller.n3486 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.VGA_VISIBLE_Y_64_LC_13_14_2 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.VGA_VISIBLE_Y_64_LC_13_14_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_VISIBLE_Y_64_LC_13_14_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \transmit_module.video_signal_controller.VGA_VISIBLE_Y_64_LC_13_14_2  (
            .in0(_gnd_net_),
            .in1(N__10521),
            .in2(_gnd_net_),
            .in3(N__10455),
            .lcout(\transmit_module.VGA_VISIBLE_Y ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23273),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_2_lut_LC_13_14_3 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_2_lut_LC_13_14_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_2_lut_LC_13_14_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \transmit_module.video_signal_controller.i1_2_lut_LC_13_14_3  (
            .in0(_gnd_net_),
            .in1(N__10133),
            .in2(_gnd_net_),
            .in3(N__11414),
            .lcout(\transmit_module.video_signal_controller.n3485 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i2288_2_lut_LC_13_14_5 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i2288_2_lut_LC_13_14_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i2288_2_lut_LC_13_14_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \transmit_module.video_signal_controller.i2288_2_lut_LC_13_14_5  (
            .in0(_gnd_net_),
            .in1(N__10177),
            .in2(_gnd_net_),
            .in3(N__10156),
            .lcout(\transmit_module.video_signal_controller.n3614 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i2306_4_lut_LC_13_14_6 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i2306_4_lut_LC_13_14_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i2306_4_lut_LC_13_14_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \transmit_module.video_signal_controller.i2306_4_lut_LC_13_14_6  (
            .in0(N__10134),
            .in1(N__10120),
            .in2(N__10099),
            .in3(N__10075),
            .lcout(\transmit_module.video_signal_controller.n3632 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i246_2_lut_4_lut_rep_31_LC_13_15_0 .C_ON=1'b0;
    defparam \transmit_module.i246_2_lut_4_lut_rep_31_LC_13_15_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i246_2_lut_4_lut_rep_31_LC_13_15_0 .LUT_INIT=16'b1101110011001100;
    LogicCell40 \transmit_module.i246_2_lut_4_lut_rep_31_LC_13_15_0  (
            .in0(N__10557),
            .in1(N__21059),
            .in2(N__10594),
            .in3(N__10614),
            .lcout(\transmit_module.n3798 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i5_3_lut_LC_13_15_1 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i5_3_lut_LC_13_15_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i5_3_lut_LC_13_15_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_12_i5_3_lut_LC_13_15_1  (
            .in0(N__17905),
            .in1(N__10963),
            .in2(_gnd_net_),
            .in3(N__13338),
            .lcout(\transmit_module.n112 ),
            .ltout(\transmit_module.n112_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1603_4_lut_LC_13_15_2 .C_ON=1'b0;
    defparam \transmit_module.i1603_4_lut_LC_13_15_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1603_4_lut_LC_13_15_2 .LUT_INIT=16'b0101000001000100;
    LogicCell40 \transmit_module.i1603_4_lut_LC_13_15_2  (
            .in0(N__21004),
            .in1(N__11317),
            .in2(N__10837),
            .in3(N__18988),
            .lcout(n24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i246_2_lut_4_lut_LC_13_15_3 .C_ON=1'b0;
    defparam \transmit_module.i246_2_lut_4_lut_LC_13_15_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i246_2_lut_4_lut_LC_13_15_3 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \transmit_module.i246_2_lut_4_lut_LC_13_15_3  (
            .in0(N__10613),
            .in1(N__10590),
            .in2(N__21167),
            .in3(N__10556),
            .lcout(\transmit_module.n2147 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.VGA_VISIBLE_65_LC_13_15_5 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.VGA_VISIBLE_65_LC_13_15_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_VISIBLE_65_LC_13_15_5 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \transmit_module.video_signal_controller.VGA_VISIBLE_65_LC_13_15_5  (
            .in0(N__10525),
            .in1(N__10510),
            .in2(N__10498),
            .in3(N__10459),
            .lcout(\transmit_module.VGA_VISIBLE ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23203),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i6_3_lut_LC_13_15_6 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i6_3_lut_LC_13_15_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i6_3_lut_LC_13_15_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_12_i6_3_lut_LC_13_15_6  (
            .in0(N__17906),
            .in1(N__10957),
            .in2(_gnd_net_),
            .in3(N__13305),
            .lcout(\transmit_module.n111 ),
            .ltout(\transmit_module.n111_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1604_4_lut_LC_13_15_7 .C_ON=1'b0;
    defparam \transmit_module.i1604_4_lut_LC_13_15_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1604_4_lut_LC_13_15_7 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \transmit_module.i1604_4_lut_LC_13_15_7  (
            .in0(N__18987),
            .in1(N__21005),
            .in2(N__10444),
            .in3(N__11295),
            .lcout(n23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.ADDR_Y_COMPONENT__i12_LC_13_16_0 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i12_LC_13_16_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i12_LC_13_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i12_LC_13_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22172),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23130),
            .ce(N__17762),
            .sr(N__21050));
    defparam \transmit_module.ADDR_Y_COMPONENT__i1_LC_13_16_1 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i1_LC_13_16_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i1_LC_13_16_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i1_LC_13_16_1  (
            .in0(N__13390),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23130),
            .ce(N__17762),
            .sr(N__21050));
    defparam \transmit_module.ADDR_Y_COMPONENT__i10_LC_13_16_2 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i10_LC_13_16_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i10_LC_13_16_2 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i10_LC_13_16_2  (
            .in0(_gnd_net_),
            .in1(N__13498),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23130),
            .ce(N__17762),
            .sr(N__21050));
    defparam \transmit_module.ADDR_Y_COMPONENT__i4_LC_13_16_6 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i4_LC_13_16_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i4_LC_13_16_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i4_LC_13_16_6  (
            .in0(N__13342),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23130),
            .ce(N__17762),
            .sr(N__21050));
    defparam \transmit_module.ADDR_Y_COMPONENT__i5_LC_13_16_7 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i5_LC_13_16_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i5_LC_13_16_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i5_LC_13_16_7  (
            .in0(N__13306),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23130),
            .ce(N__17762),
            .sr(N__21050));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2422_LC_13_17_6 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2422_LC_13_17_6 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2422_LC_13_17_6 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_2422_LC_13_17_6  (
            .in0(N__23574),
            .in1(N__10951),
            .in2(N__22232),
            .in3(N__10936),
            .lcout(\line_buffer.n3752 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n3764_bdd_4_lut_LC_13_18_6 .C_ON=1'b0;
    defparam \line_buffer.n3764_bdd_4_lut_LC_13_18_6 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3764_bdd_4_lut_LC_13_18_6 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \line_buffer.n3764_bdd_4_lut_LC_13_18_6  (
            .in0(N__10921),
            .in1(N__22215),
            .in2(N__10906),
            .in3(N__10885),
            .lcout(\line_buffer.n3767 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2320_3_lut_LC_13_21_1 .C_ON=1'b0;
    defparam \line_buffer.i2320_3_lut_LC_13_21_1 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2320_3_lut_LC_13_21_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \line_buffer.i2320_3_lut_LC_13_21_1  (
            .in0(N__23640),
            .in1(N__10879),
            .in2(_gnd_net_),
            .in3(N__10864),
            .lcout(),
            .ltout(\line_buffer.n3646_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_2397_LC_13_21_2 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_2397_LC_13_21_2 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_2397_LC_13_21_2 .LUT_INIT=16'b1110110001100100;
    LogicCell40 \line_buffer.TX_ADDR_12__bdd_4_lut_2397_LC_13_21_2  (
            .in0(N__21683),
            .in1(N__22234),
            .in2(N__10846),
            .in3(N__10843),
            .lcout(\line_buffer.n3722 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i2_2_lut_LC_14_10_0 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i2_2_lut_LC_14_10_0 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i2_2_lut_LC_14_10_0 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \receive_module.rx_counter.i2_2_lut_LC_14_10_0  (
            .in0(N__13121),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13160),
            .lcout(\receive_module.rx_counter.n10_adj_610 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i1_2_lut_adj_20_LC_14_10_1 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i1_2_lut_adj_20_LC_14_10_1 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i1_2_lut_adj_20_LC_14_10_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \receive_module.rx_counter.i1_2_lut_adj_20_LC_14_10_1  (
            .in0(N__11282),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13120),
            .lcout(\receive_module.rx_counter.n4_adj_604 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i6_4_lut_LC_14_10_2 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i6_4_lut_LC_14_10_2 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i6_4_lut_LC_14_10_2 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \receive_module.rx_counter.i6_4_lut_LC_14_10_2  (
            .in0(N__11246),
            .in1(N__11283),
            .in2(N__16863),
            .in3(N__11265),
            .lcout(\receive_module.rx_counter.n14_adj_611 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i592_2_lut_rep_24_LC_14_10_3 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i592_2_lut_rep_24_LC_14_10_3 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i592_2_lut_rep_24_LC_14_10_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \receive_module.rx_counter.i592_2_lut_rep_24_LC_14_10_3  (
            .in0(_gnd_net_),
            .in1(N__11210),
            .in2(_gnd_net_),
            .in3(N__11225),
            .lcout(\receive_module.rx_counter.n3791 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i2_4_lut_adj_21_LC_14_10_4 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i2_4_lut_adj_21_LC_14_10_4 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i2_4_lut_adj_21_LC_14_10_4 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \receive_module.rx_counter.i2_4_lut_adj_21_LC_14_10_4  (
            .in0(N__11176),
            .in1(N__11281),
            .in2(N__11248),
            .in3(N__11263),
            .lcout(\receive_module.rx_counter.n3551 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i2_3_lut_LC_14_10_5 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i2_3_lut_LC_14_10_5 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i2_3_lut_LC_14_10_5 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \receive_module.rx_counter.i2_3_lut_LC_14_10_5  (
            .in0(N__11264),
            .in1(N__11177),
            .in2(_gnd_net_),
            .in3(N__11245),
            .lcout(\receive_module.rx_counter.n3548 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i1_2_lut_3_lut_LC_14_10_6 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i1_2_lut_3_lut_LC_14_10_6 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i1_2_lut_3_lut_LC_14_10_6 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \receive_module.rx_counter.i1_2_lut_3_lut_LC_14_10_6  (
            .in0(N__11226),
            .in1(N__13159),
            .in2(_gnd_net_),
            .in3(N__11211),
            .lcout(),
            .ltout(\receive_module.rx_counter.n5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i3_4_lut_LC_14_10_7 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i3_4_lut_LC_14_10_7 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i3_4_lut_LC_14_10_7 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \receive_module.rx_counter.i3_4_lut_LC_14_10_7  (
            .in0(N__16858),
            .in1(N__11194),
            .in2(N__11188),
            .in3(N__11185),
            .lcout(\receive_module.rx_counter.n3575 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.SYNC_46_LC_14_11_3 .C_ON=1'b0;
    defparam \receive_module.rx_counter.SYNC_46_LC_14_11_3 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.SYNC_46_LC_14_11_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \receive_module.rx_counter.SYNC_46_LC_14_11_3  (
            .in0(N__11179),
            .in1(N__11158),
            .in2(N__11152),
            .in3(N__13141),
            .lcout(RX_TX_SYNC),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20142),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i8_3_lut_LC_14_11_5 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i8_3_lut_LC_14_11_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i8_3_lut_LC_14_11_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_12_i8_3_lut_LC_14_11_5  (
            .in0(N__17927),
            .in1(N__11143),
            .in2(_gnd_net_),
            .in3(N__13545),
            .lcout(\transmit_module.n109 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.X_DELTA_PATTERN_i0_LC_14_12_0 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i0_LC_14_12_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i0_LC_14_12_0 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i0_LC_14_12_0  (
            .in0(_gnd_net_),
            .in1(N__11137),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.X_DELTA_PATTERN_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23143),
            .ce(N__11123),
            .sr(N__11064));
    defparam \transmit_module.video_signal_controller.i2300_2_lut_LC_14_13_0 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i2300_2_lut_LC_14_13_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i2300_2_lut_LC_14_13_0 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \transmit_module.video_signal_controller.i2300_2_lut_LC_14_13_0  (
            .in0(N__11017),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10993),
            .lcout(),
            .ltout(\transmit_module.video_signal_controller.n3626_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i7_4_lut_LC_14_13_1 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i7_4_lut_LC_14_13_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i7_4_lut_LC_14_13_1 .LUT_INIT=16'b0000001100000010;
    LogicCell40 \transmit_module.video_signal_controller.i7_4_lut_LC_14_13_1  (
            .in0(N__11398),
            .in1(N__11380),
            .in2(N__11356),
            .in3(N__11353),
            .lcout(\transmit_module.video_signal_controller.n18_adj_616 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i0_LC_14_13_2 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i0_LC_14_13_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i0_LC_14_13_2 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \transmit_module.BRAM_ADDR__i0_LC_14_13_2  (
            .in0(N__19081),
            .in1(N__12078),
            .in2(N__21233),
            .in3(N__12051),
            .lcout(\transmit_module.TX_ADDR_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23100),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i7_LC_14_13_4 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i7_LC_14_13_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i7_LC_14_13_4 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \transmit_module.BRAM_ADDR__i7_LC_14_13_4  (
            .in0(N__19082),
            .in1(N__12801),
            .in2(N__21234),
            .in3(N__12777),
            .lcout(\transmit_module.TX_ADDR_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23100),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i5_LC_14_13_7 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i5_LC_14_13_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i5_LC_14_13_7 .LUT_INIT=16'b0010001100100000;
    LogicCell40 \transmit_module.BRAM_ADDR__i5_LC_14_13_7  (
            .in0(N__11326),
            .in1(N__21131),
            .in2(N__19099),
            .in3(N__11296),
            .lcout(\transmit_module.TX_ADDR_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23100),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i2_LC_14_14_0 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i2_LC_14_14_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i2_LC_14_14_0 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \transmit_module.BRAM_ADDR__i2_LC_14_14_0  (
            .in0(N__19078),
            .in1(N__18577),
            .in2(N__21259),
            .in3(N__18556),
            .lcout(\transmit_module.TX_ADDR_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22989),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_14_i5_3_lut_LC_14_14_1 .C_ON=1'b0;
    defparam \transmit_module.mux_14_i5_3_lut_LC_14_14_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_14_i5_3_lut_LC_14_14_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \transmit_module.mux_14_i5_3_lut_LC_14_14_1  (
            .in0(N__13337),
            .in1(N__18273),
            .in2(_gnd_net_),
            .in3(N__13315),
            .lcout(\transmit_module.n143 ),
            .ltout(\transmit_module.n143_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i4_LC_14_14_2 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i4_LC_14_14_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i4_LC_14_14_2 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \transmit_module.BRAM_ADDR__i4_LC_14_14_2  (
            .in0(N__19079),
            .in1(N__21051),
            .in2(N__11305),
            .in3(N__11302),
            .lcout(\transmit_module.TX_ADDR_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22989),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_14_i6_3_lut_LC_14_14_3 .C_ON=1'b0;
    defparam \transmit_module.mux_14_i6_3_lut_LC_14_14_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_14_i6_3_lut_LC_14_14_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \transmit_module.mux_14_i6_3_lut_LC_14_14_3  (
            .in0(N__13297),
            .in1(N__18274),
            .in2(_gnd_net_),
            .in3(N__13276),
            .lcout(\transmit_module.n142 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i1_LC_14_14_4 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i1_LC_14_14_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i1_LC_14_14_4 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \transmit_module.BRAM_ADDR__i1_LC_14_14_4  (
            .in0(N__19077),
            .in1(N__11802),
            .in2(N__21258),
            .in3(N__11812),
            .lcout(\transmit_module.TX_ADDR_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22989),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_14_i7_3_lut_LC_14_14_5 .C_ON=1'b0;
    defparam \transmit_module.mux_14_i7_3_lut_LC_14_14_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_14_i7_3_lut_LC_14_14_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_14_i7_3_lut_LC_14_14_5  (
            .in0(N__18300),
            .in1(N__13258),
            .in2(_gnd_net_),
            .in3(N__13234),
            .lcout(\transmit_module.n141 ),
            .ltout(\transmit_module.n141_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i6_LC_14_14_6 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i6_LC_14_14_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i6_LC_14_14_6 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \transmit_module.BRAM_ADDR__i6_LC_14_14_6  (
            .in0(N__19080),
            .in1(N__21052),
            .in2(N__11470),
            .in3(N__13053),
            .lcout(\transmit_module.TX_ADDR_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22989),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_14_i8_3_lut_LC_14_14_7 .C_ON=1'b0;
    defparam \transmit_module.mux_14_i8_3_lut_LC_14_14_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_14_i8_3_lut_LC_14_14_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \transmit_module.mux_14_i8_3_lut_LC_14_14_7  (
            .in0(N__18301),
            .in1(_gnd_net_),
            .in2(N__13546),
            .in3(N__13513),
            .lcout(\transmit_module.n140 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_14_i11_3_lut_LC_14_15_0 .C_ON=1'b0;
    defparam \transmit_module.mux_14_i11_3_lut_LC_14_15_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_14_i11_3_lut_LC_14_15_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_14_i11_3_lut_LC_14_15_0  (
            .in0(N__18269),
            .in1(N__13496),
            .in2(_gnd_net_),
            .in3(N__13477),
            .lcout(\transmit_module.n137 ),
            .ltout(\transmit_module.n137_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i10_LC_14_15_1 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i10_LC_14_15_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i10_LC_14_15_1 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \transmit_module.BRAM_ADDR__i10_LC_14_15_1  (
            .in0(N__19023),
            .in1(N__21003),
            .in2(N__11467),
            .in3(N__12495),
            .lcout(\transmit_module.TX_ADDR_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23107),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i2_3_lut_LC_14_15_2 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i2_3_lut_LC_14_15_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i2_3_lut_LC_14_15_2 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \transmit_module.mux_12_i2_3_lut_LC_14_15_2  (
            .in0(N__13385),
            .in1(_gnd_net_),
            .in2(N__11464),
            .in3(N__17882),
            .lcout(\transmit_module.n115 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i11_3_lut_LC_14_15_3 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i11_3_lut_LC_14_15_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i11_3_lut_LC_14_15_3 .LUT_INIT=16'b1011100010111000;
    LogicCell40 \transmit_module.mux_12_i11_3_lut_LC_14_15_3  (
            .in0(N__13497),
            .in1(N__17881),
            .in2(N__11455),
            .in3(_gnd_net_),
            .lcout(\transmit_module.n106 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_14_i1_3_lut_LC_14_15_4 .C_ON=1'b0;
    defparam \transmit_module.mux_14_i1_3_lut_LC_14_15_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_14_i1_3_lut_LC_14_15_4 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \transmit_module.mux_14_i1_3_lut_LC_14_15_4  (
            .in0(N__13399),
            .in1(_gnd_net_),
            .in2(N__18299),
            .in3(N__13454),
            .lcout(\transmit_module.n147 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.VGA_VS_67_LC_14_15_5 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.VGA_VS_67_LC_14_15_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_VS_67_LC_14_15_5 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_VS_67_LC_14_15_5  (
            .in0(N__11446),
            .in1(N__11440),
            .in2(N__11431),
            .in3(N__11422),
            .lcout(ADV_VSYNC_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23107),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_14_i2_3_lut_LC_14_15_6 .C_ON=1'b0;
    defparam \transmit_module.mux_14_i2_3_lut_LC_14_15_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_14_i2_3_lut_LC_14_15_6 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \transmit_module.mux_14_i2_3_lut_LC_14_15_6  (
            .in0(N__13384),
            .in1(_gnd_net_),
            .in2(N__13363),
            .in3(N__18294),
            .lcout(\transmit_module.n146 ),
            .ltout(\transmit_module.n146_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1600_4_lut_LC_14_15_7 .C_ON=1'b0;
    defparam \transmit_module.i1600_4_lut_LC_14_15_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1600_4_lut_LC_14_15_7 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \transmit_module.i1600_4_lut_LC_14_15_7  (
            .in0(N__19022),
            .in1(N__21002),
            .in2(N__11806),
            .in3(N__11803),
            .lcout(n27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.Y_DELTA_PATTERN_i0_LC_14_16_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i0_LC_14_16_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i0_LC_14_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i0_LC_14_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11545),
            .lcout(\transmit_module.Y_DELTA_PATTERN_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22932),
            .ce(N__21459),
            .sr(N__21048));
    defparam \transmit_module.Y_DELTA_PATTERN_i9_LC_14_16_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i9_LC_14_16_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i9_LC_14_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i9_LC_14_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11524),
            .lcout(\transmit_module.Y_DELTA_PATTERN_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22932),
            .ce(N__21459),
            .sr(N__21048));
    defparam \transmit_module.Y_DELTA_PATTERN_i1_LC_14_16_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i1_LC_14_16_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i1_LC_14_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i1_LC_14_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11554),
            .lcout(\transmit_module.Y_DELTA_PATTERN_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22932),
            .ce(N__21459),
            .sr(N__21048));
    defparam \transmit_module.Y_DELTA_PATTERN_i8_LC_14_16_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i8_LC_14_16_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i8_LC_14_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i8_LC_14_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11539),
            .lcout(\transmit_module.Y_DELTA_PATTERN_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22932),
            .ce(N__21459),
            .sr(N__21048));
    defparam \transmit_module.Y_DELTA_PATTERN_i10_LC_14_16_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i10_LC_14_16_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i10_LC_14_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i10_LC_14_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19471),
            .lcout(\transmit_module.Y_DELTA_PATTERN_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22932),
            .ce(N__21459),
            .sr(N__21048));
    defparam \transmit_module.mux_12_i7_3_lut_LC_14_17_3 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i7_3_lut_LC_14_17_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i7_3_lut_LC_14_17_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_12_i7_3_lut_LC_14_17_3  (
            .in0(N__17883),
            .in1(N__12505),
            .in2(_gnd_net_),
            .in3(N__13266),
            .lcout(\transmit_module.n110 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n3752_bdd_4_lut_LC_14_17_4 .C_ON=1'b0;
    defparam \line_buffer.n3752_bdd_4_lut_LC_14_17_4 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3752_bdd_4_lut_LC_14_17_4 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \line_buffer.n3752_bdd_4_lut_LC_14_17_4  (
            .in0(N__11518),
            .in1(N__22125),
            .in2(N__11497),
            .in3(N__11476),
            .lcout(\line_buffer.n3755 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.ADDR_Y_COMPONENT__i6_LC_14_18_1 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i6_LC_14_18_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i6_LC_14_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i6_LC_14_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13267),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22979),
            .ce(N__17770),
            .sr(N__21117));
    defparam \transmit_module.ADDR_Y_COMPONENT__i0_LC_14_18_2 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i0_LC_14_18_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i0_LC_14_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i0_LC_14_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13456),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22979),
            .ce(N__17770),
            .sr(N__21117));
    defparam \transmit_module.i1609_4_lut_LC_14_19_0 .C_ON=1'b0;
    defparam \transmit_module.i1609_4_lut_LC_14_19_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1609_4_lut_LC_14_19_0 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \transmit_module.i1609_4_lut_LC_14_19_0  (
            .in0(N__19093),
            .in1(N__12496),
            .in2(N__21205),
            .in3(N__12481),
            .lcout(n18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i1_3_lut_LC_14_19_4 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i1_3_lut_LC_14_19_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i1_3_lut_LC_14_19_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_12_i1_3_lut_LC_14_19_4  (
            .in0(N__17908),
            .in1(N__12244),
            .in2(_gnd_net_),
            .in3(N__13455),
            .lcout(\transmit_module.n116 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i6_LC_14_21_5 .C_ON=1'b0;
    defparam \line_buffer.dout_i6_LC_14_21_5 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i6_LC_14_21_5 .LUT_INIT=16'b1111110000001010;
    LogicCell40 \line_buffer.dout_i6_LC_14_21_5  (
            .in0(N__12088),
            .in1(N__15679),
            .in2(N__21694),
            .in3(N__12238),
            .lcout(TX_DATA_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22747),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.VGA_R__i7_LC_14_23_7 .C_ON=1'b0;
    defparam \transmit_module.VGA_R__i7_LC_14_23_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.VGA_R__i7_LC_14_23_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.VGA_R__i7_LC_14_23_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12232),
            .lcout(n1792),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22557),
            .ce(),
            .sr(N__22319));
    defparam \transmit_module.VGA_R__i1_LC_14_24_4 .C_ON=1'b0;
    defparam \transmit_module.VGA_R__i1_LC_14_24_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.VGA_R__i1_LC_14_24_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.VGA_R__i1_LC_14_24_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13807),
            .lcout(n1798),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22650),
            .ce(),
            .sr(N__22321));
    defparam \line_buffer.i2353_3_lut_LC_14_25_4 .C_ON=1'b0;
    defparam \line_buffer.i2353_3_lut_LC_14_25_4 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2353_3_lut_LC_14_25_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \line_buffer.i2353_3_lut_LC_14_25_4  (
            .in0(N__12121),
            .in1(N__12103),
            .in2(_gnd_net_),
            .in3(N__23668),
            .lcout(\line_buffer.n3679 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1595_4_lut_LC_14_27_0 .C_ON=1'b0;
    defparam \transmit_module.i1595_4_lut_LC_14_27_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1595_4_lut_LC_14_27_0 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \transmit_module.i1595_4_lut_LC_14_27_0  (
            .in0(N__19109),
            .in1(N__12079),
            .in2(N__21280),
            .in3(N__12052),
            .lcout(n28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1605_4_lut_LC_14_28_2 .C_ON=1'b0;
    defparam \transmit_module.i1605_4_lut_LC_14_28_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1605_4_lut_LC_14_28_2 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \transmit_module.i1605_4_lut_LC_14_28_2  (
            .in0(N__19113),
            .in1(N__13057),
            .in2(N__21281),
            .in3(N__13033),
            .lcout(n22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1606_4_lut_LC_14_31_7 .C_ON=1'b0;
    defparam \transmit_module.i1606_4_lut_LC_14_31_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1606_4_lut_LC_14_31_7 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \transmit_module.i1606_4_lut_LC_14_31_7  (
            .in0(N__19114),
            .in1(N__12805),
            .in2(N__21282),
            .in3(N__12781),
            .lcout(n21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.PULSE_1HZ_49_LC_15_4_6 .C_ON=1'b0;
    defparam \receive_module.rx_counter.PULSE_1HZ_49_LC_15_4_6 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.PULSE_1HZ_49_LC_15_4_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \receive_module.rx_counter.PULSE_1HZ_49_LC_15_4_6  (
            .in0(_gnd_net_),
            .in1(N__12543),
            .in2(_gnd_net_),
            .in3(N__12523),
            .lcout(LED_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20128),
            .ce(N__16266),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i1_2_lut_LC_15_5_0 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i1_2_lut_LC_15_5_0 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i1_2_lut_LC_15_5_0 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \receive_module.rx_counter.i1_2_lut_LC_15_5_0  (
            .in0(_gnd_net_),
            .in1(N__16296),
            .in2(_gnd_net_),
            .in3(N__16326),
            .lcout(\receive_module.rx_counter.n7_adj_609 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i2302_2_lut_LC_15_5_1 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i2302_2_lut_LC_15_5_1 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i2302_2_lut_LC_15_5_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \receive_module.rx_counter.i2302_2_lut_LC_15_5_1  (
            .in0(_gnd_net_),
            .in1(N__16278),
            .in2(_gnd_net_),
            .in3(N__16341),
            .lcout(),
            .ltout(\receive_module.rx_counter.n3628_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i5_4_lut_LC_15_5_2 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i5_4_lut_LC_15_5_2 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i5_4_lut_LC_15_5_2 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \receive_module.rx_counter.i5_4_lut_LC_15_5_2  (
            .in0(N__16356),
            .in1(N__16311),
            .in2(N__12532),
            .in3(N__12529),
            .lcout(\receive_module.rx_counter.n11 ),
            .ltout(\receive_module.rx_counter.n11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i1286_2_lut_3_lut_LC_15_5_3 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i1286_2_lut_3_lut_LC_15_5_3 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i1286_2_lut_3_lut_LC_15_5_3 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \receive_module.rx_counter.i1286_2_lut_3_lut_LC_15_5_3  (
            .in0(N__20462),
            .in1(_gnd_net_),
            .in2(N__12517),
            .in3(N__12513),
            .lcout(\receive_module.rx_counter.n2517 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.old_VS_52_LC_15_5_4 .C_ON=1'b0;
    defparam \receive_module.rx_counter.old_VS_52_LC_15_5_4 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.old_VS_52_LC_15_5_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \receive_module.rx_counter.old_VS_52_LC_15_5_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20464),
            .lcout(\receive_module.rx_counter.old_VS ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20130),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i129_2_lut_rep_25_LC_15_5_6 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i129_2_lut_rep_25_LC_15_5_6 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i129_2_lut_rep_25_LC_15_5_6 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \receive_module.rx_counter.i129_2_lut_rep_25_LC_15_5_6  (
            .in0(N__12514),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20463),
            .lcout(\receive_module.rx_counter.n3792 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.O_VS_I_0_1_lut_rep_26_LC_15_7_1 .C_ON=1'b0;
    defparam \receive_module.rx_counter.O_VS_I_0_1_lut_rep_26_LC_15_7_1 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.O_VS_I_0_1_lut_rep_26_LC_15_7_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \receive_module.rx_counter.O_VS_I_0_1_lut_rep_26_LC_15_7_1  (
            .in0(N__20465),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\receive_module.n3793 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2315_3_lut_LC_15_10_1 .C_ON=1'b0;
    defparam \line_buffer.i2315_3_lut_LC_15_10_1 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2315_3_lut_LC_15_10_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \line_buffer.i2315_3_lut_LC_15_10_1  (
            .in0(N__13198),
            .in1(N__13183),
            .in2(_gnd_net_),
            .in3(N__23659),
            .lcout(\line_buffer.n3641 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i1_4_lut_LC_15_10_2 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i1_4_lut_LC_15_10_2 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i1_4_lut_LC_15_10_2 .LUT_INIT=16'b1010100010001000;
    LogicCell40 \receive_module.rx_counter.i1_4_lut_LC_15_10_2  (
            .in0(N__13165),
            .in1(N__13140),
            .in2(N__13129),
            .in3(N__13102),
            .lcout(\receive_module.rx_counter.n4_adj_606 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i248_3_lut_3_lut_3_lut_LC_15_10_3 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i248_3_lut_3_lut_3_lut_LC_15_10_3 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i248_3_lut_3_lut_3_lut_LC_15_10_3 .LUT_INIT=16'b0111011101010101;
    LogicCell40 \receive_module.rx_counter.i248_3_lut_3_lut_3_lut_LC_15_10_3  (
            .in0(N__20483),
            .in1(N__18651),
            .in2(_gnd_net_),
            .in3(N__13075),
            .lcout(\receive_module.rx_counter.n2045 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.old_HS_51_LC_15_10_4 .C_ON=1'b0;
    defparam \receive_module.rx_counter.old_HS_51_LC_15_10_4 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.old_HS_51_LC_15_10_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \receive_module.rx_counter.old_HS_51_LC_15_10_4  (
            .in0(N__18652),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\receive_module.rx_counter.old_HS ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20137),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_2_lut_LC_15_11_0 .C_ON=1'b1;
    defparam \receive_module.add_12_2_lut_LC_15_11_0 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_2_lut_LC_15_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_2_lut_LC_15_11_0  (
            .in0(_gnd_net_),
            .in1(N__16010),
            .in2(_gnd_net_),
            .in3(N__13069),
            .lcout(\receive_module.n136 ),
            .ltout(),
            .carryin(bfn_15_11_0_),
            .carryout(\receive_module.n3245 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_3_lut_LC_15_11_1 .C_ON=1'b1;
    defparam \receive_module.add_12_3_lut_LC_15_11_1 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_3_lut_LC_15_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_3_lut_LC_15_11_1  (
            .in0(_gnd_net_),
            .in1(N__15758),
            .in2(_gnd_net_),
            .in3(N__13066),
            .lcout(\receive_module.n135 ),
            .ltout(),
            .carryin(\receive_module.n3245 ),
            .carryout(\receive_module.n3246 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_4_lut_LC_15_11_2 .C_ON=1'b1;
    defparam \receive_module.add_12_4_lut_LC_15_11_2 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_4_lut_LC_15_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_4_lut_LC_15_11_2  (
            .in0(_gnd_net_),
            .in1(N__13589),
            .in2(_gnd_net_),
            .in3(N__13063),
            .lcout(\receive_module.n134 ),
            .ltout(),
            .carryin(\receive_module.n3246 ),
            .carryout(\receive_module.n3247 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_5_lut_LC_15_11_3 .C_ON=1'b1;
    defparam \receive_module.add_12_5_lut_LC_15_11_3 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_5_lut_LC_15_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_5_lut_LC_15_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20240),
            .in3(N__13060),
            .lcout(\receive_module.n133 ),
            .ltout(),
            .carryin(\receive_module.n3247 ),
            .carryout(\receive_module.n3248 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_6_lut_LC_15_11_4 .C_ON=1'b1;
    defparam \receive_module.add_12_6_lut_LC_15_11_4 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_6_lut_LC_15_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_6_lut_LC_15_11_4  (
            .in0(_gnd_net_),
            .in1(N__15218),
            .in2(_gnd_net_),
            .in3(N__13225),
            .lcout(\receive_module.n132 ),
            .ltout(),
            .carryin(\receive_module.n3248 ),
            .carryout(\receive_module.n3249 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_7_lut_LC_15_11_5 .C_ON=1'b1;
    defparam \receive_module.add_12_7_lut_LC_15_11_5 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_7_lut_LC_15_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_7_lut_LC_15_11_5  (
            .in0(_gnd_net_),
            .in1(N__14990),
            .in2(_gnd_net_),
            .in3(N__13222),
            .lcout(\receive_module.n131 ),
            .ltout(),
            .carryin(\receive_module.n3249 ),
            .carryout(\receive_module.n3250 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_8_lut_LC_15_11_6 .C_ON=1'b1;
    defparam \receive_module.add_12_8_lut_LC_15_11_6 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_8_lut_LC_15_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_8_lut_LC_15_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14714),
            .in3(N__13219),
            .lcout(\receive_module.n130 ),
            .ltout(),
            .carryin(\receive_module.n3250 ),
            .carryout(\receive_module.n3251 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_9_lut_LC_15_11_7 .C_ON=1'b1;
    defparam \receive_module.add_12_9_lut_LC_15_11_7 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_9_lut_LC_15_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_9_lut_LC_15_11_7  (
            .in0(_gnd_net_),
            .in1(N__14462),
            .in2(_gnd_net_),
            .in3(N__13216),
            .lcout(\receive_module.n129 ),
            .ltout(),
            .carryin(\receive_module.n3251 ),
            .carryout(\receive_module.n3252 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_10_lut_LC_15_12_0 .C_ON=1'b1;
    defparam \receive_module.add_12_10_lut_LC_15_12_0 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_10_lut_LC_15_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_10_lut_LC_15_12_0  (
            .in0(_gnd_net_),
            .in1(N__14210),
            .in2(_gnd_net_),
            .in3(N__13213),
            .lcout(\receive_module.n128 ),
            .ltout(),
            .carryin(bfn_15_12_0_),
            .carryout(\receive_module.n3253 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_11_lut_LC_15_12_1 .C_ON=1'b1;
    defparam \receive_module.add_12_11_lut_LC_15_12_1 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_11_lut_LC_15_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_11_lut_LC_15_12_1  (
            .in0(_gnd_net_),
            .in1(N__13976),
            .in2(_gnd_net_),
            .in3(N__13210),
            .lcout(\receive_module.n127 ),
            .ltout(),
            .carryin(\receive_module.n3253 ),
            .carryout(\receive_module.n3254 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_12_lut_LC_15_12_2 .C_ON=1'b1;
    defparam \receive_module.add_12_12_lut_LC_15_12_2 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_12_lut_LC_15_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_12_lut_LC_15_12_2  (
            .in0(_gnd_net_),
            .in1(N__15479),
            .in2(_gnd_net_),
            .in3(N__13207),
            .lcout(\receive_module.n126 ),
            .ltout(),
            .carryin(\receive_module.n3254 ),
            .carryout(\receive_module.n3255 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.BRAM_ADDR__i11_LC_15_12_3 .C_ON=1'b1;
    defparam \receive_module.BRAM_ADDR__i11_LC_15_12_3 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i11_LC_15_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.BRAM_ADDR__i11_LC_15_12_3  (
            .in0(_gnd_net_),
            .in1(N__16685),
            .in2(_gnd_net_),
            .in3(N__13204),
            .lcout(RX_ADDR_11),
            .ltout(),
            .carryin(\receive_module.n3255 ),
            .carryout(\receive_module.n3256 ),
            .clk(N__20143),
            .ce(N__17053),
            .sr(N__21946));
    defparam \receive_module.BRAM_ADDR__i12_LC_15_12_4 .C_ON=1'b1;
    defparam \receive_module.BRAM_ADDR__i12_LC_15_12_4 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i12_LC_15_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.BRAM_ADDR__i12_LC_15_12_4  (
            .in0(_gnd_net_),
            .in1(N__16784),
            .in2(_gnd_net_),
            .in3(N__13201),
            .lcout(RX_ADDR_12),
            .ltout(),
            .carryin(\receive_module.n3256 ),
            .carryout(\receive_module.n3257 ),
            .clk(N__20143),
            .ce(N__17053),
            .sr(N__21946));
    defparam \receive_module.BRAM_ADDR__i13_LC_15_12_5 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i13_LC_15_12_5 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i13_LC_15_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.BRAM_ADDR__i13_LC_15_12_5  (
            .in0(_gnd_net_),
            .in1(N__16737),
            .in2(_gnd_net_),
            .in3(N__13459),
            .lcout(RX_ADDR_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20143),
            .ce(N__17053),
            .sr(N__21946));
    defparam \transmit_module.add_13_2_lut_LC_15_13_0 .C_ON=1'b1;
    defparam \transmit_module.add_13_2_lut_LC_15_13_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_2_lut_LC_15_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_2_lut_LC_15_13_0  (
            .in0(_gnd_net_),
            .in1(N__13439),
            .in2(N__13422),
            .in3(_gnd_net_),
            .lcout(\transmit_module.n132 ),
            .ltout(),
            .carryin(bfn_15_13_0_),
            .carryout(\transmit_module.n3258 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_3_lut_LC_15_13_1 .C_ON=1'b1;
    defparam \transmit_module.add_13_3_lut_LC_15_13_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_3_lut_LC_15_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_3_lut_LC_15_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13389),
            .in3(N__13351),
            .lcout(\transmit_module.n131 ),
            .ltout(),
            .carryin(\transmit_module.n3258 ),
            .carryout(\transmit_module.n3259 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_4_lut_LC_15_13_2 .C_ON=1'b1;
    defparam \transmit_module.add_13_4_lut_LC_15_13_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_4_lut_LC_15_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_4_lut_LC_15_13_2  (
            .in0(_gnd_net_),
            .in1(N__17955),
            .in2(_gnd_net_),
            .in3(N__13348),
            .lcout(\transmit_module.n130 ),
            .ltout(),
            .carryin(\transmit_module.n3259 ),
            .carryout(\transmit_module.n3260 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_5_lut_LC_15_13_3 .C_ON=1'b1;
    defparam \transmit_module.add_13_5_lut_LC_15_13_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_5_lut_LC_15_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_5_lut_LC_15_13_3  (
            .in0(_gnd_net_),
            .in1(N__17796),
            .in2(_gnd_net_),
            .in3(N__13345),
            .lcout(\transmit_module.n129 ),
            .ltout(),
            .carryin(\transmit_module.n3260 ),
            .carryout(\transmit_module.n3261 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_6_lut_LC_15_13_4 .C_ON=1'b1;
    defparam \transmit_module.add_13_6_lut_LC_15_13_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_6_lut_LC_15_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_6_lut_LC_15_13_4  (
            .in0(_gnd_net_),
            .in1(N__13336),
            .in2(_gnd_net_),
            .in3(N__13309),
            .lcout(\transmit_module.n128 ),
            .ltout(),
            .carryin(\transmit_module.n3261 ),
            .carryout(\transmit_module.n3262 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_7_lut_LC_15_13_5 .C_ON=1'b1;
    defparam \transmit_module.add_13_7_lut_LC_15_13_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_7_lut_LC_15_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_7_lut_LC_15_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13304),
            .in3(N__13270),
            .lcout(\transmit_module.n127 ),
            .ltout(),
            .carryin(\transmit_module.n3262 ),
            .carryout(\transmit_module.n3263 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_8_lut_LC_15_13_6 .C_ON=1'b1;
    defparam \transmit_module.add_13_8_lut_LC_15_13_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_8_lut_LC_15_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_8_lut_LC_15_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13265),
            .in3(N__13228),
            .lcout(\transmit_module.n126 ),
            .ltout(),
            .carryin(\transmit_module.n3263 ),
            .carryout(\transmit_module.n3264 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_9_lut_LC_15_13_7 .C_ON=1'b1;
    defparam \transmit_module.add_13_9_lut_LC_15_13_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_9_lut_LC_15_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_9_lut_LC_15_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13544),
            .in3(N__13507),
            .lcout(\transmit_module.n125 ),
            .ltout(),
            .carryin(\transmit_module.n3264 ),
            .carryout(\transmit_module.n3265 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_10_lut_LC_15_14_0 .C_ON=1'b1;
    defparam \transmit_module.add_13_10_lut_LC_15_14_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_10_lut_LC_15_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_10_lut_LC_15_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17353),
            .in3(N__13504),
            .lcout(\transmit_module.n124 ),
            .ltout(),
            .carryin(bfn_15_14_0_),
            .carryout(\transmit_module.n3266 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_11_lut_LC_15_14_1 .C_ON=1'b1;
    defparam \transmit_module.add_13_11_lut_LC_15_14_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_11_lut_LC_15_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_11_lut_LC_15_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17332),
            .in3(N__13501),
            .lcout(\transmit_module.n123 ),
            .ltout(),
            .carryin(\transmit_module.n3266 ),
            .carryout(\transmit_module.n3267 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_12_lut_LC_15_14_2 .C_ON=1'b1;
    defparam \transmit_module.add_13_12_lut_LC_15_14_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_12_lut_LC_15_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_12_lut_LC_15_14_2  (
            .in0(_gnd_net_),
            .in1(N__13495),
            .in2(_gnd_net_),
            .in3(N__13471),
            .lcout(\transmit_module.n122 ),
            .ltout(),
            .carryin(\transmit_module.n3267 ),
            .carryout(\transmit_module.n3268 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_13_lut_LC_15_14_3 .C_ON=1'b1;
    defparam \transmit_module.add_13_13_lut_LC_15_14_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_13_lut_LC_15_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_13_lut_LC_15_14_3  (
            .in0(_gnd_net_),
            .in1(N__23629),
            .in2(_gnd_net_),
            .in3(N__13468),
            .lcout(\transmit_module.n121 ),
            .ltout(),
            .carryin(\transmit_module.n3268 ),
            .carryout(\transmit_module.n3269 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_14_lut_LC_15_14_4 .C_ON=1'b1;
    defparam \transmit_module.add_13_14_lut_LC_15_14_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_14_lut_LC_15_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_14_lut_LC_15_14_4  (
            .in0(_gnd_net_),
            .in1(N__22173),
            .in2(_gnd_net_),
            .in3(N__13465),
            .lcout(\transmit_module.n120 ),
            .ltout(),
            .carryin(\transmit_module.n3269 ),
            .carryout(\transmit_module.n3270 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_15_lut_LC_15_14_5 .C_ON=1'b0;
    defparam \transmit_module.add_13_15_lut_LC_15_14_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_15_lut_LC_15_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_15_lut_LC_15_14_5  (
            .in0(_gnd_net_),
            .in1(N__21645),
            .in2(_gnd_net_),
            .in3(N__13462),
            .lcout(\transmit_module.n119 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.ADDR_Y_COMPONENT__i9_LC_15_14_6 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i9_LC_15_14_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i9_LC_15_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i9_LC_15_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17329),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22982),
            .ce(N__17766),
            .sr(N__21053));
    defparam \transmit_module.ADDR_Y_COMPONENT__i8_LC_15_14_7 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i8_LC_15_14_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i8_LC_15_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i8_LC_15_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17350),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22982),
            .ce(N__17766),
            .sr(N__21053));
    defparam \transmit_module.mux_12_i10_3_lut_LC_15_15_4 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i10_3_lut_LC_15_15_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i10_3_lut_LC_15_15_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_12_i10_3_lut_LC_15_15_4  (
            .in0(N__17884),
            .in1(N__13900),
            .in2(_gnd_net_),
            .in3(N__17331),
            .lcout(\transmit_module.n107 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1613_4_lut_LC_15_15_5 .C_ON=1'b0;
    defparam \transmit_module.i1613_4_lut_LC_15_15_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1613_4_lut_LC_15_15_5 .LUT_INIT=16'b1111011111110100;
    LogicCell40 \transmit_module.i1613_4_lut_LC_15_15_5  (
            .in0(N__17907),
            .in1(N__19024),
            .in2(N__21138),
            .in3(N__18307),
            .lcout(\transmit_module.n2039 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i12_LC_15_16_1 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i12_LC_15_16_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i12_LC_15_16_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \transmit_module.BRAM_ADDR__i12_LC_15_16_1  (
            .in0(N__13894),
            .in1(N__19097),
            .in2(_gnd_net_),
            .in3(N__13885),
            .lcout(TX_ADDR_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22854),
            .ce(N__13846),
            .sr(N__21049));
    defparam \transmit_module.BRAM_ADDR__i13_LC_15_16_5 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i13_LC_15_16_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i13_LC_15_16_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \transmit_module.BRAM_ADDR__i13_LC_15_16_5  (
            .in0(N__17581),
            .in1(N__19098),
            .in2(_gnd_net_),
            .in3(N__13876),
            .lcout(TX_ADDR_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22854),
            .ce(N__13846),
            .sr(N__21049));
    defparam \transmit_module.BRAM_ADDR__rep_1_i0_LC_15_17_6 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__rep_1_i0_LC_15_17_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__rep_1_i0_LC_15_17_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \transmit_module.BRAM_ADDR__rep_1_i0_LC_15_17_6  (
            .in0(N__13867),
            .in1(N__19064),
            .in2(_gnd_net_),
            .in3(N__13855),
            .lcout(TX_ADDR_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22872),
            .ce(N__13842),
            .sr(N__21235));
    defparam \transmit_module.mux_14_i3_3_lut_LC_15_18_2 .C_ON=1'b0;
    defparam \transmit_module.mux_14_i3_3_lut_LC_15_18_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_14_i3_3_lut_LC_15_18_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \transmit_module.mux_14_i3_3_lut_LC_15_18_2  (
            .in0(N__17979),
            .in1(N__18315),
            .in2(_gnd_net_),
            .in3(N__13822),
            .lcout(\transmit_module.n145 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i0_LC_15_18_4 .C_ON=1'b0;
    defparam \line_buffer.dout_i0_LC_15_18_4 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i0_LC_15_18_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \line_buffer.dout_i0_LC_15_18_4  (
            .in0(N__21652),
            .in1(N__13813),
            .in2(_gnd_net_),
            .in3(N__17521),
            .lcout(TX_DATA_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22833),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.BRAM_ADDR__i2_LC_15_19_7 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i2_LC_15_19_7 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i2_LC_15_19_7 .LUT_INIT=16'b1101110010001100;
    LogicCell40 \receive_module.BRAM_ADDR__i2_LC_15_19_7  (
            .in0(N__20672),
            .in1(N__13795),
            .in2(N__20503),
            .in3(N__13570),
            .lcout(RX_ADDR_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20152),
            .ce(),
            .sr(N__21979));
    defparam \transmit_module.video_signal_controller.i1120_1_lut_LC_15_20_3 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1120_1_lut_LC_15_20_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1120_1_lut_LC_15_20_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \transmit_module.video_signal_controller.i1120_1_lut_LC_15_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18316),
            .lcout(\transmit_module.n2354 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2354_3_lut_LC_15_21_4 .C_ON=1'b0;
    defparam \line_buffer.i2354_3_lut_LC_15_21_4 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2354_3_lut_LC_15_21_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \line_buffer.i2354_3_lut_LC_15_21_4  (
            .in0(N__15715),
            .in1(N__15700),
            .in2(_gnd_net_),
            .in3(N__23664),
            .lcout(\line_buffer.n3680 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.BRAM_ADDR__i10_LC_15_23_6 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i10_LC_15_23_6 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i10_LC_15_23_6 .LUT_INIT=16'b1110111101000000;
    LogicCell40 \receive_module.BRAM_ADDR__i10_LC_15_23_6  (
            .in0(N__20678),
            .in1(N__15442),
            .in2(N__20536),
            .in3(N__15673),
            .lcout(RX_ADDR_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20158),
            .ce(),
            .sr(N__21990));
    defparam \receive_module.BRAM_ADDR__i4_LC_15_31_1 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i4_LC_15_31_1 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i4_LC_15_31_1 .LUT_INIT=16'b1101110010001100;
    LogicCell40 \receive_module.BRAM_ADDR__i4_LC_15_31_1  (
            .in0(N__20693),
            .in1(N__15415),
            .in2(N__20567),
            .in3(N__15202),
            .lcout(RX_ADDR_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20170),
            .ce(),
            .sr(N__21997));
    defparam \receive_module.BRAM_ADDR__i5_LC_15_31_2 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i5_LC_15_31_2 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i5_LC_15_31_2 .LUT_INIT=16'b1010101011100010;
    LogicCell40 \receive_module.BRAM_ADDR__i5_LC_15_31_2  (
            .in0(N__15178),
            .in1(N__20557),
            .in2(N__14956),
            .in3(N__20696),
            .lcout(RX_ADDR_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20170),
            .ce(),
            .sr(N__21997));
    defparam \receive_module.BRAM_ADDR__i6_LC_15_31_3 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i6_LC_15_31_3 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i6_LC_15_31_3 .LUT_INIT=16'b1110111101000000;
    LogicCell40 \receive_module.BRAM_ADDR__i6_LC_15_31_3  (
            .in0(N__20694),
            .in1(N__14686),
            .in2(N__20568),
            .in3(N__14914),
            .lcout(RX_ADDR_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20170),
            .ce(),
            .sr(N__21997));
    defparam \receive_module.BRAM_ADDR__i7_LC_15_31_4 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i7_LC_15_31_4 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i7_LC_15_31_4 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \receive_module.BRAM_ADDR__i7_LC_15_31_4  (
            .in0(N__20564),
            .in1(N__20697),
            .in2(N__14446),
            .in3(N__14662),
            .lcout(RX_ADDR_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20170),
            .ce(),
            .sr(N__21997));
    defparam \receive_module.BRAM_ADDR__i8_LC_15_31_5 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i8_LC_15_31_5 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i8_LC_15_31_5 .LUT_INIT=16'b1110111101000000;
    LogicCell40 \receive_module.BRAM_ADDR__i8_LC_15_31_5  (
            .in0(N__20695),
            .in1(N__14182),
            .in2(N__20569),
            .in3(N__14407),
            .lcout(RX_ADDR_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20170),
            .ce(),
            .sr(N__21997));
    defparam \receive_module.BRAM_ADDR__i9_LC_15_31_6 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i9_LC_15_31_6 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i9_LC_15_31_6 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \receive_module.BRAM_ADDR__i9_LC_15_31_6  (
            .in0(N__20565),
            .in1(N__20698),
            .in2(N__13942),
            .in3(N__14158),
            .lcout(RX_ADDR_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20170),
            .ce(),
            .sr(N__21997));
    defparam \receive_module.rx_counter.FRAME_COUNTER_243__i0_LC_16_5_0 .C_ON=1'b1;
    defparam \receive_module.rx_counter.FRAME_COUNTER_243__i0_LC_16_5_0 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.FRAME_COUNTER_243__i0_LC_16_5_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.FRAME_COUNTER_243__i0_LC_16_5_0  (
            .in0(_gnd_net_),
            .in1(N__16357),
            .in2(_gnd_net_),
            .in3(N__16345),
            .lcout(\receive_module.rx_counter.FRAME_COUNTER_0 ),
            .ltout(),
            .carryin(bfn_16_5_0_),
            .carryout(\receive_module.rx_counter.n3310 ),
            .clk(N__20129),
            .ce(N__16267),
            .sr(N__16243));
    defparam \receive_module.rx_counter.FRAME_COUNTER_243__i1_LC_16_5_1 .C_ON=1'b1;
    defparam \receive_module.rx_counter.FRAME_COUNTER_243__i1_LC_16_5_1 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.FRAME_COUNTER_243__i1_LC_16_5_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.FRAME_COUNTER_243__i1_LC_16_5_1  (
            .in0(_gnd_net_),
            .in1(N__16342),
            .in2(_gnd_net_),
            .in3(N__16330),
            .lcout(\receive_module.rx_counter.FRAME_COUNTER_1 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3310 ),
            .carryout(\receive_module.rx_counter.n3311 ),
            .clk(N__20129),
            .ce(N__16267),
            .sr(N__16243));
    defparam \receive_module.rx_counter.FRAME_COUNTER_243__i2_LC_16_5_2 .C_ON=1'b1;
    defparam \receive_module.rx_counter.FRAME_COUNTER_243__i2_LC_16_5_2 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.FRAME_COUNTER_243__i2_LC_16_5_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.FRAME_COUNTER_243__i2_LC_16_5_2  (
            .in0(_gnd_net_),
            .in1(N__16327),
            .in2(_gnd_net_),
            .in3(N__16315),
            .lcout(\receive_module.rx_counter.FRAME_COUNTER_2 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3311 ),
            .carryout(\receive_module.rx_counter.n3312 ),
            .clk(N__20129),
            .ce(N__16267),
            .sr(N__16243));
    defparam \receive_module.rx_counter.FRAME_COUNTER_243__i3_LC_16_5_3 .C_ON=1'b1;
    defparam \receive_module.rx_counter.FRAME_COUNTER_243__i3_LC_16_5_3 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.FRAME_COUNTER_243__i3_LC_16_5_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.FRAME_COUNTER_243__i3_LC_16_5_3  (
            .in0(_gnd_net_),
            .in1(N__16312),
            .in2(_gnd_net_),
            .in3(N__16300),
            .lcout(\receive_module.rx_counter.FRAME_COUNTER_3 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3312 ),
            .carryout(\receive_module.rx_counter.n3313 ),
            .clk(N__20129),
            .ce(N__16267),
            .sr(N__16243));
    defparam \receive_module.rx_counter.FRAME_COUNTER_243__i4_LC_16_5_4 .C_ON=1'b1;
    defparam \receive_module.rx_counter.FRAME_COUNTER_243__i4_LC_16_5_4 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.FRAME_COUNTER_243__i4_LC_16_5_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.FRAME_COUNTER_243__i4_LC_16_5_4  (
            .in0(_gnd_net_),
            .in1(N__16297),
            .in2(_gnd_net_),
            .in3(N__16285),
            .lcout(\receive_module.rx_counter.FRAME_COUNTER_4 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3313 ),
            .carryout(\receive_module.rx_counter.n3314 ),
            .clk(N__20129),
            .ce(N__16267),
            .sr(N__16243));
    defparam \receive_module.rx_counter.FRAME_COUNTER_243__i5_LC_16_5_5 .C_ON=1'b0;
    defparam \receive_module.rx_counter.FRAME_COUNTER_243__i5_LC_16_5_5 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.FRAME_COUNTER_243__i5_LC_16_5_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.FRAME_COUNTER_243__i5_LC_16_5_5  (
            .in0(_gnd_net_),
            .in1(N__16279),
            .in2(_gnd_net_),
            .in3(N__16282),
            .lcout(\receive_module.rx_counter.FRAME_COUNTER_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20129),
            .ce(N__16267),
            .sr(N__16243));
    defparam \receive_module.BRAM_ADDR__i0_LC_16_7_0 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i0_LC_16_7_0 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i0_LC_16_7_0 .LUT_INIT=16'b1101110010001100;
    LogicCell40 \receive_module.BRAM_ADDR__i0_LC_16_7_0  (
            .in0(N__20673),
            .in1(N__16231),
            .in2(N__20535),
            .in3(N__15994),
            .lcout(RX_ADDR_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20131),
            .ce(),
            .sr(N__21933));
    defparam \receive_module.BRAM_ADDR__i1_LC_16_7_1 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i1_LC_16_7_1 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i1_LC_16_7_1 .LUT_INIT=16'b1111000010111000;
    LogicCell40 \receive_module.BRAM_ADDR__i1_LC_16_7_1  (
            .in0(N__15751),
            .in1(N__20521),
            .in2(N__15973),
            .in3(N__20674),
            .lcout(RX_ADDR_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20131),
            .ce(),
            .sr(N__21933));
    defparam \line_buffer.i2308_3_lut_LC_16_8_6 .C_ON=1'b0;
    defparam \line_buffer.i2308_3_lut_LC_16_8_6 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2308_3_lut_LC_16_8_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \line_buffer.i2308_3_lut_LC_16_8_6  (
            .in0(N__23667),
            .in1(N__16573),
            .in2(_gnd_net_),
            .in3(N__16555),
            .lcout(\line_buffer.n3634 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2350_3_lut_LC_16_9_5 .C_ON=1'b0;
    defparam \line_buffer.i2350_3_lut_LC_16_9_5 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2350_3_lut_LC_16_9_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \line_buffer.i2350_3_lut_LC_16_9_5  (
            .in0(N__23655),
            .in1(N__16543),
            .in2(_gnd_net_),
            .in3(N__16525),
            .lcout(\line_buffer.n3676 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i1_2_lut_adj_22_LC_16_10_2 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i1_2_lut_adj_22_LC_16_10_2 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i1_2_lut_adj_22_LC_16_10_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \receive_module.rx_counter.i1_2_lut_adj_22_LC_16_10_2  (
            .in0(_gnd_net_),
            .in1(N__18593),
            .in2(_gnd_net_),
            .in3(N__19337),
            .lcout(),
            .ltout(\receive_module.rx_counter.n4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i2_4_lut_LC_16_10_3 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i2_4_lut_LC_16_10_3 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i2_4_lut_LC_16_10_3 .LUT_INIT=16'b1100100000000000;
    LogicCell40 \receive_module.rx_counter.i2_4_lut_LC_16_10_3  (
            .in0(N__19320),
            .in1(N__19301),
            .in2(N__16510),
            .in3(N__19283),
            .lcout(\receive_module.rx_counter.n3581 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i2_2_lut_adj_19_LC_16_10_4 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i2_2_lut_adj_19_LC_16_10_4 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i2_2_lut_adj_19_LC_16_10_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \receive_module.rx_counter.i2_2_lut_adj_19_LC_16_10_4  (
            .in0(_gnd_net_),
            .in1(N__19319),
            .in2(_gnd_net_),
            .in3(N__19338),
            .lcout(),
            .ltout(\receive_module.rx_counter.n6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i2208_4_lut_LC_16_10_5 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i2208_4_lut_LC_16_10_5 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i2208_4_lut_LC_16_10_5 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \receive_module.rx_counter.i2208_4_lut_LC_16_10_5  (
            .in0(N__18594),
            .in1(N__19302),
            .in2(N__16507),
            .in3(N__19284),
            .lcout(\receive_module.rx_counter.n3534 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i59_4_lut_LC_16_11_1 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i59_4_lut_LC_16_11_1 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i59_4_lut_LC_16_11_1 .LUT_INIT=16'b1111000110100001;
    LogicCell40 \receive_module.rx_counter.i59_4_lut_LC_16_11_1  (
            .in0(N__19266),
            .in1(N__16504),
            .in2(N__19249),
            .in3(N__16498),
            .lcout(\receive_module.rx_counter.n55_adj_607 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_12_LC_16_11_3 .C_ON=1'b0;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_12_LC_16_11_3 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_12_LC_16_11_3 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \line_buffer.i1_2_lut_3_lut_4_lut_adj_12_LC_16_11_3  (
            .in0(N__16782),
            .in1(N__20635),
            .in2(N__16686),
            .in3(N__16735),
            .lcout(\line_buffer.n517 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_17_LC_16_11_4 .C_ON=1'b0;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_17_LC_16_11_4 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_17_LC_16_11_4 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \line_buffer.i1_2_lut_3_lut_4_lut_adj_17_LC_16_11_4  (
            .in0(N__16678),
            .in1(N__16781),
            .in2(N__16741),
            .in3(N__20634),
            .lcout(\line_buffer.n452 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_15_LC_16_11_5 .C_ON=1'b0;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_15_LC_16_11_5 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_15_LC_16_11_5 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \line_buffer.i1_2_lut_3_lut_4_lut_adj_15_LC_16_11_5  (
            .in0(N__16783),
            .in1(N__20636),
            .in2(N__16687),
            .in3(N__16736),
            .lcout(\line_buffer.n548 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.i245_2_lut_rep_28_LC_16_12_0 .C_ON=1'b0;
    defparam \receive_module.i245_2_lut_rep_28_LC_16_12_0 .SEQ_MODE=4'b0000;
    defparam \receive_module.i245_2_lut_rep_28_LC_16_12_0 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \receive_module.i245_2_lut_rep_28_LC_16_12_0  (
            .in0(N__20631),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20534),
            .lcout(\receive_module.n3795 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_14_LC_16_12_2 .C_ON=1'b0;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_14_LC_16_12_2 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_14_LC_16_12_2 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \line_buffer.i1_2_lut_3_lut_4_lut_adj_14_LC_16_12_2  (
            .in0(N__20629),
            .in1(N__16674),
            .in2(N__16785),
            .in3(N__16724),
            .lcout(\line_buffer.n451 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_16_LC_16_12_4 .C_ON=1'b0;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_16_LC_16_12_4 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_16_LC_16_12_4 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \line_buffer.i1_2_lut_3_lut_4_lut_adj_16_LC_16_12_4  (
            .in0(N__20630),
            .in1(N__16675),
            .in2(N__16786),
            .in3(N__16725),
            .lcout(\line_buffer.n549 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_13_LC_16_12_5 .C_ON=1'b0;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_13_LC_16_12_5 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_13_LC_16_12_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \line_buffer.i1_2_lut_3_lut_4_lut_adj_13_LC_16_12_5  (
            .in0(N__16673),
            .in1(N__16772),
            .in2(N__16738),
            .in3(N__20628),
            .lcout(\line_buffer.n516 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.O_VISIBLE_53_LC_16_12_7 .C_ON=1'b0;
    defparam \receive_module.rx_counter.O_VISIBLE_53_LC_16_12_7 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.O_VISIBLE_53_LC_16_12_7 .LUT_INIT=16'b0000000000101010;
    LogicCell40 \receive_module.rx_counter.O_VISIBLE_53_LC_16_12_7  (
            .in0(N__16891),
            .in1(N__16879),
            .in2(N__16870),
            .in3(N__16834),
            .lcout(RX_WE),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20139),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_11_LC_16_13_0 .C_ON=1'b0;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_11_LC_16_13_0 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_11_LC_16_13_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \line_buffer.i1_2_lut_3_lut_4_lut_adj_11_LC_16_13_0  (
            .in0(N__16677),
            .in1(N__16780),
            .in2(N__16740),
            .in3(N__20633),
            .lcout(\line_buffer.n581 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_LC_16_13_1 .C_ON=1'b0;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_LC_16_13_1 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_LC_16_13_1 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \line_buffer.i1_2_lut_3_lut_4_lut_LC_16_13_1  (
            .in0(N__16779),
            .in1(N__20632),
            .in2(N__16739),
            .in3(N__16676),
            .lcout(\line_buffer.n580 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i3_LC_16_13_3 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i3_LC_16_13_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i3_LC_16_13_3 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \transmit_module.BRAM_ADDR__i3_LC_16_13_3  (
            .in0(N__19068),
            .in1(N__17827),
            .in2(N__21268),
            .in3(N__18208),
            .lcout(\transmit_module.TX_ADDR_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22825),
            .ce(),
            .sr(_gnd_net_));
    defparam \sync_buffer.WIRE_OUT_8_LC_16_14_1 .C_ON=1'b0;
    defparam \sync_buffer.WIRE_OUT_8_LC_16_14_1 .SEQ_MODE=4'b1000;
    defparam \sync_buffer.WIRE_OUT_8_LC_16_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sync_buffer.WIRE_OUT_8_LC_16_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17374),
            .lcout(RX_TX_SYNC_BUFF),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVsync_buffer.WIRE_OUT_8C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \sync_buffer.BUFFER_i0_LC_16_14_5 .C_ON=1'b0;
    defparam \sync_buffer.BUFFER_i0_LC_16_14_5 .SEQ_MODE=4'b1000;
    defparam \sync_buffer.BUFFER_i0_LC_16_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sync_buffer.BUFFER_i0_LC_16_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17392),
            .lcout(\sync_buffer.BUFFER_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVsync_buffer.WIRE_OUT_8C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \sync_buffer.BUFFER_i1_LC_16_14_7 .C_ON=1'b0;
    defparam \sync_buffer.BUFFER_i1_LC_16_14_7 .SEQ_MODE=4'b1000;
    defparam \sync_buffer.BUFFER_i1_LC_16_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sync_buffer.BUFFER_i1_LC_16_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17380),
            .lcout(\sync_buffer.BUFFER_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVsync_buffer.WIRE_OUT_8C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_14_i9_3_lut_LC_16_15_1 .C_ON=1'b0;
    defparam \transmit_module.mux_14_i9_3_lut_LC_16_15_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_14_i9_3_lut_LC_16_15_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_14_i9_3_lut_LC_16_15_1  (
            .in0(N__18302),
            .in1(N__17351),
            .in2(_gnd_net_),
            .in3(N__17368),
            .lcout(\transmit_module.n139 ),
            .ltout(\transmit_module.n139_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i8_LC_16_15_2 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i8_LC_16_15_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i8_LC_16_15_2 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \transmit_module.BRAM_ADDR__i8_LC_16_15_2  (
            .in0(N__21055),
            .in1(N__19066),
            .in2(N__17362),
            .in3(N__18912),
            .lcout(\transmit_module.TX_ADDR_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22809),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i9_3_lut_LC_16_15_3 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i9_3_lut_LC_16_15_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i9_3_lut_LC_16_15_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_12_i9_3_lut_LC_16_15_3  (
            .in0(N__17928),
            .in1(N__17359),
            .in2(_gnd_net_),
            .in3(N__17352),
            .lcout(\transmit_module.n108 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i9_LC_16_15_4 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i9_LC_16_15_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i9_LC_16_15_4 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \transmit_module.BRAM_ADDR__i9_LC_16_15_4  (
            .in0(N__19067),
            .in1(N__17293),
            .in2(N__21166),
            .in3(N__17302),
            .lcout(\transmit_module.TX_ADDR_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22809),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_14_i10_3_lut_LC_16_15_5 .C_ON=1'b0;
    defparam \transmit_module.mux_14_i10_3_lut_LC_16_15_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_14_i10_3_lut_LC_16_15_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_14_i10_3_lut_LC_16_15_5  (
            .in0(N__18303),
            .in1(N__17330),
            .in2(_gnd_net_),
            .in3(N__17308),
            .lcout(\transmit_module.n138 ),
            .ltout(\transmit_module.n138_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1608_4_lut_LC_16_15_6 .C_ON=1'b0;
    defparam \transmit_module.i1608_4_lut_LC_16_15_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1608_4_lut_LC_16_15_6 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \transmit_module.i1608_4_lut_LC_16_15_6  (
            .in0(N__21054),
            .in1(N__19065),
            .in2(N__17296),
            .in3(N__17292),
            .lcout(n19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.ADDR_Y_COMPONENT__i13_LC_16_16_3 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i13_LC_16_16_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i13_LC_16_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i13_LC_16_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21644),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22853),
            .ce(N__17779),
            .sr(N__21266));
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_LC_16_17_0 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_LC_16_17_0 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_LC_16_17_0 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \line_buffer.TX_ADDR_12__bdd_4_lut_LC_16_17_0  (
            .in0(N__22124),
            .in1(N__19345),
            .in2(N__21675),
            .in3(N__17575),
            .lcout(\line_buffer.n3728 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n3746_bdd_4_lut_LC_16_17_2 .C_ON=1'b0;
    defparam \line_buffer.n3746_bdd_4_lut_LC_16_17_2 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3746_bdd_4_lut_LC_16_17_2 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \line_buffer.n3746_bdd_4_lut_LC_16_17_2  (
            .in0(N__17563),
            .in1(N__22123),
            .in2(N__17545),
            .in3(N__19414),
            .lcout(\line_buffer.n3749 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2348_3_lut_LC_16_17_3 .C_ON=1'b0;
    defparam \line_buffer.i2348_3_lut_LC_16_17_3 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2348_3_lut_LC_16_17_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \line_buffer.i2348_3_lut_LC_16_17_3  (
            .in0(N__17515),
            .in1(N__17497),
            .in2(_gnd_net_),
            .in3(N__23543),
            .lcout(\line_buffer.n3674 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_2392_LC_16_17_6 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_2392_LC_16_17_6 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_2392_LC_16_17_6 .LUT_INIT=16'b1011110010001100;
    LogicCell40 \line_buffer.TX_ADDR_12__bdd_4_lut_2392_LC_16_17_6  (
            .in0(N__19378),
            .in1(N__22122),
            .in2(N__21674),
            .in3(N__17479),
            .lcout(\line_buffer.n3716 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i2_LC_16_18_3 .C_ON=1'b0;
    defparam \line_buffer.dout_i2_LC_16_18_3 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i2_LC_16_18_3 .LUT_INIT=16'b1111110000001010;
    LogicCell40 \line_buffer.dout_i2_LC_16_18_3  (
            .in0(N__19123),
            .in1(N__17467),
            .in2(N__21682),
            .in3(N__17461),
            .lcout(TX_DATA_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22883),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2314_3_lut_LC_16_18_4 .C_ON=1'b0;
    defparam \line_buffer.i2314_3_lut_LC_16_18_4 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2314_3_lut_LC_16_18_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \line_buffer.i2314_3_lut_LC_16_18_4  (
            .in0(N__17455),
            .in1(N__17440),
            .in2(_gnd_net_),
            .in3(N__23544),
            .lcout(),
            .ltout(\line_buffer.n3640_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i4_LC_16_18_5 .C_ON=1'b0;
    defparam \line_buffer.dout_i4_LC_16_18_5 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i4_LC_16_18_5 .LUT_INIT=16'b1101110010011000;
    LogicCell40 \line_buffer.dout_i4_LC_16_18_5  (
            .in0(N__21661),
            .in1(N__17425),
            .in2(N__17419),
            .in3(N__17416),
            .lcout(TX_DATA_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22883),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i3_3_lut_LC_16_18_7 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i3_3_lut_LC_16_18_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i3_3_lut_LC_16_18_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_12_i3_3_lut_LC_16_18_7  (
            .in0(N__17929),
            .in1(N__17944),
            .in2(_gnd_net_),
            .in3(N__17972),
            .lcout(\transmit_module.n114 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1601_4_lut_LC_16_19_0 .C_ON=1'b0;
    defparam \transmit_module.i1601_4_lut_LC_16_19_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1601_4_lut_LC_16_19_0 .LUT_INIT=16'b0000101100001000;
    LogicCell40 \transmit_module.i1601_4_lut_LC_16_19_0  (
            .in0(N__18567),
            .in1(N__19059),
            .in2(N__21265),
            .in3(N__18549),
            .lcout(n26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_14_i4_3_lut_LC_16_19_2 .C_ON=1'b0;
    defparam \transmit_module.mux_14_i4_3_lut_LC_16_19_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_14_i4_3_lut_LC_16_19_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_14_i4_3_lut_LC_16_19_2  (
            .in0(N__18314),
            .in1(N__17808),
            .in2(_gnd_net_),
            .in3(N__18220),
            .lcout(\transmit_module.n144 ),
            .ltout(\transmit_module.n144_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1602_4_lut_LC_16_19_3 .C_ON=1'b0;
    defparam \transmit_module.i1602_4_lut_LC_16_19_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1602_4_lut_LC_16_19_3 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \transmit_module.i1602_4_lut_LC_16_19_3  (
            .in0(N__19060),
            .in1(N__21178),
            .in2(N__18196),
            .in3(N__17820),
            .lcout(n25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.ADDR_Y_COMPONENT__i2_LC_16_19_4 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i2_LC_16_19_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i2_LC_16_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i2_LC_16_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17980),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22694),
            .ce(N__17778),
            .sr(N__21283));
    defparam \transmit_module.mux_12_i4_3_lut_LC_16_19_5 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i4_3_lut_LC_16_19_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i4_3_lut_LC_16_19_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \transmit_module.mux_12_i4_3_lut_LC_16_19_5  (
            .in0(N__17807),
            .in1(N__17937),
            .in2(_gnd_net_),
            .in3(N__17785),
            .lcout(\transmit_module.n113 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.ADDR_Y_COMPONENT__i3_LC_16_19_6 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i3_LC_16_19_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i3_LC_16_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i3_LC_16_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17809),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22694),
            .ce(N__17778),
            .sr(N__21283));
    defparam \transmit_module.VGA_R__i5_LC_16_20_2 .C_ON=1'b0;
    defparam \transmit_module.VGA_R__i5_LC_16_20_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.VGA_R__i5_LC_16_20_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.VGA_R__i5_LC_16_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17707),
            .lcout(n1794),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22558),
            .ce(),
            .sr(N__22315));
    defparam \transmit_module.VGA_R__i3_LC_16_20_7 .C_ON=1'b0;
    defparam \transmit_module.VGA_R__i3_LC_16_20_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.VGA_R__i3_LC_16_20_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.VGA_R__i3_LC_16_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17638),
            .lcout(n1796),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22558),
            .ce(),
            .sr(N__22315));
    defparam \line_buffer.i2347_3_lut_LC_16_21_7 .C_ON=1'b0;
    defparam \line_buffer.i2347_3_lut_LC_16_21_7 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2347_3_lut_LC_16_21_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \line_buffer.i2347_3_lut_LC_16_21_7  (
            .in0(N__19156),
            .in1(N__19141),
            .in2(_gnd_net_),
            .in3(N__23665),
            .lcout(\line_buffer.n3673 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1607_4_lut_LC_16_23_1 .C_ON=1'b0;
    defparam \transmit_module.i1607_4_lut_LC_16_23_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1607_4_lut_LC_16_23_1 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \transmit_module.i1607_4_lut_LC_16_23_1  (
            .in0(N__19086),
            .in1(N__18916),
            .in2(N__21318),
            .in3(N__18898),
            .lcout(n20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_TVP_CLK_c_THRU_LUT4_0_LC_16_32_3.C_ON=1'b0;
    defparam GB_BUFFER_TVP_CLK_c_THRU_LUT4_0_LC_16_32_3.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_TVP_CLK_c_THRU_LUT4_0_LC_16_32_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_TVP_CLK_c_THRU_LUT4_0_LC_16_32_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20182),
            .lcout(GB_BUFFER_TVP_CLK_c_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i5_1_lut_rep_23_LC_17_9_6 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i5_1_lut_rep_23_LC_17_9_6 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i5_1_lut_rep_23_LC_17_9_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \receive_module.rx_counter.i5_1_lut_rep_23_LC_17_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18645),
            .lcout(\receive_module.rx_counter.n3790 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.X_242__i0_LC_17_10_0 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_242__i0_LC_17_10_0 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_242__i0_LC_17_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_242__i0_LC_17_10_0  (
            .in0(_gnd_net_),
            .in1(N__18622),
            .in2(_gnd_net_),
            .in3(N__18616),
            .lcout(\receive_module.rx_counter.n10 ),
            .ltout(),
            .carryin(bfn_17_10_0_),
            .carryout(\receive_module.rx_counter.n3301 ),
            .clk(N__20133),
            .ce(),
            .sr(N__19234));
    defparam \receive_module.rx_counter.X_242__i1_LC_17_10_1 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_242__i1_LC_17_10_1 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_242__i1_LC_17_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_242__i1_LC_17_10_1  (
            .in0(_gnd_net_),
            .in1(N__18613),
            .in2(_gnd_net_),
            .in3(N__18607),
            .lcout(\receive_module.rx_counter.n9 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3301 ),
            .carryout(\receive_module.rx_counter.n3302 ),
            .clk(N__20133),
            .ce(),
            .sr(N__19234));
    defparam \receive_module.rx_counter.X_242__i2_LC_17_10_2 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_242__i2_LC_17_10_2 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_242__i2_LC_17_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_242__i2_LC_17_10_2  (
            .in0(_gnd_net_),
            .in1(N__18604),
            .in2(_gnd_net_),
            .in3(N__18598),
            .lcout(\receive_module.rx_counter.n8 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3302 ),
            .carryout(\receive_module.rx_counter.n3303 ),
            .clk(N__20133),
            .ce(),
            .sr(N__19234));
    defparam \receive_module.rx_counter.X_242__i3_LC_17_10_3 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_242__i3_LC_17_10_3 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_242__i3_LC_17_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_242__i3_LC_17_10_3  (
            .in0(_gnd_net_),
            .in1(N__18595),
            .in2(_gnd_net_),
            .in3(N__18580),
            .lcout(\receive_module.rx_counter.X_3 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3303 ),
            .carryout(\receive_module.rx_counter.n3304 ),
            .clk(N__20133),
            .ce(),
            .sr(N__19234));
    defparam \receive_module.rx_counter.X_242__i4_LC_17_10_4 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_242__i4_LC_17_10_4 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_242__i4_LC_17_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_242__i4_LC_17_10_4  (
            .in0(_gnd_net_),
            .in1(N__19339),
            .in2(_gnd_net_),
            .in3(N__19324),
            .lcout(\receive_module.rx_counter.X_4 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3304 ),
            .carryout(\receive_module.rx_counter.n3305 ),
            .clk(N__20133),
            .ce(),
            .sr(N__19234));
    defparam \receive_module.rx_counter.X_242__i5_LC_17_10_5 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_242__i5_LC_17_10_5 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_242__i5_LC_17_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_242__i5_LC_17_10_5  (
            .in0(_gnd_net_),
            .in1(N__19321),
            .in2(_gnd_net_),
            .in3(N__19306),
            .lcout(\receive_module.rx_counter.X_5 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3305 ),
            .carryout(\receive_module.rx_counter.n3306 ),
            .clk(N__20133),
            .ce(),
            .sr(N__19234));
    defparam \receive_module.rx_counter.X_242__i6_LC_17_10_6 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_242__i6_LC_17_10_6 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_242__i6_LC_17_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_242__i6_LC_17_10_6  (
            .in0(_gnd_net_),
            .in1(N__19303),
            .in2(_gnd_net_),
            .in3(N__19288),
            .lcout(\receive_module.rx_counter.X_6 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3306 ),
            .carryout(\receive_module.rx_counter.n3307 ),
            .clk(N__20133),
            .ce(),
            .sr(N__19234));
    defparam \receive_module.rx_counter.X_242__i7_LC_17_10_7 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_242__i7_LC_17_10_7 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_242__i7_LC_17_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_242__i7_LC_17_10_7  (
            .in0(_gnd_net_),
            .in1(N__19285),
            .in2(_gnd_net_),
            .in3(N__19270),
            .lcout(\receive_module.rx_counter.X_7 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3307 ),
            .carryout(\receive_module.rx_counter.n3308 ),
            .clk(N__20133),
            .ce(),
            .sr(N__19234));
    defparam \receive_module.rx_counter.X_242__i8_LC_17_11_0 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_242__i8_LC_17_11_0 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_242__i8_LC_17_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_242__i8_LC_17_11_0  (
            .in0(_gnd_net_),
            .in1(N__19267),
            .in2(_gnd_net_),
            .in3(N__19255),
            .lcout(\receive_module.rx_counter.X_8 ),
            .ltout(),
            .carryin(bfn_17_11_0_),
            .carryout(\receive_module.rx_counter.n3309 ),
            .clk(N__20135),
            .ce(),
            .sr(N__19233));
    defparam \receive_module.rx_counter.X_242__i9_LC_17_11_1 .C_ON=1'b0;
    defparam \receive_module.rx_counter.X_242__i9_LC_17_11_1 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_242__i9_LC_17_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_242__i9_LC_17_11_1  (
            .in0(_gnd_net_),
            .in1(N__19248),
            .in2(_gnd_net_),
            .in3(N__19252),
            .lcout(\receive_module.rx_counter.X_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20135),
            .ce(),
            .sr(N__19233));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2407_LC_17_13_4 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2407_LC_17_13_4 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2407_LC_17_13_4 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_2407_LC_17_13_4  (
            .in0(N__23663),
            .in1(N__19213),
            .in2(N__22216),
            .in3(N__19204),
            .lcout(),
            .ltout(\line_buffer.n3734_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n3734_bdd_4_lut_LC_17_13_5 .C_ON=1'b0;
    defparam \line_buffer.n3734_bdd_4_lut_LC_17_13_5 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3734_bdd_4_lut_LC_17_13_5 .LUT_INIT=16'b1111000011001010;
    LogicCell40 \line_buffer.n3734_bdd_4_lut_LC_17_13_5  (
            .in0(N__19189),
            .in1(N__19174),
            .in2(N__19159),
            .in3(N__22178),
            .lcout(\line_buffer.n3737 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.Y_DELTA_PATTERN_i24_LC_17_14_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i24_LC_17_14_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i24_LC_17_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i24_LC_17_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19459),
            .lcout(\transmit_module.Y_DELTA_PATTERN_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22994),
            .ce(N__21482),
            .sr(N__21303));
    defparam \transmit_module.Y_DELTA_PATTERN_i12_LC_17_15_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i12_LC_17_15_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i12_LC_17_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i12_LC_17_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19447),
            .lcout(\transmit_module.Y_DELTA_PATTERN_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23073),
            .ce(N__21461),
            .sr(N__21171));
    defparam \transmit_module.Y_DELTA_PATTERN_i11_LC_17_15_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i11_LC_17_15_2 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i11_LC_17_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i11_LC_17_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19477),
            .lcout(\transmit_module.Y_DELTA_PATTERN_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23073),
            .ce(N__21461),
            .sr(N__21171));
    defparam \transmit_module.Y_DELTA_PATTERN_i25_LC_17_15_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i25_LC_17_15_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i25_LC_17_15_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i25_LC_17_15_3  (
            .in0(N__19453),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.Y_DELTA_PATTERN_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23073),
            .ce(N__21461),
            .sr(N__21171));
    defparam \transmit_module.Y_DELTA_PATTERN_i26_LC_17_15_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i26_LC_17_15_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i26_LC_17_15_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i26_LC_17_15_4  (
            .in0(N__19504),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.Y_DELTA_PATTERN_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23073),
            .ce(N__21461),
            .sr(N__21171));
    defparam \transmit_module.Y_DELTA_PATTERN_i13_LC_17_15_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i13_LC_17_15_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i13_LC_17_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i13_LC_17_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21565),
            .lcout(\transmit_module.Y_DELTA_PATTERN_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23073),
            .ce(N__21461),
            .sr(N__21171));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2417_LC_17_16_6 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2417_LC_17_16_6 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2417_LC_17_16_6 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_2417_LC_17_16_6  (
            .in0(N__23602),
            .in1(N__19441),
            .in2(N__22174),
            .in3(N__19429),
            .lcout(\line_buffer.n3746 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2351_3_lut_LC_17_17_3 .C_ON=1'b0;
    defparam \line_buffer.i2351_3_lut_LC_17_17_3 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2351_3_lut_LC_17_17_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \line_buffer.i2351_3_lut_LC_17_17_3  (
            .in0(N__23638),
            .in1(N__19408),
            .in2(_gnd_net_),
            .in3(N__19393),
            .lcout(\line_buffer.n3677 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2309_3_lut_LC_17_17_7 .C_ON=1'b0;
    defparam \line_buffer.i2309_3_lut_LC_17_17_7 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2309_3_lut_LC_17_17_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \line_buffer.i2309_3_lut_LC_17_17_7  (
            .in0(N__19372),
            .in1(N__23637),
            .in2(_gnd_net_),
            .in3(N__19360),
            .lcout(\line_buffer.n3635 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i5_LC_17_18_3 .C_ON=1'b0;
    defparam \line_buffer.dout_i5_LC_17_18_3 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i5_LC_17_18_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \line_buffer.dout_i5_LC_17_18_3  (
            .in0(N__21684),
            .in1(N__19969),
            .in2(_gnd_net_),
            .in3(N__19924),
            .lcout(TX_DATA_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22843),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n3698_bdd_4_lut_LC_17_19_6 .C_ON=1'b0;
    defparam \line_buffer.n3698_bdd_4_lut_LC_17_19_6 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3698_bdd_4_lut_LC_17_19_6 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \line_buffer.n3698_bdd_4_lut_LC_17_19_6  (
            .in0(N__19960),
            .in1(N__22179),
            .in2(N__19945),
            .in3(N__20803),
            .lcout(\line_buffer.n3701 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.VGA_R__i6_LC_17_22_3 .C_ON=1'b0;
    defparam \transmit_module.VGA_R__i6_LC_17_22_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.VGA_R__i6_LC_17_22_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.VGA_R__i6_LC_17_22_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19918),
            .lcout(n1793),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22690),
            .ce(),
            .sr(N__22320));
    defparam CONSTANT_ONE_LUT4_LC_17_25_3.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_17_25_3.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_17_25_3.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_17_25_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.Y_DELTA_PATTERN_i32_LC_18_13_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i32_LC_18_13_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i32_LC_18_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i32_LC_18_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19519),
            .lcout(\transmit_module.Y_DELTA_PATTERN_32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23105),
            .ce(N__21490),
            .sr(N__21260));
    defparam \transmit_module.Y_DELTA_PATTERN_i27_LC_18_13_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i27_LC_18_13_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i27_LC_18_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i27_LC_18_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19495),
            .lcout(\transmit_module.Y_DELTA_PATTERN_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23105),
            .ce(N__21490),
            .sr(N__21260));
    defparam \transmit_module.Y_DELTA_PATTERN_i28_LC_18_13_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i28_LC_18_13_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i28_LC_18_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i28_LC_18_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19489),
            .lcout(\transmit_module.Y_DELTA_PATTERN_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23105),
            .ce(N__21490),
            .sr(N__21260));
    defparam \transmit_module.Y_DELTA_PATTERN_i29_LC_18_13_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i29_LC_18_13_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i29_LC_18_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i29_LC_18_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19483),
            .lcout(\transmit_module.Y_DELTA_PATTERN_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23105),
            .ce(N__21490),
            .sr(N__21260));
    defparam \transmit_module.Y_DELTA_PATTERN_i30_LC_18_13_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i30_LC_18_13_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i30_LC_18_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i30_LC_18_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20017),
            .lcout(\transmit_module.Y_DELTA_PATTERN_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23105),
            .ce(N__21490),
            .sr(N__21260));
    defparam \transmit_module.Y_DELTA_PATTERN_i31_LC_18_13_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i31_LC_18_13_7 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i31_LC_18_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i31_LC_18_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20023),
            .lcout(\transmit_module.Y_DELTA_PATTERN_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23105),
            .ce(N__21490),
            .sr(N__21260));
    defparam \transmit_module.Y_DELTA_PATTERN_i22_LC_18_14_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i22_LC_18_14_2 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i22_LC_18_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i22_LC_18_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19999),
            .lcout(\transmit_module.Y_DELTA_PATTERN_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22996),
            .ce(N__21483),
            .sr(N__21301));
    defparam \transmit_module.Y_DELTA_PATTERN_i21_LC_18_14_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i21_LC_18_14_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i21_LC_18_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i21_LC_18_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20011),
            .lcout(\transmit_module.Y_DELTA_PATTERN_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22996),
            .ce(N__21483),
            .sr(N__21301));
    defparam \transmit_module.Y_DELTA_PATTERN_i23_LC_18_14_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i23_LC_18_14_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i23_LC_18_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i23_LC_18_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20005),
            .lcout(\transmit_module.Y_DELTA_PATTERN_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22996),
            .ce(N__21483),
            .sr(N__21301));
    defparam \transmit_module.Y_DELTA_PATTERN_i15_LC_18_15_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i15_LC_18_15_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i15_LC_18_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i15_LC_18_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19993),
            .lcout(\transmit_module.Y_DELTA_PATTERN_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22824),
            .ce(N__21453),
            .sr(N__21185));
    defparam \transmit_module.Y_DELTA_PATTERN_i19_LC_18_15_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i19_LC_18_15_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i19_LC_18_15_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i19_LC_18_15_3  (
            .in0(N__21496),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.Y_DELTA_PATTERN_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22824),
            .ce(N__21453),
            .sr(N__21185));
    defparam \transmit_module.Y_DELTA_PATTERN_i16_LC_18_15_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i16_LC_18_15_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i16_LC_18_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i16_LC_18_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19987),
            .lcout(\transmit_module.Y_DELTA_PATTERN_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22824),
            .ce(N__21453),
            .sr(N__21185));
    defparam \transmit_module.Y_DELTA_PATTERN_i17_LC_18_15_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i17_LC_18_15_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i17_LC_18_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i17_LC_18_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19975),
            .lcout(\transmit_module.Y_DELTA_PATTERN_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22824),
            .ce(N__21453),
            .sr(N__21185));
    defparam \transmit_module.Y_DELTA_PATTERN_i18_LC_18_15_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i18_LC_18_15_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i18_LC_18_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i18_LC_18_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19981),
            .lcout(\transmit_module.Y_DELTA_PATTERN_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22824),
            .ce(N__21453),
            .sr(N__21185));
    defparam \transmit_module.Y_DELTA_PATTERN_i14_LC_18_16_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i14_LC_18_16_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i14_LC_18_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i14_LC_18_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21571),
            .lcout(\transmit_module.Y_DELTA_PATTERN_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22947),
            .ce(N__21484),
            .sr(N__21302));
    defparam \transmit_module.VGA_R__i2_LC_18_21_4 .C_ON=1'b0;
    defparam \transmit_module.VGA_R__i2_LC_18_21_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.VGA_R__i2_LC_18_21_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.VGA_R__i2_LC_18_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20752),
            .lcout(n1797),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22751),
            .ce(),
            .sr(N__22322));
    defparam \transmit_module.Y_DELTA_PATTERN_i20_LC_19_14_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i20_LC_19_14_2 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i20_LC_19_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i20_LC_19_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21502),
            .lcout(\transmit_module.Y_DELTA_PATTERN_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22995),
            .ce(N__21489),
            .sr(N__21267));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2378_LC_19_15_1 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2378_LC_19_15_1 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2378_LC_19_15_1 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_2378_LC_19_15_1  (
            .in0(N__23647),
            .in1(N__20833),
            .in2(N__22217),
            .in3(N__20818),
            .lcout(\line_buffer.n3698 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n3692_bdd_4_lut_LC_19_17_5 .C_ON=1'b0;
    defparam \line_buffer.n3692_bdd_4_lut_LC_19_17_5 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3692_bdd_4_lut_LC_19_17_5 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \line_buffer.n3692_bdd_4_lut_LC_19_17_5  (
            .in0(N__20791),
            .in1(N__22186),
            .in2(N__20776),
            .in3(N__20704),
            .lcout(),
            .ltout(\line_buffer.n3695_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i1_LC_19_17_6 .C_ON=1'b0;
    defparam \line_buffer.dout_i1_LC_19_17_6 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i1_LC_19_17_6 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \line_buffer.dout_i1_LC_19_17_6  (
            .in0(_gnd_net_),
            .in1(N__21693),
            .in2(N__20755),
            .in3(N__21712),
            .lcout(TX_DATA_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22998),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2373_LC_19_18_7 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2373_LC_19_18_7 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2373_LC_19_18_7 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_2373_LC_19_18_7  (
            .in0(N__23653),
            .in1(N__20740),
            .in2(N__22218),
            .in3(N__20725),
            .lcout(\line_buffer.n3692 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.BRAM_ADDR__i3_LC_19_19_7 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i3_LC_19_19_7 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i3_LC_19_19_7 .LUT_INIT=16'b1101110010001100;
    LogicCell40 \receive_module.BRAM_ADDR__i3_LC_19_19_7  (
            .in0(N__20679),
            .in1(N__20584),
            .in2(N__20566),
            .in3(N__20209),
            .lcout(RX_ADDR_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__20153),
            .ce(),
            .sr(N__21989));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2402_LC_20_15_4 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2402_LC_20_15_4 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2402_LC_20_15_4 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_2402_LC_20_15_4  (
            .in0(N__23654),
            .in1(N__21904),
            .in2(N__22235),
            .in3(N__21892),
            .lcout(\line_buffer.n3710 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n3710_bdd_4_lut_LC_20_16_6 .C_ON=1'b0;
    defparam \line_buffer.n3710_bdd_4_lut_LC_20_16_6 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3710_bdd_4_lut_LC_20_16_6 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \line_buffer.n3710_bdd_4_lut_LC_20_16_6  (
            .in0(N__21883),
            .in1(N__22199),
            .in2(N__21868),
            .in3(N__21844),
            .lcout(\line_buffer.n3713 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2427_LC_20_17_0 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2427_LC_20_17_0 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2427_LC_20_17_0 .LUT_INIT=16'b1111100001011000;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_2427_LC_20_17_0  (
            .in0(N__22225),
            .in1(N__21838),
            .in2(N__23666),
            .in3(N__21820),
            .lcout(),
            .ltout(\line_buffer.n3758_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n3758_bdd_4_lut_LC_20_17_1 .C_ON=1'b0;
    defparam \line_buffer.n3758_bdd_4_lut_LC_20_17_1 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3758_bdd_4_lut_LC_20_17_1 .LUT_INIT=16'b1111000011001010;
    LogicCell40 \line_buffer.n3758_bdd_4_lut_LC_20_17_1  (
            .in0(N__21808),
            .in1(N__21790),
            .in2(N__21772),
            .in3(N__22227),
            .lcout(\line_buffer.n3761 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2412_LC_20_17_2 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2412_LC_20_17_2 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2412_LC_20_17_2 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_2412_LC_20_17_2  (
            .in0(N__23649),
            .in1(N__21769),
            .in2(N__22236),
            .in3(N__21757),
            .lcout(),
            .ltout(\line_buffer.n3740_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n3740_bdd_4_lut_LC_20_17_3 .C_ON=1'b0;
    defparam \line_buffer.n3740_bdd_4_lut_LC_20_17_3 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3740_bdd_4_lut_LC_20_17_3 .LUT_INIT=16'b1111000011001010;
    LogicCell40 \line_buffer.n3740_bdd_4_lut_LC_20_17_3  (
            .in0(N__21748),
            .in1(N__21730),
            .in2(N__21715),
            .in3(N__22226),
            .lcout(\line_buffer.n3743 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i3_LC_20_17_5 .C_ON=1'b0;
    defparam \line_buffer.dout_i3_LC_20_17_5 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i3_LC_20_17_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \line_buffer.dout_i3_LC_20_17_5  (
            .in0(N__21691),
            .in1(N__21706),
            .in2(_gnd_net_),
            .in3(N__21700),
            .lcout(TX_DATA_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23096),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i7_LC_20_18_2 .C_ON=1'b0;
    defparam \line_buffer.dout_i7_LC_20_18_2 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i7_LC_20_18_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \line_buffer.dout_i7_LC_20_18_2  (
            .in0(N__21692),
            .in1(N__21580),
            .in2(_gnd_net_),
            .in3(N__22003),
            .lcout(TX_DATA_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22981),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2383_LC_20_19_1 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2383_LC_20_19_1 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2383_LC_20_19_1 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_2383_LC_20_19_1  (
            .in0(N__23648),
            .in1(N__23473),
            .in2(N__22237),
            .in3(N__23458),
            .lcout(\line_buffer.n3704 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.VGA_R__i4_LC_20_20_3 .C_ON=1'b0;
    defparam \transmit_module.VGA_R__i4_LC_20_20_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.VGA_R__i4_LC_20_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.VGA_R__i4_LC_20_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23443),
            .lcout(n1795),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22980),
            .ce(),
            .sr(N__22326));
    defparam \transmit_module.VGA_R__i8_LC_20_22_3 .C_ON=1'b0;
    defparam \transmit_module.VGA_R__i8_LC_20_22_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.VGA_R__i8_LC_20_22_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \transmit_module.VGA_R__i8_LC_20_22_3  (
            .in0(N__23374),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(ADV_B_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22832),
            .ce(),
            .sr(N__22327));
    defparam \line_buffer.n3704_bdd_4_lut_LC_21_19_7 .C_ON=1'b0;
    defparam \line_buffer.n3704_bdd_4_lut_LC_21_19_7 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3704_bdd_4_lut_LC_21_19_7 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \line_buffer.n3704_bdd_4_lut_LC_21_19_7  (
            .in0(N__22252),
            .in1(N__22231),
            .in2(N__22030),
            .in3(N__22009),
            .lcout(\line_buffer.n3707 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // main
