// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     Oct 7 2018 23:14:10

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "main" view "INTERFACE"

module main (
    TVP_VIDEO,
    ADV_B,
    ADV_G,
    ADV_R,
    DEBUG,
    TVP_CLK,
    ADV_CLK,
    TVP_HSYNC,
    ADV_HSYNC,
    TVP_VSYNC,
    ADV_VSYNC,
    ADV_BLANK_N,
    LED,
    ADV_SYNC_N);

    input [9:0] TVP_VIDEO;
    output [7:0] ADV_B;
    output [7:0] ADV_G;
    output [7:0] ADV_R;
    inout [7:0] DEBUG;
    input TVP_CLK;
    output ADV_CLK;
    input TVP_HSYNC;
    output ADV_HSYNC;
    input TVP_VSYNC;
    output ADV_VSYNC;
    output ADV_BLANK_N;
    output LED;
    output ADV_SYNC_N;

    wire N__24834;
    wire N__24833;
    wire N__24832;
    wire N__24823;
    wire N__24822;
    wire N__24821;
    wire N__24814;
    wire N__24813;
    wire N__24812;
    wire N__24805;
    wire N__24804;
    wire N__24803;
    wire N__24796;
    wire N__24795;
    wire N__24794;
    wire N__24787;
    wire N__24786;
    wire N__24785;
    wire N__24778;
    wire N__24777;
    wire N__24776;
    wire N__24769;
    wire N__24768;
    wire N__24767;
    wire N__24760;
    wire N__24759;
    wire N__24758;
    wire N__24751;
    wire N__24750;
    wire N__24749;
    wire N__24742;
    wire N__24741;
    wire N__24740;
    wire N__24733;
    wire N__24732;
    wire N__24731;
    wire N__24724;
    wire N__24723;
    wire N__24722;
    wire N__24715;
    wire N__24714;
    wire N__24713;
    wire N__24706;
    wire N__24705;
    wire N__24704;
    wire N__24697;
    wire N__24696;
    wire N__24695;
    wire N__24688;
    wire N__24687;
    wire N__24686;
    wire N__24679;
    wire N__24678;
    wire N__24677;
    wire N__24670;
    wire N__24669;
    wire N__24668;
    wire N__24661;
    wire N__24660;
    wire N__24659;
    wire N__24652;
    wire N__24651;
    wire N__24650;
    wire N__24643;
    wire N__24642;
    wire N__24641;
    wire N__24634;
    wire N__24633;
    wire N__24632;
    wire N__24625;
    wire N__24624;
    wire N__24623;
    wire N__24616;
    wire N__24615;
    wire N__24614;
    wire N__24607;
    wire N__24606;
    wire N__24605;
    wire N__24598;
    wire N__24597;
    wire N__24596;
    wire N__24589;
    wire N__24588;
    wire N__24587;
    wire N__24580;
    wire N__24579;
    wire N__24578;
    wire N__24571;
    wire N__24570;
    wire N__24569;
    wire N__24562;
    wire N__24561;
    wire N__24560;
    wire N__24553;
    wire N__24552;
    wire N__24551;
    wire N__24544;
    wire N__24543;
    wire N__24542;
    wire N__24535;
    wire N__24534;
    wire N__24533;
    wire N__24526;
    wire N__24525;
    wire N__24524;
    wire N__24517;
    wire N__24516;
    wire N__24515;
    wire N__24508;
    wire N__24507;
    wire N__24506;
    wire N__24499;
    wire N__24498;
    wire N__24497;
    wire N__24490;
    wire N__24489;
    wire N__24488;
    wire N__24481;
    wire N__24480;
    wire N__24479;
    wire N__24472;
    wire N__24471;
    wire N__24470;
    wire N__24463;
    wire N__24462;
    wire N__24461;
    wire N__24454;
    wire N__24453;
    wire N__24452;
    wire N__24445;
    wire N__24444;
    wire N__24443;
    wire N__24436;
    wire N__24435;
    wire N__24434;
    wire N__24427;
    wire N__24426;
    wire N__24425;
    wire N__24418;
    wire N__24417;
    wire N__24416;
    wire N__24409;
    wire N__24408;
    wire N__24407;
    wire N__24400;
    wire N__24399;
    wire N__24398;
    wire N__24381;
    wire N__24378;
    wire N__24375;
    wire N__24372;
    wire N__24369;
    wire N__24366;
    wire N__24363;
    wire N__24362;
    wire N__24359;
    wire N__24356;
    wire N__24355;
    wire N__24354;
    wire N__24353;
    wire N__24352;
    wire N__24351;
    wire N__24350;
    wire N__24349;
    wire N__24344;
    wire N__24341;
    wire N__24338;
    wire N__24337;
    wire N__24336;
    wire N__24335;
    wire N__24334;
    wire N__24333;
    wire N__24332;
    wire N__24331;
    wire N__24328;
    wire N__24325;
    wire N__24322;
    wire N__24319;
    wire N__24316;
    wire N__24315;
    wire N__24314;
    wire N__24313;
    wire N__24312;
    wire N__24305;
    wire N__24302;
    wire N__24301;
    wire N__24300;
    wire N__24299;
    wire N__24296;
    wire N__24295;
    wire N__24294;
    wire N__24293;
    wire N__24292;
    wire N__24291;
    wire N__24288;
    wire N__24287;
    wire N__24284;
    wire N__24283;
    wire N__24280;
    wire N__24277;
    wire N__24274;
    wire N__24273;
    wire N__24272;
    wire N__24271;
    wire N__24270;
    wire N__24267;
    wire N__24258;
    wire N__24255;
    wire N__24252;
    wire N__24251;
    wire N__24250;
    wire N__24249;
    wire N__24248;
    wire N__24245;
    wire N__24242;
    wire N__24241;
    wire N__24236;
    wire N__24233;
    wire N__24230;
    wire N__24229;
    wire N__24228;
    wire N__24227;
    wire N__24224;
    wire N__24223;
    wire N__24222;
    wire N__24221;
    wire N__24220;
    wire N__24217;
    wire N__24214;
    wire N__24213;
    wire N__24210;
    wire N__24209;
    wire N__24208;
    wire N__24205;
    wire N__24204;
    wire N__24201;
    wire N__24198;
    wire N__24197;
    wire N__24194;
    wire N__24191;
    wire N__24188;
    wire N__24185;
    wire N__24184;
    wire N__24181;
    wire N__24176;
    wire N__24173;
    wire N__24170;
    wire N__24167;
    wire N__24164;
    wire N__24159;
    wire N__24156;
    wire N__24153;
    wire N__24150;
    wire N__24147;
    wire N__24146;
    wire N__24143;
    wire N__24140;
    wire N__24139;
    wire N__24138;
    wire N__24133;
    wire N__24130;
    wire N__24125;
    wire N__24122;
    wire N__24119;
    wire N__24116;
    wire N__24115;
    wire N__24114;
    wire N__24113;
    wire N__24112;
    wire N__24109;
    wire N__24106;
    wire N__24103;
    wire N__24102;
    wire N__24099;
    wire N__24096;
    wire N__24093;
    wire N__24092;
    wire N__24087;
    wire N__24084;
    wire N__24081;
    wire N__24078;
    wire N__24075;
    wire N__24074;
    wire N__24071;
    wire N__24068;
    wire N__24067;
    wire N__24066;
    wire N__24065;
    wire N__24064;
    wire N__24061;
    wire N__24058;
    wire N__24055;
    wire N__24050;
    wire N__24045;
    wire N__24042;
    wire N__24033;
    wire N__24028;
    wire N__24017;
    wire N__24014;
    wire N__24011;
    wire N__24008;
    wire N__24005;
    wire N__24002;
    wire N__24001;
    wire N__23996;
    wire N__23987;
    wire N__23984;
    wire N__23981;
    wire N__23980;
    wire N__23979;
    wire N__23978;
    wire N__23977;
    wire N__23974;
    wire N__23973;
    wire N__23972;
    wire N__23969;
    wire N__23966;
    wire N__23961;
    wire N__23958;
    wire N__23957;
    wire N__23952;
    wire N__23951;
    wire N__23950;
    wire N__23949;
    wire N__23948;
    wire N__23945;
    wire N__23942;
    wire N__23937;
    wire N__23934;
    wire N__23931;
    wire N__23928;
    wire N__23925;
    wire N__23920;
    wire N__23917;
    wire N__23914;
    wire N__23911;
    wire N__23910;
    wire N__23909;
    wire N__23906;
    wire N__23899;
    wire N__23892;
    wire N__23883;
    wire N__23876;
    wire N__23873;
    wire N__23870;
    wire N__23869;
    wire N__23862;
    wire N__23859;
    wire N__23856;
    wire N__23853;
    wire N__23852;
    wire N__23849;
    wire N__23846;
    wire N__23845;
    wire N__23842;
    wire N__23839;
    wire N__23836;
    wire N__23835;
    wire N__23832;
    wire N__23825;
    wire N__23822;
    wire N__23819;
    wire N__23816;
    wire N__23815;
    wire N__23812;
    wire N__23811;
    wire N__23808;
    wire N__23807;
    wire N__23804;
    wire N__23799;
    wire N__23798;
    wire N__23795;
    wire N__23786;
    wire N__23779;
    wire N__23776;
    wire N__23773;
    wire N__23772;
    wire N__23771;
    wire N__23768;
    wire N__23765;
    wire N__23764;
    wire N__23759;
    wire N__23756;
    wire N__23749;
    wire N__23746;
    wire N__23745;
    wire N__23742;
    wire N__23739;
    wire N__23736;
    wire N__23735;
    wire N__23732;
    wire N__23729;
    wire N__23726;
    wire N__23723;
    wire N__23720;
    wire N__23713;
    wire N__23710;
    wire N__23705;
    wire N__23702;
    wire N__23697;
    wire N__23694;
    wire N__23691;
    wire N__23688;
    wire N__23685;
    wire N__23682;
    wire N__23681;
    wire N__23678;
    wire N__23675;
    wire N__23672;
    wire N__23665;
    wire N__23660;
    wire N__23657;
    wire N__23654;
    wire N__23653;
    wire N__23650;
    wire N__23647;
    wire N__23644;
    wire N__23643;
    wire N__23640;
    wire N__23637;
    wire N__23634;
    wire N__23631;
    wire N__23628;
    wire N__23625;
    wire N__23620;
    wire N__23617;
    wire N__23616;
    wire N__23611;
    wire N__23604;
    wire N__23599;
    wire N__23590;
    wire N__23587;
    wire N__23584;
    wire N__23579;
    wire N__23576;
    wire N__23573;
    wire N__23568;
    wire N__23559;
    wire N__23556;
    wire N__23553;
    wire N__23550;
    wire N__23547;
    wire N__23544;
    wire N__23541;
    wire N__23538;
    wire N__23533;
    wire N__23530;
    wire N__23527;
    wire N__23522;
    wire N__23519;
    wire N__23516;
    wire N__23509;
    wire N__23504;
    wire N__23499;
    wire N__23490;
    wire N__23483;
    wire N__23480;
    wire N__23477;
    wire N__23474;
    wire N__23469;
    wire N__23464;
    wire N__23461;
    wire N__23458;
    wire N__23455;
    wire N__23452;
    wire N__23449;
    wire N__23446;
    wire N__23443;
    wire N__23440;
    wire N__23437;
    wire N__23434;
    wire N__23425;
    wire N__23422;
    wire N__23415;
    wire N__23410;
    wire N__23397;
    wire N__23396;
    wire N__23395;
    wire N__23392;
    wire N__23391;
    wire N__23388;
    wire N__23387;
    wire N__23384;
    wire N__23381;
    wire N__23378;
    wire N__23375;
    wire N__23372;
    wire N__23369;
    wire N__23364;
    wire N__23359;
    wire N__23356;
    wire N__23351;
    wire N__23346;
    wire N__23343;
    wire N__23340;
    wire N__23337;
    wire N__23336;
    wire N__23335;
    wire N__23334;
    wire N__23333;
    wire N__23332;
    wire N__23331;
    wire N__23328;
    wire N__23327;
    wire N__23326;
    wire N__23325;
    wire N__23324;
    wire N__23323;
    wire N__23320;
    wire N__23317;
    wire N__23314;
    wire N__23311;
    wire N__23310;
    wire N__23307;
    wire N__23304;
    wire N__23303;
    wire N__23302;
    wire N__23301;
    wire N__23300;
    wire N__23299;
    wire N__23298;
    wire N__23297;
    wire N__23296;
    wire N__23293;
    wire N__23290;
    wire N__23287;
    wire N__23286;
    wire N__23285;
    wire N__23284;
    wire N__23283;
    wire N__23282;
    wire N__23281;
    wire N__23280;
    wire N__23277;
    wire N__23276;
    wire N__23275;
    wire N__23274;
    wire N__23271;
    wire N__23268;
    wire N__23265;
    wire N__23262;
    wire N__23257;
    wire N__23254;
    wire N__23253;
    wire N__23252;
    wire N__23247;
    wire N__23244;
    wire N__23243;
    wire N__23242;
    wire N__23241;
    wire N__23240;
    wire N__23239;
    wire N__23238;
    wire N__23235;
    wire N__23234;
    wire N__23233;
    wire N__23230;
    wire N__23229;
    wire N__23228;
    wire N__23225;
    wire N__23224;
    wire N__23223;
    wire N__23220;
    wire N__23217;
    wire N__23214;
    wire N__23213;
    wire N__23212;
    wire N__23209;
    wire N__23202;
    wire N__23199;
    wire N__23198;
    wire N__23197;
    wire N__23196;
    wire N__23193;
    wire N__23190;
    wire N__23187;
    wire N__23184;
    wire N__23181;
    wire N__23178;
    wire N__23175;
    wire N__23174;
    wire N__23171;
    wire N__23168;
    wire N__23165;
    wire N__23158;
    wire N__23151;
    wire N__23148;
    wire N__23145;
    wire N__23144;
    wire N__23143;
    wire N__23142;
    wire N__23141;
    wire N__23140;
    wire N__23135;
    wire N__23132;
    wire N__23129;
    wire N__23126;
    wire N__23125;
    wire N__23122;
    wire N__23121;
    wire N__23120;
    wire N__23119;
    wire N__23116;
    wire N__23111;
    wire N__23108;
    wire N__23101;
    wire N__23098;
    wire N__23095;
    wire N__23092;
    wire N__23091;
    wire N__23088;
    wire N__23083;
    wire N__23080;
    wire N__23075;
    wire N__23068;
    wire N__23065;
    wire N__23062;
    wire N__23059;
    wire N__23056;
    wire N__23053;
    wire N__23050;
    wire N__23047;
    wire N__23040;
    wire N__23037;
    wire N__23034;
    wire N__23031;
    wire N__23026;
    wire N__23025;
    wire N__23024;
    wire N__23019;
    wire N__23016;
    wire N__23007;
    wire N__23004;
    wire N__23001;
    wire N__22998;
    wire N__22991;
    wire N__22982;
    wire N__22973;
    wire N__22970;
    wire N__22965;
    wire N__22960;
    wire N__22951;
    wire N__22946;
    wire N__22941;
    wire N__22932;
    wire N__22929;
    wire N__22922;
    wire N__22917;
    wire N__22910;
    wire N__22897;
    wire N__22888;
    wire N__22869;
    wire N__22866;
    wire N__22863;
    wire N__22860;
    wire N__22857;
    wire N__22854;
    wire N__22851;
    wire N__22848;
    wire N__22845;
    wire N__22842;
    wire N__22839;
    wire N__22836;
    wire N__22833;
    wire N__22832;
    wire N__22831;
    wire N__22830;
    wire N__22829;
    wire N__22828;
    wire N__22827;
    wire N__22826;
    wire N__22825;
    wire N__22822;
    wire N__22821;
    wire N__22818;
    wire N__22815;
    wire N__22812;
    wire N__22809;
    wire N__22808;
    wire N__22807;
    wire N__22804;
    wire N__22799;
    wire N__22798;
    wire N__22795;
    wire N__22792;
    wire N__22789;
    wire N__22786;
    wire N__22783;
    wire N__22778;
    wire N__22775;
    wire N__22772;
    wire N__22771;
    wire N__22770;
    wire N__22769;
    wire N__22768;
    wire N__22767;
    wire N__22764;
    wire N__22763;
    wire N__22760;
    wire N__22759;
    wire N__22756;
    wire N__22755;
    wire N__22754;
    wire N__22753;
    wire N__22748;
    wire N__22745;
    wire N__22736;
    wire N__22733;
    wire N__22730;
    wire N__22727;
    wire N__22724;
    wire N__22723;
    wire N__22720;
    wire N__22717;
    wire N__22714;
    wire N__22711;
    wire N__22708;
    wire N__22707;
    wire N__22704;
    wire N__22701;
    wire N__22698;
    wire N__22695;
    wire N__22692;
    wire N__22689;
    wire N__22684;
    wire N__22675;
    wire N__22672;
    wire N__22669;
    wire N__22662;
    wire N__22659;
    wire N__22656;
    wire N__22651;
    wire N__22648;
    wire N__22643;
    wire N__22634;
    wire N__22633;
    wire N__22620;
    wire N__22617;
    wire N__22614;
    wire N__22611;
    wire N__22602;
    wire N__22599;
    wire N__22596;
    wire N__22593;
    wire N__22590;
    wire N__22587;
    wire N__22584;
    wire N__22581;
    wire N__22578;
    wire N__22575;
    wire N__22572;
    wire N__22569;
    wire N__22566;
    wire N__22563;
    wire N__22560;
    wire N__22557;
    wire N__22554;
    wire N__22551;
    wire N__22548;
    wire N__22545;
    wire N__22542;
    wire N__22539;
    wire N__22538;
    wire N__22535;
    wire N__22532;
    wire N__22531;
    wire N__22526;
    wire N__22523;
    wire N__22520;
    wire N__22517;
    wire N__22514;
    wire N__22511;
    wire N__22508;
    wire N__22505;
    wire N__22502;
    wire N__22499;
    wire N__22494;
    wire N__22491;
    wire N__22488;
    wire N__22485;
    wire N__22482;
    wire N__22481;
    wire N__22478;
    wire N__22477;
    wire N__22474;
    wire N__22471;
    wire N__22468;
    wire N__22465;
    wire N__22462;
    wire N__22459;
    wire N__22456;
    wire N__22451;
    wire N__22448;
    wire N__22445;
    wire N__22442;
    wire N__22439;
    wire N__22434;
    wire N__22431;
    wire N__22428;
    wire N__22427;
    wire N__22426;
    wire N__22425;
    wire N__22424;
    wire N__22421;
    wire N__22418;
    wire N__22415;
    wire N__22414;
    wire N__22411;
    wire N__22408;
    wire N__22401;
    wire N__22398;
    wire N__22397;
    wire N__22394;
    wire N__22391;
    wire N__22386;
    wire N__22383;
    wire N__22380;
    wire N__22377;
    wire N__22374;
    wire N__22371;
    wire N__22362;
    wire N__22359;
    wire N__22356;
    wire N__22353;
    wire N__22350;
    wire N__22347;
    wire N__22344;
    wire N__22341;
    wire N__22338;
    wire N__22335;
    wire N__22332;
    wire N__22329;
    wire N__22326;
    wire N__22323;
    wire N__22322;
    wire N__22319;
    wire N__22316;
    wire N__22315;
    wire N__22310;
    wire N__22307;
    wire N__22306;
    wire N__22301;
    wire N__22298;
    wire N__22297;
    wire N__22292;
    wire N__22289;
    wire N__22288;
    wire N__22283;
    wire N__22280;
    wire N__22279;
    wire N__22274;
    wire N__22271;
    wire N__22270;
    wire N__22269;
    wire N__22264;
    wire N__22261;
    wire N__22260;
    wire N__22257;
    wire N__22256;
    wire N__22255;
    wire N__22250;
    wire N__22247;
    wire N__22246;
    wire N__22243;
    wire N__22240;
    wire N__22237;
    wire N__22236;
    wire N__22235;
    wire N__22230;
    wire N__22227;
    wire N__22226;
    wire N__22219;
    wire N__22216;
    wire N__22213;
    wire N__22212;
    wire N__22211;
    wire N__22206;
    wire N__22203;
    wire N__22202;
    wire N__22195;
    wire N__22192;
    wire N__22189;
    wire N__22188;
    wire N__22187;
    wire N__22182;
    wire N__22179;
    wire N__22178;
    wire N__22171;
    wire N__22168;
    wire N__22165;
    wire N__22164;
    wire N__22163;
    wire N__22158;
    wire N__22155;
    wire N__22154;
    wire N__22153;
    wire N__22146;
    wire N__22143;
    wire N__22140;
    wire N__22139;
    wire N__22138;
    wire N__22133;
    wire N__22130;
    wire N__22127;
    wire N__22126;
    wire N__22119;
    wire N__22116;
    wire N__22113;
    wire N__22112;
    wire N__22111;
    wire N__22106;
    wire N__22103;
    wire N__22100;
    wire N__22099;
    wire N__22092;
    wire N__22089;
    wire N__22086;
    wire N__22079;
    wire N__22076;
    wire N__22071;
    wire N__22068;
    wire N__22065;
    wire N__22064;
    wire N__22061;
    wire N__22060;
    wire N__22055;
    wire N__22052;
    wire N__22049;
    wire N__22046;
    wire N__22043;
    wire N__22040;
    wire N__22031;
    wire N__22026;
    wire N__22023;
    wire N__22020;
    wire N__22017;
    wire N__22014;
    wire N__22011;
    wire N__22008;
    wire N__22005;
    wire N__22002;
    wire N__21999;
    wire N__21996;
    wire N__21995;
    wire N__21994;
    wire N__21993;
    wire N__21992;
    wire N__21991;
    wire N__21990;
    wire N__21989;
    wire N__21988;
    wire N__21987;
    wire N__21986;
    wire N__21985;
    wire N__21984;
    wire N__21983;
    wire N__21982;
    wire N__21981;
    wire N__21978;
    wire N__21977;
    wire N__21976;
    wire N__21975;
    wire N__21974;
    wire N__21973;
    wire N__21972;
    wire N__21971;
    wire N__21970;
    wire N__21969;
    wire N__21968;
    wire N__21967;
    wire N__21966;
    wire N__21965;
    wire N__21964;
    wire N__21963;
    wire N__21962;
    wire N__21961;
    wire N__21960;
    wire N__21959;
    wire N__21958;
    wire N__21957;
    wire N__21956;
    wire N__21955;
    wire N__21954;
    wire N__21953;
    wire N__21952;
    wire N__21951;
    wire N__21950;
    wire N__21949;
    wire N__21948;
    wire N__21947;
    wire N__21946;
    wire N__21945;
    wire N__21944;
    wire N__21943;
    wire N__21942;
    wire N__21941;
    wire N__21940;
    wire N__21939;
    wire N__21938;
    wire N__21937;
    wire N__21936;
    wire N__21935;
    wire N__21934;
    wire N__21933;
    wire N__21932;
    wire N__21931;
    wire N__21930;
    wire N__21929;
    wire N__21928;
    wire N__21927;
    wire N__21926;
    wire N__21789;
    wire N__21786;
    wire N__21783;
    wire N__21780;
    wire N__21777;
    wire N__21774;
    wire N__21771;
    wire N__21768;
    wire N__21765;
    wire N__21762;
    wire N__21759;
    wire N__21756;
    wire N__21753;
    wire N__21750;
    wire N__21747;
    wire N__21744;
    wire N__21741;
    wire N__21738;
    wire N__21737;
    wire N__21734;
    wire N__21731;
    wire N__21728;
    wire N__21727;
    wire N__21726;
    wire N__21725;
    wire N__21724;
    wire N__21721;
    wire N__21718;
    wire N__21715;
    wire N__21714;
    wire N__21711;
    wire N__21708;
    wire N__21705;
    wire N__21704;
    wire N__21701;
    wire N__21696;
    wire N__21693;
    wire N__21692;
    wire N__21689;
    wire N__21686;
    wire N__21683;
    wire N__21680;
    wire N__21673;
    wire N__21670;
    wire N__21667;
    wire N__21664;
    wire N__21659;
    wire N__21656;
    wire N__21653;
    wire N__21650;
    wire N__21645;
    wire N__21640;
    wire N__21633;
    wire N__21630;
    wire N__21627;
    wire N__21624;
    wire N__21623;
    wire N__21620;
    wire N__21617;
    wire N__21614;
    wire N__21611;
    wire N__21608;
    wire N__21605;
    wire N__21602;
    wire N__21599;
    wire N__21596;
    wire N__21593;
    wire N__21588;
    wire N__21585;
    wire N__21582;
    wire N__21579;
    wire N__21576;
    wire N__21573;
    wire N__21570;
    wire N__21567;
    wire N__21564;
    wire N__21561;
    wire N__21558;
    wire N__21555;
    wire N__21552;
    wire N__21549;
    wire N__21546;
    wire N__21543;
    wire N__21540;
    wire N__21537;
    wire N__21534;
    wire N__21531;
    wire N__21528;
    wire N__21525;
    wire N__21522;
    wire N__21519;
    wire N__21516;
    wire N__21513;
    wire N__21510;
    wire N__21507;
    wire N__21506;
    wire N__21505;
    wire N__21504;
    wire N__21503;
    wire N__21502;
    wire N__21501;
    wire N__21500;
    wire N__21499;
    wire N__21498;
    wire N__21497;
    wire N__21494;
    wire N__21491;
    wire N__21488;
    wire N__21485;
    wire N__21484;
    wire N__21483;
    wire N__21480;
    wire N__21479;
    wire N__21478;
    wire N__21475;
    wire N__21474;
    wire N__21471;
    wire N__21468;
    wire N__21465;
    wire N__21464;
    wire N__21463;
    wire N__21460;
    wire N__21459;
    wire N__21458;
    wire N__21455;
    wire N__21452;
    wire N__21449;
    wire N__21446;
    wire N__21443;
    wire N__21440;
    wire N__21439;
    wire N__21436;
    wire N__21433;
    wire N__21426;
    wire N__21421;
    wire N__21418;
    wire N__21415;
    wire N__21414;
    wire N__21411;
    wire N__21408;
    wire N__21405;
    wire N__21402;
    wire N__21397;
    wire N__21394;
    wire N__21389;
    wire N__21386;
    wire N__21383;
    wire N__21380;
    wire N__21367;
    wire N__21362;
    wire N__21359;
    wire N__21356;
    wire N__21351;
    wire N__21344;
    wire N__21337;
    wire N__21324;
    wire N__21321;
    wire N__21318;
    wire N__21315;
    wire N__21312;
    wire N__21309;
    wire N__21306;
    wire N__21305;
    wire N__21304;
    wire N__21301;
    wire N__21300;
    wire N__21299;
    wire N__21296;
    wire N__21295;
    wire N__21294;
    wire N__21293;
    wire N__21290;
    wire N__21287;
    wire N__21284;
    wire N__21283;
    wire N__21280;
    wire N__21277;
    wire N__21274;
    wire N__21271;
    wire N__21270;
    wire N__21269;
    wire N__21268;
    wire N__21267;
    wire N__21264;
    wire N__21261;
    wire N__21258;
    wire N__21255;
    wire N__21252;
    wire N__21249;
    wire N__21246;
    wire N__21243;
    wire N__21240;
    wire N__21237;
    wire N__21232;
    wire N__21229;
    wire N__21228;
    wire N__21225;
    wire N__21220;
    wire N__21217;
    wire N__21212;
    wire N__21207;
    wire N__21202;
    wire N__21197;
    wire N__21194;
    wire N__21189;
    wire N__21186;
    wire N__21181;
    wire N__21174;
    wire N__21165;
    wire N__21162;
    wire N__21159;
    wire N__21156;
    wire N__21153;
    wire N__21150;
    wire N__21147;
    wire N__21144;
    wire N__21141;
    wire N__21138;
    wire N__21135;
    wire N__21132;
    wire N__21129;
    wire N__21126;
    wire N__21123;
    wire N__21120;
    wire N__21117;
    wire N__21114;
    wire N__21111;
    wire N__21108;
    wire N__21105;
    wire N__21102;
    wire N__21099;
    wire N__21096;
    wire N__21093;
    wire N__21090;
    wire N__21087;
    wire N__21084;
    wire N__21081;
    wire N__21078;
    wire N__21075;
    wire N__21072;
    wire N__21069;
    wire N__21066;
    wire N__21063;
    wire N__21060;
    wire N__21057;
    wire N__21054;
    wire N__21053;
    wire N__21052;
    wire N__21051;
    wire N__21050;
    wire N__21049;
    wire N__21046;
    wire N__21043;
    wire N__21040;
    wire N__21037;
    wire N__21034;
    wire N__21033;
    wire N__21030;
    wire N__21029;
    wire N__21026;
    wire N__21017;
    wire N__21014;
    wire N__21011;
    wire N__21008;
    wire N__21007;
    wire N__21004;
    wire N__20999;
    wire N__20994;
    wire N__20991;
    wire N__20988;
    wire N__20985;
    wire N__20982;
    wire N__20979;
    wire N__20974;
    wire N__20971;
    wire N__20968;
    wire N__20961;
    wire N__20958;
    wire N__20955;
    wire N__20952;
    wire N__20949;
    wire N__20946;
    wire N__20943;
    wire N__20940;
    wire N__20937;
    wire N__20934;
    wire N__20931;
    wire N__20928;
    wire N__20925;
    wire N__20922;
    wire N__20919;
    wire N__20916;
    wire N__20913;
    wire N__20910;
    wire N__20907;
    wire N__20904;
    wire N__20901;
    wire N__20898;
    wire N__20895;
    wire N__20892;
    wire N__20889;
    wire N__20886;
    wire N__20883;
    wire N__20880;
    wire N__20877;
    wire N__20874;
    wire N__20871;
    wire N__20868;
    wire N__20865;
    wire N__20862;
    wire N__20859;
    wire N__20856;
    wire N__20853;
    wire N__20850;
    wire N__20847;
    wire N__20844;
    wire N__20841;
    wire N__20838;
    wire N__20835;
    wire N__20832;
    wire N__20829;
    wire N__20826;
    wire N__20823;
    wire N__20820;
    wire N__20817;
    wire N__20814;
    wire N__20811;
    wire N__20808;
    wire N__20805;
    wire N__20802;
    wire N__20799;
    wire N__20796;
    wire N__20793;
    wire N__20790;
    wire N__20787;
    wire N__20784;
    wire N__20781;
    wire N__20778;
    wire N__20775;
    wire N__20772;
    wire N__20769;
    wire N__20766;
    wire N__20763;
    wire N__20762;
    wire N__20759;
    wire N__20756;
    wire N__20753;
    wire N__20750;
    wire N__20747;
    wire N__20744;
    wire N__20743;
    wire N__20740;
    wire N__20737;
    wire N__20734;
    wire N__20731;
    wire N__20728;
    wire N__20725;
    wire N__20720;
    wire N__20717;
    wire N__20714;
    wire N__20709;
    wire N__20706;
    wire N__20703;
    wire N__20700;
    wire N__20697;
    wire N__20696;
    wire N__20693;
    wire N__20690;
    wire N__20687;
    wire N__20684;
    wire N__20679;
    wire N__20678;
    wire N__20675;
    wire N__20672;
    wire N__20669;
    wire N__20666;
    wire N__20661;
    wire N__20658;
    wire N__20655;
    wire N__20652;
    wire N__20649;
    wire N__20646;
    wire N__20643;
    wire N__20640;
    wire N__20637;
    wire N__20634;
    wire N__20633;
    wire N__20630;
    wire N__20629;
    wire N__20628;
    wire N__20627;
    wire N__20626;
    wire N__20625;
    wire N__20622;
    wire N__20619;
    wire N__20614;
    wire N__20609;
    wire N__20606;
    wire N__20605;
    wire N__20604;
    wire N__20601;
    wire N__20596;
    wire N__20593;
    wire N__20592;
    wire N__20591;
    wire N__20590;
    wire N__20587;
    wire N__20584;
    wire N__20581;
    wire N__20580;
    wire N__20579;
    wire N__20576;
    wire N__20573;
    wire N__20570;
    wire N__20567;
    wire N__20564;
    wire N__20561;
    wire N__20554;
    wire N__20549;
    wire N__20532;
    wire N__20529;
    wire N__20526;
    wire N__20525;
    wire N__20522;
    wire N__20519;
    wire N__20518;
    wire N__20517;
    wire N__20516;
    wire N__20515;
    wire N__20514;
    wire N__20511;
    wire N__20510;
    wire N__20507;
    wire N__20504;
    wire N__20503;
    wire N__20500;
    wire N__20499;
    wire N__20496;
    wire N__20493;
    wire N__20492;
    wire N__20489;
    wire N__20488;
    wire N__20487;
    wire N__20486;
    wire N__20483;
    wire N__20480;
    wire N__20475;
    wire N__20472;
    wire N__20469;
    wire N__20466;
    wire N__20463;
    wire N__20460;
    wire N__20457;
    wire N__20454;
    wire N__20451;
    wire N__20448;
    wire N__20445;
    wire N__20440;
    wire N__20437;
    wire N__20434;
    wire N__20429;
    wire N__20426;
    wire N__20423;
    wire N__20420;
    wire N__20419;
    wire N__20414;
    wire N__20411;
    wire N__20408;
    wire N__20405;
    wire N__20400;
    wire N__20391;
    wire N__20388;
    wire N__20381;
    wire N__20370;
    wire N__20367;
    wire N__20364;
    wire N__20361;
    wire N__20358;
    wire N__20355;
    wire N__20352;
    wire N__20349;
    wire N__20346;
    wire N__20343;
    wire N__20340;
    wire N__20337;
    wire N__20334;
    wire N__20331;
    wire N__20328;
    wire N__20325;
    wire N__20322;
    wire N__20319;
    wire N__20316;
    wire N__20313;
    wire N__20310;
    wire N__20307;
    wire N__20304;
    wire N__20301;
    wire N__20298;
    wire N__20295;
    wire N__20292;
    wire N__20289;
    wire N__20286;
    wire N__20283;
    wire N__20280;
    wire N__20277;
    wire N__20274;
    wire N__20271;
    wire N__20268;
    wire N__20265;
    wire N__20262;
    wire N__20259;
    wire N__20256;
    wire N__20253;
    wire N__20250;
    wire N__20247;
    wire N__20244;
    wire N__20241;
    wire N__20238;
    wire N__20235;
    wire N__20232;
    wire N__20229;
    wire N__20226;
    wire N__20223;
    wire N__20220;
    wire N__20217;
    wire N__20214;
    wire N__20211;
    wire N__20208;
    wire N__20205;
    wire N__20202;
    wire N__20199;
    wire N__20196;
    wire N__20193;
    wire N__20190;
    wire N__20187;
    wire N__20184;
    wire N__20181;
    wire N__20178;
    wire N__20175;
    wire N__20172;
    wire N__20169;
    wire N__20168;
    wire N__20165;
    wire N__20162;
    wire N__20157;
    wire N__20154;
    wire N__20151;
    wire N__20148;
    wire N__20145;
    wire N__20142;
    wire N__20139;
    wire N__20138;
    wire N__20137;
    wire N__20136;
    wire N__20135;
    wire N__20134;
    wire N__20133;
    wire N__20132;
    wire N__20131;
    wire N__20130;
    wire N__20129;
    wire N__20126;
    wire N__20119;
    wire N__20112;
    wire N__20105;
    wire N__20104;
    wire N__20101;
    wire N__20100;
    wire N__20097;
    wire N__20096;
    wire N__20089;
    wire N__20086;
    wire N__20083;
    wire N__20080;
    wire N__20079;
    wire N__20076;
    wire N__20073;
    wire N__20068;
    wire N__20067;
    wire N__20066;
    wire N__20063;
    wire N__20060;
    wire N__20057;
    wire N__20056;
    wire N__20051;
    wire N__20048;
    wire N__20043;
    wire N__20036;
    wire N__20033;
    wire N__20022;
    wire N__20019;
    wire N__20018;
    wire N__20015;
    wire N__20012;
    wire N__20009;
    wire N__20006;
    wire N__20001;
    wire N__20000;
    wire N__19999;
    wire N__19996;
    wire N__19991;
    wire N__19988;
    wire N__19983;
    wire N__19980;
    wire N__19977;
    wire N__19974;
    wire N__19971;
    wire N__19968;
    wire N__19965;
    wire N__19962;
    wire N__19959;
    wire N__19956;
    wire N__19955;
    wire N__19952;
    wire N__19949;
    wire N__19946;
    wire N__19943;
    wire N__19940;
    wire N__19937;
    wire N__19934;
    wire N__19931;
    wire N__19926;
    wire N__19923;
    wire N__19922;
    wire N__19921;
    wire N__19918;
    wire N__19915;
    wire N__19914;
    wire N__19911;
    wire N__19910;
    wire N__19909;
    wire N__19904;
    wire N__19901;
    wire N__19898;
    wire N__19895;
    wire N__19892;
    wire N__19891;
    wire N__19888;
    wire N__19885;
    wire N__19878;
    wire N__19875;
    wire N__19874;
    wire N__19873;
    wire N__19870;
    wire N__19867;
    wire N__19862;
    wire N__19859;
    wire N__19856;
    wire N__19853;
    wire N__19850;
    wire N__19845;
    wire N__19842;
    wire N__19837;
    wire N__19834;
    wire N__19831;
    wire N__19826;
    wire N__19823;
    wire N__19818;
    wire N__19815;
    wire N__19812;
    wire N__19809;
    wire N__19806;
    wire N__19803;
    wire N__19800;
    wire N__19797;
    wire N__19794;
    wire N__19791;
    wire N__19788;
    wire N__19785;
    wire N__19782;
    wire N__19779;
    wire N__19776;
    wire N__19773;
    wire N__19770;
    wire N__19767;
    wire N__19764;
    wire N__19761;
    wire N__19758;
    wire N__19755;
    wire N__19752;
    wire N__19749;
    wire N__19746;
    wire N__19743;
    wire N__19740;
    wire N__19737;
    wire N__19734;
    wire N__19731;
    wire N__19728;
    wire N__19725;
    wire N__19722;
    wire N__19719;
    wire N__19716;
    wire N__19713;
    wire N__19710;
    wire N__19707;
    wire N__19704;
    wire N__19701;
    wire N__19698;
    wire N__19697;
    wire N__19694;
    wire N__19691;
    wire N__19690;
    wire N__19687;
    wire N__19686;
    wire N__19685;
    wire N__19684;
    wire N__19681;
    wire N__19680;
    wire N__19677;
    wire N__19676;
    wire N__19673;
    wire N__19672;
    wire N__19671;
    wire N__19670;
    wire N__19669;
    wire N__19668;
    wire N__19667;
    wire N__19664;
    wire N__19661;
    wire N__19660;
    wire N__19659;
    wire N__19656;
    wire N__19653;
    wire N__19650;
    wire N__19649;
    wire N__19646;
    wire N__19645;
    wire N__19642;
    wire N__19641;
    wire N__19638;
    wire N__19631;
    wire N__19626;
    wire N__19613;
    wire N__19608;
    wire N__19605;
    wire N__19602;
    wire N__19595;
    wire N__19594;
    wire N__19593;
    wire N__19592;
    wire N__19591;
    wire N__19586;
    wire N__19583;
    wire N__19576;
    wire N__19571;
    wire N__19568;
    wire N__19565;
    wire N__19560;
    wire N__19555;
    wire N__19542;
    wire N__19541;
    wire N__19538;
    wire N__19535;
    wire N__19532;
    wire N__19529;
    wire N__19526;
    wire N__19523;
    wire N__19520;
    wire N__19517;
    wire N__19514;
    wire N__19511;
    wire N__19508;
    wire N__19505;
    wire N__19502;
    wire N__19499;
    wire N__19496;
    wire N__19493;
    wire N__19490;
    wire N__19487;
    wire N__19484;
    wire N__19481;
    wire N__19478;
    wire N__19475;
    wire N__19472;
    wire N__19469;
    wire N__19466;
    wire N__19463;
    wire N__19460;
    wire N__19457;
    wire N__19454;
    wire N__19451;
    wire N__19448;
    wire N__19445;
    wire N__19442;
    wire N__19439;
    wire N__19436;
    wire N__19433;
    wire N__19430;
    wire N__19427;
    wire N__19424;
    wire N__19421;
    wire N__19418;
    wire N__19415;
    wire N__19412;
    wire N__19409;
    wire N__19406;
    wire N__19403;
    wire N__19400;
    wire N__19397;
    wire N__19394;
    wire N__19391;
    wire N__19388;
    wire N__19385;
    wire N__19382;
    wire N__19379;
    wire N__19376;
    wire N__19373;
    wire N__19370;
    wire N__19367;
    wire N__19364;
    wire N__19361;
    wire N__19358;
    wire N__19355;
    wire N__19352;
    wire N__19349;
    wire N__19348;
    wire N__19345;
    wire N__19342;
    wire N__19339;
    wire N__19336;
    wire N__19333;
    wire N__19330;
    wire N__19329;
    wire N__19326;
    wire N__19323;
    wire N__19320;
    wire N__19317;
    wire N__19314;
    wire N__19311;
    wire N__19302;
    wire N__19301;
    wire N__19300;
    wire N__19299;
    wire N__19298;
    wire N__19295;
    wire N__19292;
    wire N__19291;
    wire N__19288;
    wire N__19285;
    wire N__19282;
    wire N__19279;
    wire N__19276;
    wire N__19273;
    wire N__19272;
    wire N__19269;
    wire N__19266;
    wire N__19263;
    wire N__19260;
    wire N__19255;
    wire N__19252;
    wire N__19249;
    wire N__19246;
    wire N__19243;
    wire N__19236;
    wire N__19227;
    wire N__19224;
    wire N__19221;
    wire N__19218;
    wire N__19215;
    wire N__19212;
    wire N__19209;
    wire N__19206;
    wire N__19203;
    wire N__19200;
    wire N__19197;
    wire N__19194;
    wire N__19191;
    wire N__19190;
    wire N__19187;
    wire N__19184;
    wire N__19181;
    wire N__19180;
    wire N__19179;
    wire N__19174;
    wire N__19169;
    wire N__19164;
    wire N__19161;
    wire N__19158;
    wire N__19155;
    wire N__19152;
    wire N__19149;
    wire N__19148;
    wire N__19145;
    wire N__19142;
    wire N__19141;
    wire N__19140;
    wire N__19135;
    wire N__19134;
    wire N__19133;
    wire N__19130;
    wire N__19129;
    wire N__19126;
    wire N__19123;
    wire N__19120;
    wire N__19119;
    wire N__19116;
    wire N__19113;
    wire N__19110;
    wire N__19107;
    wire N__19102;
    wire N__19099;
    wire N__19096;
    wire N__19093;
    wire N__19090;
    wire N__19087;
    wire N__19082;
    wire N__19079;
    wire N__19074;
    wire N__19069;
    wire N__19064;
    wire N__19061;
    wire N__19056;
    wire N__19055;
    wire N__19052;
    wire N__19049;
    wire N__19044;
    wire N__19043;
    wire N__19040;
    wire N__19037;
    wire N__19032;
    wire N__19031;
    wire N__19028;
    wire N__19025;
    wire N__19020;
    wire N__19019;
    wire N__19016;
    wire N__19013;
    wire N__19008;
    wire N__19005;
    wire N__19002;
    wire N__18999;
    wire N__18998;
    wire N__18995;
    wire N__18992;
    wire N__18989;
    wire N__18984;
    wire N__18981;
    wire N__18978;
    wire N__18975;
    wire N__18972;
    wire N__18969;
    wire N__18966;
    wire N__18963;
    wire N__18960;
    wire N__18959;
    wire N__18956;
    wire N__18953;
    wire N__18948;
    wire N__18947;
    wire N__18944;
    wire N__18941;
    wire N__18938;
    wire N__18935;
    wire N__18930;
    wire N__18929;
    wire N__18926;
    wire N__18923;
    wire N__18922;
    wire N__18921;
    wire N__18920;
    wire N__18919;
    wire N__18918;
    wire N__18917;
    wire N__18916;
    wire N__18913;
    wire N__18910;
    wire N__18903;
    wire N__18900;
    wire N__18895;
    wire N__18892;
    wire N__18889;
    wire N__18884;
    wire N__18873;
    wire N__18872;
    wire N__18871;
    wire N__18868;
    wire N__18867;
    wire N__18866;
    wire N__18863;
    wire N__18860;
    wire N__18857;
    wire N__18854;
    wire N__18851;
    wire N__18850;
    wire N__18849;
    wire N__18846;
    wire N__18843;
    wire N__18840;
    wire N__18835;
    wire N__18834;
    wire N__18833;
    wire N__18830;
    wire N__18827;
    wire N__18824;
    wire N__18817;
    wire N__18814;
    wire N__18809;
    wire N__18806;
    wire N__18803;
    wire N__18800;
    wire N__18789;
    wire N__18788;
    wire N__18785;
    wire N__18782;
    wire N__18781;
    wire N__18780;
    wire N__18779;
    wire N__18778;
    wire N__18777;
    wire N__18776;
    wire N__18773;
    wire N__18770;
    wire N__18763;
    wire N__18762;
    wire N__18759;
    wire N__18754;
    wire N__18751;
    wire N__18748;
    wire N__18745;
    wire N__18742;
    wire N__18729;
    wire N__18726;
    wire N__18725;
    wire N__18722;
    wire N__18719;
    wire N__18718;
    wire N__18717;
    wire N__18712;
    wire N__18709;
    wire N__18706;
    wire N__18699;
    wire N__18696;
    wire N__18693;
    wire N__18690;
    wire N__18687;
    wire N__18686;
    wire N__18683;
    wire N__18680;
    wire N__18675;
    wire N__18672;
    wire N__18669;
    wire N__18666;
    wire N__18663;
    wire N__18662;
    wire N__18659;
    wire N__18656;
    wire N__18655;
    wire N__18652;
    wire N__18649;
    wire N__18646;
    wire N__18645;
    wire N__18642;
    wire N__18639;
    wire N__18636;
    wire N__18633;
    wire N__18624;
    wire N__18623;
    wire N__18622;
    wire N__18621;
    wire N__18618;
    wire N__18613;
    wire N__18610;
    wire N__18603;
    wire N__18600;
    wire N__18599;
    wire N__18596;
    wire N__18595;
    wire N__18594;
    wire N__18591;
    wire N__18588;
    wire N__18583;
    wire N__18576;
    wire N__18573;
    wire N__18572;
    wire N__18571;
    wire N__18570;
    wire N__18567;
    wire N__18562;
    wire N__18559;
    wire N__18552;
    wire N__18549;
    wire N__18546;
    wire N__18545;
    wire N__18544;
    wire N__18543;
    wire N__18540;
    wire N__18537;
    wire N__18532;
    wire N__18525;
    wire N__18522;
    wire N__18521;
    wire N__18520;
    wire N__18519;
    wire N__18516;
    wire N__18509;
    wire N__18504;
    wire N__18501;
    wire N__18500;
    wire N__18499;
    wire N__18496;
    wire N__18491;
    wire N__18486;
    wire N__18483;
    wire N__18482;
    wire N__18481;
    wire N__18478;
    wire N__18475;
    wire N__18472;
    wire N__18465;
    wire N__18462;
    wire N__18461;
    wire N__18460;
    wire N__18459;
    wire N__18456;
    wire N__18451;
    wire N__18448;
    wire N__18441;
    wire N__18438;
    wire N__18435;
    wire N__18432;
    wire N__18429;
    wire N__18426;
    wire N__18423;
    wire N__18420;
    wire N__18417;
    wire N__18414;
    wire N__18411;
    wire N__18408;
    wire N__18405;
    wire N__18402;
    wire N__18399;
    wire N__18396;
    wire N__18393;
    wire N__18390;
    wire N__18387;
    wire N__18384;
    wire N__18381;
    wire N__18378;
    wire N__18375;
    wire N__18372;
    wire N__18369;
    wire N__18366;
    wire N__18363;
    wire N__18360;
    wire N__18357;
    wire N__18354;
    wire N__18351;
    wire N__18348;
    wire N__18345;
    wire N__18342;
    wire N__18339;
    wire N__18338;
    wire N__18337;
    wire N__18334;
    wire N__18331;
    wire N__18328;
    wire N__18325;
    wire N__18322;
    wire N__18319;
    wire N__18316;
    wire N__18313;
    wire N__18310;
    wire N__18307;
    wire N__18304;
    wire N__18301;
    wire N__18298;
    wire N__18295;
    wire N__18292;
    wire N__18289;
    wire N__18286;
    wire N__18283;
    wire N__18276;
    wire N__18275;
    wire N__18272;
    wire N__18271;
    wire N__18270;
    wire N__18267;
    wire N__18264;
    wire N__18261;
    wire N__18258;
    wire N__18255;
    wire N__18248;
    wire N__18245;
    wire N__18242;
    wire N__18239;
    wire N__18236;
    wire N__18233;
    wire N__18230;
    wire N__18225;
    wire N__18222;
    wire N__18219;
    wire N__18216;
    wire N__18215;
    wire N__18212;
    wire N__18209;
    wire N__18206;
    wire N__18203;
    wire N__18200;
    wire N__18197;
    wire N__18194;
    wire N__18191;
    wire N__18186;
    wire N__18183;
    wire N__18180;
    wire N__18177;
    wire N__18176;
    wire N__18173;
    wire N__18170;
    wire N__18167;
    wire N__18164;
    wire N__18163;
    wire N__18160;
    wire N__18157;
    wire N__18154;
    wire N__18147;
    wire N__18144;
    wire N__18141;
    wire N__18138;
    wire N__18135;
    wire N__18132;
    wire N__18129;
    wire N__18126;
    wire N__18123;
    wire N__18120;
    wire N__18117;
    wire N__18114;
    wire N__18111;
    wire N__18108;
    wire N__18105;
    wire N__18104;
    wire N__18101;
    wire N__18098;
    wire N__18097;
    wire N__18092;
    wire N__18091;
    wire N__18088;
    wire N__18085;
    wire N__18082;
    wire N__18075;
    wire N__18072;
    wire N__18069;
    wire N__18066;
    wire N__18063;
    wire N__18060;
    wire N__18059;
    wire N__18056;
    wire N__18053;
    wire N__18050;
    wire N__18047;
    wire N__18044;
    wire N__18041;
    wire N__18038;
    wire N__18035;
    wire N__18032;
    wire N__18029;
    wire N__18026;
    wire N__18023;
    wire N__18020;
    wire N__18017;
    wire N__18014;
    wire N__18011;
    wire N__18008;
    wire N__18005;
    wire N__18002;
    wire N__17999;
    wire N__17996;
    wire N__17993;
    wire N__17990;
    wire N__17987;
    wire N__17984;
    wire N__17981;
    wire N__17978;
    wire N__17975;
    wire N__17972;
    wire N__17969;
    wire N__17966;
    wire N__17963;
    wire N__17960;
    wire N__17957;
    wire N__17954;
    wire N__17951;
    wire N__17948;
    wire N__17945;
    wire N__17942;
    wire N__17939;
    wire N__17936;
    wire N__17933;
    wire N__17930;
    wire N__17927;
    wire N__17924;
    wire N__17921;
    wire N__17918;
    wire N__17915;
    wire N__17912;
    wire N__17909;
    wire N__17906;
    wire N__17903;
    wire N__17900;
    wire N__17897;
    wire N__17894;
    wire N__17891;
    wire N__17888;
    wire N__17885;
    wire N__17882;
    wire N__17879;
    wire N__17876;
    wire N__17873;
    wire N__17870;
    wire N__17867;
    wire N__17864;
    wire N__17861;
    wire N__17858;
    wire N__17855;
    wire N__17854;
    wire N__17853;
    wire N__17850;
    wire N__17847;
    wire N__17844;
    wire N__17841;
    wire N__17838;
    wire N__17835;
    wire N__17832;
    wire N__17829;
    wire N__17824;
    wire N__17817;
    wire N__17814;
    wire N__17811;
    wire N__17808;
    wire N__17805;
    wire N__17804;
    wire N__17801;
    wire N__17798;
    wire N__17795;
    wire N__17792;
    wire N__17789;
    wire N__17786;
    wire N__17783;
    wire N__17780;
    wire N__17777;
    wire N__17774;
    wire N__17771;
    wire N__17768;
    wire N__17765;
    wire N__17762;
    wire N__17759;
    wire N__17756;
    wire N__17753;
    wire N__17750;
    wire N__17747;
    wire N__17744;
    wire N__17741;
    wire N__17738;
    wire N__17735;
    wire N__17732;
    wire N__17729;
    wire N__17726;
    wire N__17723;
    wire N__17720;
    wire N__17717;
    wire N__17714;
    wire N__17711;
    wire N__17708;
    wire N__17705;
    wire N__17702;
    wire N__17699;
    wire N__17696;
    wire N__17693;
    wire N__17690;
    wire N__17687;
    wire N__17684;
    wire N__17681;
    wire N__17678;
    wire N__17675;
    wire N__17672;
    wire N__17669;
    wire N__17666;
    wire N__17663;
    wire N__17660;
    wire N__17657;
    wire N__17654;
    wire N__17651;
    wire N__17648;
    wire N__17645;
    wire N__17642;
    wire N__17639;
    wire N__17636;
    wire N__17633;
    wire N__17630;
    wire N__17627;
    wire N__17624;
    wire N__17621;
    wire N__17618;
    wire N__17617;
    wire N__17614;
    wire N__17611;
    wire N__17608;
    wire N__17605;
    wire N__17602;
    wire N__17599;
    wire N__17598;
    wire N__17595;
    wire N__17592;
    wire N__17589;
    wire N__17586;
    wire N__17583;
    wire N__17580;
    wire N__17571;
    wire N__17568;
    wire N__17565;
    wire N__17562;
    wire N__17561;
    wire N__17558;
    wire N__17555;
    wire N__17552;
    wire N__17549;
    wire N__17546;
    wire N__17543;
    wire N__17540;
    wire N__17537;
    wire N__17534;
    wire N__17531;
    wire N__17528;
    wire N__17525;
    wire N__17522;
    wire N__17519;
    wire N__17516;
    wire N__17513;
    wire N__17510;
    wire N__17507;
    wire N__17504;
    wire N__17501;
    wire N__17498;
    wire N__17495;
    wire N__17492;
    wire N__17489;
    wire N__17486;
    wire N__17483;
    wire N__17480;
    wire N__17477;
    wire N__17474;
    wire N__17471;
    wire N__17468;
    wire N__17465;
    wire N__17462;
    wire N__17459;
    wire N__17456;
    wire N__17453;
    wire N__17450;
    wire N__17447;
    wire N__17444;
    wire N__17441;
    wire N__17438;
    wire N__17435;
    wire N__17432;
    wire N__17429;
    wire N__17426;
    wire N__17423;
    wire N__17420;
    wire N__17417;
    wire N__17414;
    wire N__17411;
    wire N__17408;
    wire N__17405;
    wire N__17402;
    wire N__17399;
    wire N__17396;
    wire N__17393;
    wire N__17390;
    wire N__17387;
    wire N__17384;
    wire N__17381;
    wire N__17378;
    wire N__17375;
    wire N__17372;
    wire N__17369;
    wire N__17366;
    wire N__17363;
    wire N__17362;
    wire N__17361;
    wire N__17358;
    wire N__17355;
    wire N__17352;
    wire N__17349;
    wire N__17346;
    wire N__17343;
    wire N__17340;
    wire N__17337;
    wire N__17332;
    wire N__17329;
    wire N__17324;
    wire N__17319;
    wire N__17316;
    wire N__17313;
    wire N__17310;
    wire N__17309;
    wire N__17306;
    wire N__17303;
    wire N__17300;
    wire N__17297;
    wire N__17294;
    wire N__17291;
    wire N__17288;
    wire N__17285;
    wire N__17282;
    wire N__17279;
    wire N__17276;
    wire N__17273;
    wire N__17270;
    wire N__17267;
    wire N__17264;
    wire N__17261;
    wire N__17258;
    wire N__17255;
    wire N__17252;
    wire N__17249;
    wire N__17246;
    wire N__17243;
    wire N__17240;
    wire N__17237;
    wire N__17234;
    wire N__17231;
    wire N__17228;
    wire N__17225;
    wire N__17222;
    wire N__17219;
    wire N__17216;
    wire N__17213;
    wire N__17210;
    wire N__17207;
    wire N__17204;
    wire N__17201;
    wire N__17198;
    wire N__17195;
    wire N__17192;
    wire N__17189;
    wire N__17186;
    wire N__17183;
    wire N__17180;
    wire N__17177;
    wire N__17174;
    wire N__17171;
    wire N__17168;
    wire N__17165;
    wire N__17162;
    wire N__17159;
    wire N__17156;
    wire N__17153;
    wire N__17150;
    wire N__17147;
    wire N__17144;
    wire N__17141;
    wire N__17138;
    wire N__17135;
    wire N__17132;
    wire N__17129;
    wire N__17126;
    wire N__17123;
    wire N__17120;
    wire N__17117;
    wire N__17116;
    wire N__17113;
    wire N__17110;
    wire N__17107;
    wire N__17104;
    wire N__17101;
    wire N__17100;
    wire N__17097;
    wire N__17094;
    wire N__17091;
    wire N__17088;
    wire N__17083;
    wire N__17080;
    wire N__17073;
    wire N__17070;
    wire N__17067;
    wire N__17064;
    wire N__17061;
    wire N__17060;
    wire N__17057;
    wire N__17054;
    wire N__17051;
    wire N__17048;
    wire N__17045;
    wire N__17042;
    wire N__17039;
    wire N__17036;
    wire N__17033;
    wire N__17030;
    wire N__17027;
    wire N__17024;
    wire N__17021;
    wire N__17018;
    wire N__17015;
    wire N__17012;
    wire N__17009;
    wire N__17006;
    wire N__17003;
    wire N__17000;
    wire N__16997;
    wire N__16994;
    wire N__16991;
    wire N__16988;
    wire N__16985;
    wire N__16982;
    wire N__16979;
    wire N__16976;
    wire N__16973;
    wire N__16970;
    wire N__16967;
    wire N__16964;
    wire N__16961;
    wire N__16958;
    wire N__16955;
    wire N__16952;
    wire N__16949;
    wire N__16946;
    wire N__16943;
    wire N__16940;
    wire N__16937;
    wire N__16934;
    wire N__16931;
    wire N__16928;
    wire N__16925;
    wire N__16922;
    wire N__16919;
    wire N__16916;
    wire N__16913;
    wire N__16910;
    wire N__16907;
    wire N__16904;
    wire N__16901;
    wire N__16898;
    wire N__16895;
    wire N__16892;
    wire N__16889;
    wire N__16886;
    wire N__16883;
    wire N__16880;
    wire N__16877;
    wire N__16874;
    wire N__16871;
    wire N__16868;
    wire N__16865;
    wire N__16864;
    wire N__16861;
    wire N__16858;
    wire N__16857;
    wire N__16854;
    wire N__16851;
    wire N__16848;
    wire N__16845;
    wire N__16842;
    wire N__16839;
    wire N__16836;
    wire N__16833;
    wire N__16830;
    wire N__16825;
    wire N__16818;
    wire N__16815;
    wire N__16812;
    wire N__16809;
    wire N__16808;
    wire N__16805;
    wire N__16802;
    wire N__16799;
    wire N__16796;
    wire N__16793;
    wire N__16790;
    wire N__16787;
    wire N__16784;
    wire N__16781;
    wire N__16778;
    wire N__16775;
    wire N__16772;
    wire N__16769;
    wire N__16766;
    wire N__16763;
    wire N__16760;
    wire N__16757;
    wire N__16754;
    wire N__16751;
    wire N__16748;
    wire N__16745;
    wire N__16742;
    wire N__16739;
    wire N__16736;
    wire N__16733;
    wire N__16730;
    wire N__16727;
    wire N__16724;
    wire N__16721;
    wire N__16718;
    wire N__16715;
    wire N__16712;
    wire N__16709;
    wire N__16706;
    wire N__16703;
    wire N__16700;
    wire N__16697;
    wire N__16694;
    wire N__16691;
    wire N__16688;
    wire N__16685;
    wire N__16682;
    wire N__16679;
    wire N__16676;
    wire N__16673;
    wire N__16670;
    wire N__16667;
    wire N__16664;
    wire N__16661;
    wire N__16658;
    wire N__16655;
    wire N__16652;
    wire N__16649;
    wire N__16646;
    wire N__16643;
    wire N__16640;
    wire N__16637;
    wire N__16634;
    wire N__16631;
    wire N__16628;
    wire N__16625;
    wire N__16622;
    wire N__16619;
    wire N__16618;
    wire N__16615;
    wire N__16612;
    wire N__16609;
    wire N__16606;
    wire N__16603;
    wire N__16600;
    wire N__16599;
    wire N__16596;
    wire N__16593;
    wire N__16590;
    wire N__16587;
    wire N__16584;
    wire N__16581;
    wire N__16572;
    wire N__16569;
    wire N__16566;
    wire N__16563;
    wire N__16560;
    wire N__16557;
    wire N__16554;
    wire N__16551;
    wire N__16548;
    wire N__16545;
    wire N__16542;
    wire N__16539;
    wire N__16536;
    wire N__16533;
    wire N__16532;
    wire N__16529;
    wire N__16528;
    wire N__16527;
    wire N__16524;
    wire N__16521;
    wire N__16518;
    wire N__16515;
    wire N__16512;
    wire N__16509;
    wire N__16506;
    wire N__16503;
    wire N__16500;
    wire N__16497;
    wire N__16492;
    wire N__16489;
    wire N__16486;
    wire N__16481;
    wire N__16476;
    wire N__16473;
    wire N__16470;
    wire N__16467;
    wire N__16466;
    wire N__16465;
    wire N__16464;
    wire N__16461;
    wire N__16458;
    wire N__16455;
    wire N__16452;
    wire N__16447;
    wire N__16442;
    wire N__16437;
    wire N__16434;
    wire N__16431;
    wire N__16428;
    wire N__16427;
    wire N__16424;
    wire N__16423;
    wire N__16420;
    wire N__16417;
    wire N__16414;
    wire N__16413;
    wire N__16410;
    wire N__16405;
    wire N__16402;
    wire N__16399;
    wire N__16394;
    wire N__16391;
    wire N__16388;
    wire N__16385;
    wire N__16382;
    wire N__16377;
    wire N__16374;
    wire N__16371;
    wire N__16368;
    wire N__16365;
    wire N__16362;
    wire N__16359;
    wire N__16356;
    wire N__16353;
    wire N__16350;
    wire N__16347;
    wire N__16344;
    wire N__16341;
    wire N__16338;
    wire N__16335;
    wire N__16332;
    wire N__16329;
    wire N__16326;
    wire N__16323;
    wire N__16322;
    wire N__16321;
    wire N__16320;
    wire N__16319;
    wire N__16318;
    wire N__16317;
    wire N__16316;
    wire N__16315;
    wire N__16314;
    wire N__16309;
    wire N__16308;
    wire N__16307;
    wire N__16306;
    wire N__16305;
    wire N__16304;
    wire N__16301;
    wire N__16300;
    wire N__16299;
    wire N__16298;
    wire N__16291;
    wire N__16282;
    wire N__16279;
    wire N__16276;
    wire N__16267;
    wire N__16266;
    wire N__16265;
    wire N__16264;
    wire N__16261;
    wire N__16254;
    wire N__16251;
    wire N__16242;
    wire N__16241;
    wire N__16240;
    wire N__16239;
    wire N__16238;
    wire N__16237;
    wire N__16234;
    wire N__16233;
    wire N__16230;
    wire N__16227;
    wire N__16222;
    wire N__16217;
    wire N__16210;
    wire N__16201;
    wire N__16188;
    wire N__16185;
    wire N__16182;
    wire N__16179;
    wire N__16176;
    wire N__16173;
    wire N__16170;
    wire N__16167;
    wire N__16164;
    wire N__16161;
    wire N__16158;
    wire N__16155;
    wire N__16152;
    wire N__16149;
    wire N__16148;
    wire N__16145;
    wire N__16142;
    wire N__16141;
    wire N__16140;
    wire N__16135;
    wire N__16132;
    wire N__16129;
    wire N__16124;
    wire N__16121;
    wire N__16118;
    wire N__16115;
    wire N__16112;
    wire N__16107;
    wire N__16104;
    wire N__16103;
    wire N__16100;
    wire N__16097;
    wire N__16096;
    wire N__16091;
    wire N__16088;
    wire N__16087;
    wire N__16082;
    wire N__16079;
    wire N__16076;
    wire N__16073;
    wire N__16070;
    wire N__16067;
    wire N__16064;
    wire N__16061;
    wire N__16058;
    wire N__16055;
    wire N__16050;
    wire N__16047;
    wire N__16044;
    wire N__16041;
    wire N__16038;
    wire N__16035;
    wire N__16032;
    wire N__16031;
    wire N__16028;
    wire N__16025;
    wire N__16020;
    wire N__16019;
    wire N__16016;
    wire N__16013;
    wire N__16008;
    wire N__16005;
    wire N__16004;
    wire N__16003;
    wire N__16000;
    wire N__15997;
    wire N__15994;
    wire N__15991;
    wire N__15988;
    wire N__15981;
    wire N__15978;
    wire N__15977;
    wire N__15976;
    wire N__15973;
    wire N__15970;
    wire N__15967;
    wire N__15964;
    wire N__15961;
    wire N__15954;
    wire N__15951;
    wire N__15950;
    wire N__15947;
    wire N__15946;
    wire N__15943;
    wire N__15940;
    wire N__15937;
    wire N__15934;
    wire N__15931;
    wire N__15924;
    wire N__15923;
    wire N__15920;
    wire N__15917;
    wire N__15912;
    wire N__15909;
    wire N__15908;
    wire N__15905;
    wire N__15902;
    wire N__15901;
    wire N__15898;
    wire N__15895;
    wire N__15892;
    wire N__15889;
    wire N__15886;
    wire N__15879;
    wire N__15876;
    wire N__15873;
    wire N__15872;
    wire N__15871;
    wire N__15868;
    wire N__15865;
    wire N__15862;
    wire N__15859;
    wire N__15856;
    wire N__15849;
    wire N__15848;
    wire N__15843;
    wire N__15842;
    wire N__15839;
    wire N__15836;
    wire N__15833;
    wire N__15828;
    wire N__15825;
    wire N__15824;
    wire N__15821;
    wire N__15818;
    wire N__15815;
    wire N__15810;
    wire N__15807;
    wire N__15804;
    wire N__15801;
    wire N__15798;
    wire N__15795;
    wire N__15792;
    wire N__15789;
    wire N__15786;
    wire N__15783;
    wire N__15780;
    wire N__15777;
    wire N__15774;
    wire N__15771;
    wire N__15768;
    wire N__15765;
    wire N__15762;
    wire N__15761;
    wire N__15758;
    wire N__15755;
    wire N__15750;
    wire N__15747;
    wire N__15746;
    wire N__15743;
    wire N__15740;
    wire N__15737;
    wire N__15734;
    wire N__15729;
    wire N__15728;
    wire N__15725;
    wire N__15722;
    wire N__15717;
    wire N__15716;
    wire N__15713;
    wire N__15710;
    wire N__15705;
    wire N__15704;
    wire N__15701;
    wire N__15698;
    wire N__15693;
    wire N__15690;
    wire N__15687;
    wire N__15684;
    wire N__15681;
    wire N__15678;
    wire N__15675;
    wire N__15672;
    wire N__15669;
    wire N__15666;
    wire N__15663;
    wire N__15660;
    wire N__15657;
    wire N__15654;
    wire N__15653;
    wire N__15650;
    wire N__15647;
    wire N__15644;
    wire N__15641;
    wire N__15640;
    wire N__15637;
    wire N__15636;
    wire N__15635;
    wire N__15632;
    wire N__15631;
    wire N__15628;
    wire N__15625;
    wire N__15622;
    wire N__15619;
    wire N__15616;
    wire N__15613;
    wire N__15610;
    wire N__15605;
    wire N__15602;
    wire N__15597;
    wire N__15594;
    wire N__15593;
    wire N__15590;
    wire N__15587;
    wire N__15586;
    wire N__15583;
    wire N__15580;
    wire N__15577;
    wire N__15572;
    wire N__15569;
    wire N__15562;
    wire N__15557;
    wire N__15552;
    wire N__15549;
    wire N__15546;
    wire N__15543;
    wire N__15540;
    wire N__15537;
    wire N__15534;
    wire N__15531;
    wire N__15528;
    wire N__15525;
    wire N__15524;
    wire N__15521;
    wire N__15518;
    wire N__15515;
    wire N__15514;
    wire N__15513;
    wire N__15508;
    wire N__15505;
    wire N__15502;
    wire N__15495;
    wire N__15492;
    wire N__15489;
    wire N__15488;
    wire N__15487;
    wire N__15484;
    wire N__15481;
    wire N__15478;
    wire N__15477;
    wire N__15474;
    wire N__15469;
    wire N__15466;
    wire N__15463;
    wire N__15460;
    wire N__15457;
    wire N__15450;
    wire N__15447;
    wire N__15444;
    wire N__15443;
    wire N__15440;
    wire N__15439;
    wire N__15436;
    wire N__15433;
    wire N__15432;
    wire N__15429;
    wire N__15426;
    wire N__15423;
    wire N__15420;
    wire N__15417;
    wire N__15408;
    wire N__15405;
    wire N__15402;
    wire N__15401;
    wire N__15398;
    wire N__15397;
    wire N__15394;
    wire N__15391;
    wire N__15390;
    wire N__15389;
    wire N__15388;
    wire N__15385;
    wire N__15382;
    wire N__15379;
    wire N__15376;
    wire N__15373;
    wire N__15370;
    wire N__15367;
    wire N__15364;
    wire N__15361;
    wire N__15358;
    wire N__15355;
    wire N__15350;
    wire N__15345;
    wire N__15342;
    wire N__15339;
    wire N__15336;
    wire N__15327;
    wire N__15324;
    wire N__15321;
    wire N__15318;
    wire N__15317;
    wire N__15314;
    wire N__15311;
    wire N__15308;
    wire N__15305;
    wire N__15302;
    wire N__15299;
    wire N__15296;
    wire N__15293;
    wire N__15290;
    wire N__15287;
    wire N__15284;
    wire N__15281;
    wire N__15278;
    wire N__15275;
    wire N__15272;
    wire N__15269;
    wire N__15266;
    wire N__15263;
    wire N__15260;
    wire N__15257;
    wire N__15254;
    wire N__15251;
    wire N__15248;
    wire N__15245;
    wire N__15242;
    wire N__15239;
    wire N__15236;
    wire N__15233;
    wire N__15230;
    wire N__15227;
    wire N__15224;
    wire N__15221;
    wire N__15218;
    wire N__15215;
    wire N__15212;
    wire N__15209;
    wire N__15206;
    wire N__15203;
    wire N__15200;
    wire N__15197;
    wire N__15194;
    wire N__15191;
    wire N__15188;
    wire N__15185;
    wire N__15182;
    wire N__15179;
    wire N__15176;
    wire N__15173;
    wire N__15170;
    wire N__15167;
    wire N__15164;
    wire N__15161;
    wire N__15158;
    wire N__15155;
    wire N__15152;
    wire N__15149;
    wire N__15146;
    wire N__15143;
    wire N__15140;
    wire N__15137;
    wire N__15134;
    wire N__15131;
    wire N__15128;
    wire N__15125;
    wire N__15124;
    wire N__15123;
    wire N__15120;
    wire N__15117;
    wire N__15114;
    wire N__15111;
    wire N__15106;
    wire N__15103;
    wire N__15100;
    wire N__15097;
    wire N__15090;
    wire N__15087;
    wire N__15084;
    wire N__15081;
    wire N__15080;
    wire N__15077;
    wire N__15074;
    wire N__15071;
    wire N__15068;
    wire N__15065;
    wire N__15062;
    wire N__15059;
    wire N__15056;
    wire N__15053;
    wire N__15050;
    wire N__15047;
    wire N__15044;
    wire N__15041;
    wire N__15038;
    wire N__15035;
    wire N__15032;
    wire N__15029;
    wire N__15026;
    wire N__15023;
    wire N__15020;
    wire N__15017;
    wire N__15014;
    wire N__15011;
    wire N__15008;
    wire N__15005;
    wire N__15002;
    wire N__14999;
    wire N__14996;
    wire N__14993;
    wire N__14990;
    wire N__14987;
    wire N__14984;
    wire N__14981;
    wire N__14978;
    wire N__14975;
    wire N__14972;
    wire N__14969;
    wire N__14966;
    wire N__14963;
    wire N__14960;
    wire N__14957;
    wire N__14954;
    wire N__14951;
    wire N__14948;
    wire N__14945;
    wire N__14942;
    wire N__14939;
    wire N__14936;
    wire N__14933;
    wire N__14930;
    wire N__14927;
    wire N__14924;
    wire N__14921;
    wire N__14918;
    wire N__14915;
    wire N__14912;
    wire N__14909;
    wire N__14906;
    wire N__14903;
    wire N__14900;
    wire N__14897;
    wire N__14894;
    wire N__14891;
    wire N__14888;
    wire N__14885;
    wire N__14882;
    wire N__14881;
    wire N__14880;
    wire N__14877;
    wire N__14874;
    wire N__14871;
    wire N__14868;
    wire N__14865;
    wire N__14862;
    wire N__14859;
    wire N__14856;
    wire N__14851;
    wire N__14844;
    wire N__14841;
    wire N__14838;
    wire N__14835;
    wire N__14834;
    wire N__14831;
    wire N__14828;
    wire N__14825;
    wire N__14822;
    wire N__14819;
    wire N__14816;
    wire N__14813;
    wire N__14810;
    wire N__14807;
    wire N__14804;
    wire N__14801;
    wire N__14798;
    wire N__14795;
    wire N__14792;
    wire N__14789;
    wire N__14786;
    wire N__14783;
    wire N__14780;
    wire N__14777;
    wire N__14774;
    wire N__14771;
    wire N__14768;
    wire N__14765;
    wire N__14762;
    wire N__14759;
    wire N__14756;
    wire N__14753;
    wire N__14750;
    wire N__14747;
    wire N__14744;
    wire N__14741;
    wire N__14738;
    wire N__14735;
    wire N__14732;
    wire N__14729;
    wire N__14726;
    wire N__14723;
    wire N__14720;
    wire N__14717;
    wire N__14714;
    wire N__14711;
    wire N__14708;
    wire N__14705;
    wire N__14702;
    wire N__14699;
    wire N__14696;
    wire N__14693;
    wire N__14690;
    wire N__14687;
    wire N__14684;
    wire N__14681;
    wire N__14678;
    wire N__14675;
    wire N__14672;
    wire N__14669;
    wire N__14666;
    wire N__14663;
    wire N__14660;
    wire N__14657;
    wire N__14654;
    wire N__14651;
    wire N__14648;
    wire N__14645;
    wire N__14642;
    wire N__14639;
    wire N__14638;
    wire N__14637;
    wire N__14634;
    wire N__14631;
    wire N__14628;
    wire N__14625;
    wire N__14622;
    wire N__14619;
    wire N__14616;
    wire N__14613;
    wire N__14610;
    wire N__14607;
    wire N__14598;
    wire N__14597;
    wire N__14594;
    wire N__14593;
    wire N__14590;
    wire N__14587;
    wire N__14584;
    wire N__14581;
    wire N__14578;
    wire N__14575;
    wire N__14570;
    wire N__14567;
    wire N__14564;
    wire N__14561;
    wire N__14556;
    wire N__14553;
    wire N__14550;
    wire N__14547;
    wire N__14544;
    wire N__14541;
    wire N__14538;
    wire N__14537;
    wire N__14534;
    wire N__14531;
    wire N__14528;
    wire N__14525;
    wire N__14522;
    wire N__14519;
    wire N__14516;
    wire N__14513;
    wire N__14510;
    wire N__14507;
    wire N__14504;
    wire N__14501;
    wire N__14498;
    wire N__14495;
    wire N__14492;
    wire N__14489;
    wire N__14486;
    wire N__14483;
    wire N__14480;
    wire N__14477;
    wire N__14474;
    wire N__14471;
    wire N__14468;
    wire N__14465;
    wire N__14462;
    wire N__14459;
    wire N__14456;
    wire N__14453;
    wire N__14450;
    wire N__14447;
    wire N__14444;
    wire N__14441;
    wire N__14438;
    wire N__14435;
    wire N__14432;
    wire N__14429;
    wire N__14426;
    wire N__14423;
    wire N__14420;
    wire N__14417;
    wire N__14414;
    wire N__14411;
    wire N__14408;
    wire N__14405;
    wire N__14402;
    wire N__14399;
    wire N__14396;
    wire N__14393;
    wire N__14390;
    wire N__14387;
    wire N__14384;
    wire N__14381;
    wire N__14378;
    wire N__14375;
    wire N__14372;
    wire N__14369;
    wire N__14366;
    wire N__14363;
    wire N__14360;
    wire N__14357;
    wire N__14356;
    wire N__14353;
    wire N__14350;
    wire N__14347;
    wire N__14344;
    wire N__14341;
    wire N__14338;
    wire N__14335;
    wire N__14332;
    wire N__14329;
    wire N__14328;
    wire N__14325;
    wire N__14322;
    wire N__14319;
    wire N__14316;
    wire N__14313;
    wire N__14310;
    wire N__14301;
    wire N__14298;
    wire N__14295;
    wire N__14292;
    wire N__14289;
    wire N__14286;
    wire N__14283;
    wire N__14280;
    wire N__14277;
    wire N__14274;
    wire N__14271;
    wire N__14268;
    wire N__14265;
    wire N__14262;
    wire N__14259;
    wire N__14258;
    wire N__14255;
    wire N__14252;
    wire N__14249;
    wire N__14246;
    wire N__14243;
    wire N__14240;
    wire N__14237;
    wire N__14234;
    wire N__14231;
    wire N__14228;
    wire N__14225;
    wire N__14222;
    wire N__14219;
    wire N__14216;
    wire N__14213;
    wire N__14210;
    wire N__14207;
    wire N__14204;
    wire N__14201;
    wire N__14198;
    wire N__14195;
    wire N__14192;
    wire N__14189;
    wire N__14186;
    wire N__14183;
    wire N__14180;
    wire N__14177;
    wire N__14174;
    wire N__14171;
    wire N__14168;
    wire N__14165;
    wire N__14162;
    wire N__14159;
    wire N__14156;
    wire N__14153;
    wire N__14150;
    wire N__14147;
    wire N__14144;
    wire N__14141;
    wire N__14138;
    wire N__14135;
    wire N__14132;
    wire N__14129;
    wire N__14126;
    wire N__14123;
    wire N__14120;
    wire N__14117;
    wire N__14114;
    wire N__14111;
    wire N__14108;
    wire N__14105;
    wire N__14102;
    wire N__14099;
    wire N__14096;
    wire N__14093;
    wire N__14090;
    wire N__14087;
    wire N__14084;
    wire N__14081;
    wire N__14078;
    wire N__14075;
    wire N__14072;
    wire N__14069;
    wire N__14066;
    wire N__14063;
    wire N__14060;
    wire N__14057;
    wire N__14054;
    wire N__14051;
    wire N__14048;
    wire N__14043;
    wire N__14042;
    wire N__14041;
    wire N__14040;
    wire N__14039;
    wire N__14036;
    wire N__14033;
    wire N__14030;
    wire N__14029;
    wire N__14028;
    wire N__14027;
    wire N__14026;
    wire N__14025;
    wire N__14024;
    wire N__14021;
    wire N__14018;
    wire N__14011;
    wire N__14006;
    wire N__14003;
    wire N__14002;
    wire N__14001;
    wire N__14000;
    wire N__13995;
    wire N__13992;
    wire N__13987;
    wire N__13980;
    wire N__13973;
    wire N__13962;
    wire N__13959;
    wire N__13956;
    wire N__13953;
    wire N__13950;
    wire N__13947;
    wire N__13944;
    wire N__13941;
    wire N__13938;
    wire N__13935;
    wire N__13932;
    wire N__13929;
    wire N__13928;
    wire N__13923;
    wire N__13920;
    wire N__13917;
    wire N__13914;
    wire N__13913;
    wire N__13910;
    wire N__13909;
    wire N__13908;
    wire N__13905;
    wire N__13902;
    wire N__13899;
    wire N__13896;
    wire N__13893;
    wire N__13884;
    wire N__13881;
    wire N__13878;
    wire N__13875;
    wire N__13872;
    wire N__13869;
    wire N__13866;
    wire N__13863;
    wire N__13860;
    wire N__13857;
    wire N__13854;
    wire N__13851;
    wire N__13848;
    wire N__13845;
    wire N__13842;
    wire N__13839;
    wire N__13836;
    wire N__13833;
    wire N__13830;
    wire N__13827;
    wire N__13824;
    wire N__13821;
    wire N__13818;
    wire N__13815;
    wire N__13812;
    wire N__13809;
    wire N__13806;
    wire N__13803;
    wire N__13800;
    wire N__13797;
    wire N__13794;
    wire N__13791;
    wire N__13788;
    wire N__13785;
    wire N__13782;
    wire N__13779;
    wire N__13778;
    wire N__13775;
    wire N__13772;
    wire N__13767;
    wire N__13764;
    wire N__13761;
    wire N__13758;
    wire N__13757;
    wire N__13754;
    wire N__13753;
    wire N__13750;
    wire N__13747;
    wire N__13744;
    wire N__13737;
    wire N__13736;
    wire N__13733;
    wire N__13730;
    wire N__13729;
    wire N__13724;
    wire N__13721;
    wire N__13716;
    wire N__13713;
    wire N__13710;
    wire N__13709;
    wire N__13706;
    wire N__13703;
    wire N__13698;
    wire N__13695;
    wire N__13694;
    wire N__13691;
    wire N__13690;
    wire N__13687;
    wire N__13684;
    wire N__13681;
    wire N__13674;
    wire N__13673;
    wire N__13670;
    wire N__13667;
    wire N__13662;
    wire N__13659;
    wire N__13656;
    wire N__13653;
    wire N__13650;
    wire N__13647;
    wire N__13644;
    wire N__13641;
    wire N__13638;
    wire N__13635;
    wire N__13632;
    wire N__13629;
    wire N__13626;
    wire N__13623;
    wire N__13620;
    wire N__13617;
    wire N__13614;
    wire N__13611;
    wire N__13610;
    wire N__13607;
    wire N__13604;
    wire N__13601;
    wire N__13598;
    wire N__13593;
    wire N__13590;
    wire N__13587;
    wire N__13584;
    wire N__13581;
    wire N__13580;
    wire N__13577;
    wire N__13574;
    wire N__13573;
    wire N__13572;
    wire N__13571;
    wire N__13570;
    wire N__13567;
    wire N__13564;
    wire N__13561;
    wire N__13558;
    wire N__13555;
    wire N__13554;
    wire N__13553;
    wire N__13550;
    wire N__13549;
    wire N__13546;
    wire N__13541;
    wire N__13536;
    wire N__13533;
    wire N__13530;
    wire N__13527;
    wire N__13524;
    wire N__13521;
    wire N__13518;
    wire N__13515;
    wire N__13512;
    wire N__13509;
    wire N__13506;
    wire N__13503;
    wire N__13500;
    wire N__13491;
    wire N__13488;
    wire N__13485;
    wire N__13476;
    wire N__13473;
    wire N__13470;
    wire N__13467;
    wire N__13464;
    wire N__13461;
    wire N__13460;
    wire N__13457;
    wire N__13454;
    wire N__13451;
    wire N__13448;
    wire N__13445;
    wire N__13442;
    wire N__13439;
    wire N__13436;
    wire N__13433;
    wire N__13430;
    wire N__13427;
    wire N__13424;
    wire N__13421;
    wire N__13418;
    wire N__13415;
    wire N__13412;
    wire N__13409;
    wire N__13406;
    wire N__13403;
    wire N__13400;
    wire N__13397;
    wire N__13394;
    wire N__13391;
    wire N__13388;
    wire N__13385;
    wire N__13382;
    wire N__13379;
    wire N__13376;
    wire N__13373;
    wire N__13370;
    wire N__13367;
    wire N__13364;
    wire N__13361;
    wire N__13358;
    wire N__13355;
    wire N__13352;
    wire N__13349;
    wire N__13346;
    wire N__13343;
    wire N__13340;
    wire N__13337;
    wire N__13334;
    wire N__13331;
    wire N__13328;
    wire N__13325;
    wire N__13322;
    wire N__13319;
    wire N__13316;
    wire N__13313;
    wire N__13310;
    wire N__13307;
    wire N__13304;
    wire N__13301;
    wire N__13298;
    wire N__13295;
    wire N__13292;
    wire N__13289;
    wire N__13286;
    wire N__13283;
    wire N__13280;
    wire N__13277;
    wire N__13274;
    wire N__13271;
    wire N__13268;
    wire N__13265;
    wire N__13262;
    wire N__13259;
    wire N__13256;
    wire N__13253;
    wire N__13250;
    wire N__13247;
    wire N__13242;
    wire N__13239;
    wire N__13236;
    wire N__13235;
    wire N__13232;
    wire N__13229;
    wire N__13226;
    wire N__13223;
    wire N__13220;
    wire N__13217;
    wire N__13214;
    wire N__13211;
    wire N__13208;
    wire N__13205;
    wire N__13202;
    wire N__13199;
    wire N__13196;
    wire N__13193;
    wire N__13190;
    wire N__13187;
    wire N__13184;
    wire N__13181;
    wire N__13178;
    wire N__13175;
    wire N__13172;
    wire N__13169;
    wire N__13166;
    wire N__13163;
    wire N__13160;
    wire N__13157;
    wire N__13154;
    wire N__13151;
    wire N__13148;
    wire N__13145;
    wire N__13142;
    wire N__13139;
    wire N__13136;
    wire N__13133;
    wire N__13130;
    wire N__13127;
    wire N__13124;
    wire N__13121;
    wire N__13118;
    wire N__13115;
    wire N__13112;
    wire N__13109;
    wire N__13106;
    wire N__13103;
    wire N__13100;
    wire N__13097;
    wire N__13094;
    wire N__13091;
    wire N__13088;
    wire N__13085;
    wire N__13082;
    wire N__13079;
    wire N__13076;
    wire N__13073;
    wire N__13070;
    wire N__13067;
    wire N__13064;
    wire N__13061;
    wire N__13058;
    wire N__13055;
    wire N__13052;
    wire N__13049;
    wire N__13046;
    wire N__13043;
    wire N__13040;
    wire N__13037;
    wire N__13032;
    wire N__13029;
    wire N__13026;
    wire N__13023;
    wire N__13020;
    wire N__13017;
    wire N__13014;
    wire N__13011;
    wire N__13008;
    wire N__13005;
    wire N__13002;
    wire N__12999;
    wire N__12996;
    wire N__12995;
    wire N__12992;
    wire N__12989;
    wire N__12984;
    wire N__12981;
    wire N__12980;
    wire N__12977;
    wire N__12974;
    wire N__12971;
    wire N__12968;
    wire N__12965;
    wire N__12962;
    wire N__12959;
    wire N__12956;
    wire N__12953;
    wire N__12950;
    wire N__12947;
    wire N__12944;
    wire N__12941;
    wire N__12938;
    wire N__12935;
    wire N__12932;
    wire N__12929;
    wire N__12926;
    wire N__12923;
    wire N__12920;
    wire N__12917;
    wire N__12914;
    wire N__12911;
    wire N__12908;
    wire N__12905;
    wire N__12902;
    wire N__12899;
    wire N__12896;
    wire N__12893;
    wire N__12890;
    wire N__12887;
    wire N__12884;
    wire N__12881;
    wire N__12878;
    wire N__12875;
    wire N__12872;
    wire N__12869;
    wire N__12866;
    wire N__12863;
    wire N__12860;
    wire N__12857;
    wire N__12854;
    wire N__12851;
    wire N__12848;
    wire N__12845;
    wire N__12842;
    wire N__12839;
    wire N__12836;
    wire N__12833;
    wire N__12830;
    wire N__12827;
    wire N__12824;
    wire N__12821;
    wire N__12818;
    wire N__12815;
    wire N__12812;
    wire N__12809;
    wire N__12806;
    wire N__12803;
    wire N__12800;
    wire N__12797;
    wire N__12794;
    wire N__12791;
    wire N__12788;
    wire N__12785;
    wire N__12782;
    wire N__12779;
    wire N__12776;
    wire N__12773;
    wire N__12770;
    wire N__12767;
    wire N__12764;
    wire N__12759;
    wire N__12756;
    wire N__12755;
    wire N__12752;
    wire N__12749;
    wire N__12744;
    wire N__12743;
    wire N__12740;
    wire N__12737;
    wire N__12732;
    wire N__12729;
    wire N__12728;
    wire N__12725;
    wire N__12722;
    wire N__12719;
    wire N__12716;
    wire N__12713;
    wire N__12710;
    wire N__12707;
    wire N__12704;
    wire N__12701;
    wire N__12698;
    wire N__12695;
    wire N__12692;
    wire N__12689;
    wire N__12686;
    wire N__12683;
    wire N__12680;
    wire N__12677;
    wire N__12674;
    wire N__12671;
    wire N__12668;
    wire N__12665;
    wire N__12662;
    wire N__12659;
    wire N__12656;
    wire N__12653;
    wire N__12650;
    wire N__12647;
    wire N__12644;
    wire N__12641;
    wire N__12638;
    wire N__12635;
    wire N__12632;
    wire N__12629;
    wire N__12626;
    wire N__12623;
    wire N__12620;
    wire N__12617;
    wire N__12614;
    wire N__12611;
    wire N__12608;
    wire N__12605;
    wire N__12602;
    wire N__12599;
    wire N__12596;
    wire N__12593;
    wire N__12590;
    wire N__12587;
    wire N__12584;
    wire N__12581;
    wire N__12578;
    wire N__12575;
    wire N__12572;
    wire N__12569;
    wire N__12566;
    wire N__12563;
    wire N__12560;
    wire N__12557;
    wire N__12554;
    wire N__12551;
    wire N__12548;
    wire N__12545;
    wire N__12542;
    wire N__12539;
    wire N__12536;
    wire N__12533;
    wire N__12530;
    wire N__12527;
    wire N__12524;
    wire N__12521;
    wire N__12518;
    wire N__12515;
    wire N__12512;
    wire N__12507;
    wire N__12504;
    wire N__12501;
    wire N__12500;
    wire N__12499;
    wire N__12498;
    wire N__12495;
    wire N__12492;
    wire N__12489;
    wire N__12484;
    wire N__12477;
    wire N__12474;
    wire N__12471;
    wire N__12468;
    wire N__12465;
    wire N__12462;
    wire N__12461;
    wire N__12460;
    wire N__12457;
    wire N__12454;
    wire N__12453;
    wire N__12450;
    wire N__12445;
    wire N__12442;
    wire N__12435;
    wire N__12432;
    wire N__12429;
    wire N__12428;
    wire N__12427;
    wire N__12426;
    wire N__12423;
    wire N__12420;
    wire N__12415;
    wire N__12412;
    wire N__12405;
    wire N__12402;
    wire N__12399;
    wire N__12398;
    wire N__12397;
    wire N__12396;
    wire N__12393;
    wire N__12390;
    wire N__12385;
    wire N__12382;
    wire N__12375;
    wire N__12372;
    wire N__12369;
    wire N__12366;
    wire N__12363;
    wire N__12362;
    wire N__12361;
    wire N__12360;
    wire N__12357;
    wire N__12354;
    wire N__12351;
    wire N__12348;
    wire N__12339;
    wire N__12336;
    wire N__12333;
    wire N__12330;
    wire N__12327;
    wire N__12324;
    wire N__12321;
    wire N__12318;
    wire N__12315;
    wire N__12312;
    wire N__12309;
    wire N__12306;
    wire N__12303;
    wire N__12300;
    wire N__12297;
    wire N__12294;
    wire N__12291;
    wire N__12288;
    wire N__12285;
    wire N__12282;
    wire N__12279;
    wire N__12276;
    wire N__12273;
    wire N__12272;
    wire N__12269;
    wire N__12266;
    wire N__12263;
    wire N__12258;
    wire N__12257;
    wire N__12256;
    wire N__12255;
    wire N__12252;
    wire N__12249;
    wire N__12246;
    wire N__12243;
    wire N__12242;
    wire N__12237;
    wire N__12234;
    wire N__12231;
    wire N__12228;
    wire N__12225;
    wire N__12220;
    wire N__12213;
    wire N__12210;
    wire N__12209;
    wire N__12204;
    wire N__12201;
    wire N__12200;
    wire N__12199;
    wire N__12194;
    wire N__12193;
    wire N__12190;
    wire N__12189;
    wire N__12186;
    wire N__12183;
    wire N__12180;
    wire N__12177;
    wire N__12174;
    wire N__12169;
    wire N__12162;
    wire N__12161;
    wire N__12160;
    wire N__12159;
    wire N__12156;
    wire N__12151;
    wire N__12150;
    wire N__12147;
    wire N__12144;
    wire N__12141;
    wire N__12138;
    wire N__12133;
    wire N__12130;
    wire N__12123;
    wire N__12120;
    wire N__12117;
    wire N__12114;
    wire N__12111;
    wire N__12108;
    wire N__12107;
    wire N__12106;
    wire N__12101;
    wire N__12100;
    wire N__12097;
    wire N__12094;
    wire N__12091;
    wire N__12084;
    wire N__12081;
    wire N__12078;
    wire N__12075;
    wire N__12074;
    wire N__12073;
    wire N__12070;
    wire N__12065;
    wire N__12064;
    wire N__12061;
    wire N__12058;
    wire N__12055;
    wire N__12048;
    wire N__12045;
    wire N__12042;
    wire N__12039;
    wire N__12036;
    wire N__12033;
    wire N__12030;
    wire N__12027;
    wire N__12026;
    wire N__12025;
    wire N__12024;
    wire N__12021;
    wire N__12018;
    wire N__12013;
    wire N__12006;
    wire N__12003;
    wire N__12000;
    wire N__11997;
    wire N__11994;
    wire N__11993;
    wire N__11992;
    wire N__11991;
    wire N__11988;
    wire N__11985;
    wire N__11980;
    wire N__11973;
    wire N__11972;
    wire N__11969;
    wire N__11966;
    wire N__11961;
    wire N__11958;
    wire N__11955;
    wire N__11954;
    wire N__11953;
    wire N__11950;
    wire N__11949;
    wire N__11944;
    wire N__11941;
    wire N__11938;
    wire N__11933;
    wire N__11928;
    wire N__11927;
    wire N__11924;
    wire N__11921;
    wire N__11918;
    wire N__11913;
    wire N__11910;
    wire N__11907;
    wire N__11904;
    wire N__11901;
    wire N__11900;
    wire N__11899;
    wire N__11898;
    wire N__11895;
    wire N__11892;
    wire N__11891;
    wire N__11888;
    wire N__11885;
    wire N__11882;
    wire N__11879;
    wire N__11876;
    wire N__11873;
    wire N__11864;
    wire N__11859;
    wire N__11858;
    wire N__11857;
    wire N__11854;
    wire N__11851;
    wire N__11850;
    wire N__11847;
    wire N__11842;
    wire N__11839;
    wire N__11832;
    wire N__11829;
    wire N__11826;
    wire N__11823;
    wire N__11820;
    wire N__11817;
    wire N__11816;
    wire N__11815;
    wire N__11814;
    wire N__11813;
    wire N__11812;
    wire N__11809;
    wire N__11804;
    wire N__11799;
    wire N__11796;
    wire N__11787;
    wire N__11786;
    wire N__11785;
    wire N__11784;
    wire N__11781;
    wire N__11776;
    wire N__11773;
    wire N__11766;
    wire N__11763;
    wire N__11760;
    wire N__11759;
    wire N__11758;
    wire N__11757;
    wire N__11754;
    wire N__11747;
    wire N__11742;
    wire N__11741;
    wire N__11740;
    wire N__11739;
    wire N__11736;
    wire N__11733;
    wire N__11728;
    wire N__11721;
    wire N__11718;
    wire N__11717;
    wire N__11716;
    wire N__11713;
    wire N__11708;
    wire N__11703;
    wire N__11702;
    wire N__11701;
    wire N__11698;
    wire N__11693;
    wire N__11688;
    wire N__11685;
    wire N__11684;
    wire N__11679;
    wire N__11676;
    wire N__11675;
    wire N__11672;
    wire N__11669;
    wire N__11664;
    wire N__11663;
    wire N__11660;
    wire N__11657;
    wire N__11652;
    wire N__11649;
    wire N__11646;
    wire N__11643;
    wire N__11640;
    wire N__11637;
    wire N__11634;
    wire N__11631;
    wire N__11628;
    wire N__11625;
    wire N__11622;
    wire N__11619;
    wire N__11616;
    wire N__11613;
    wire N__11610;
    wire N__11607;
    wire N__11604;
    wire N__11601;
    wire N__11598;
    wire N__11595;
    wire N__11592;
    wire N__11589;
    wire N__11586;
    wire N__11583;
    wire N__11580;
    wire N__11577;
    wire N__11574;
    wire N__11571;
    wire N__11568;
    wire N__11565;
    wire N__11562;
    wire N__11559;
    wire N__11556;
    wire N__11553;
    wire N__11550;
    wire N__11547;
    wire N__11544;
    wire N__11541;
    wire N__11538;
    wire N__11535;
    wire N__11532;
    wire N__11529;
    wire N__11526;
    wire N__11523;
    wire N__11520;
    wire N__11519;
    wire N__11518;
    wire N__11515;
    wire N__11512;
    wire N__11509;
    wire N__11506;
    wire N__11503;
    wire N__11500;
    wire N__11497;
    wire N__11494;
    wire N__11491;
    wire N__11488;
    wire N__11485;
    wire N__11482;
    wire N__11479;
    wire N__11476;
    wire N__11469;
    wire N__11466;
    wire N__11463;
    wire N__11460;
    wire N__11457;
    wire N__11454;
    wire N__11451;
    wire N__11448;
    wire N__11445;
    wire N__11442;
    wire N__11439;
    wire N__11438;
    wire N__11435;
    wire N__11432;
    wire N__11427;
    wire N__11424;
    wire N__11421;
    wire N__11420;
    wire N__11417;
    wire N__11414;
    wire N__11411;
    wire N__11408;
    wire N__11405;
    wire N__11402;
    wire N__11399;
    wire N__11396;
    wire N__11393;
    wire N__11390;
    wire N__11387;
    wire N__11384;
    wire N__11381;
    wire N__11378;
    wire N__11375;
    wire N__11372;
    wire N__11369;
    wire N__11366;
    wire N__11363;
    wire N__11360;
    wire N__11357;
    wire N__11354;
    wire N__11351;
    wire N__11348;
    wire N__11345;
    wire N__11342;
    wire N__11339;
    wire N__11336;
    wire N__11333;
    wire N__11330;
    wire N__11327;
    wire N__11324;
    wire N__11321;
    wire N__11318;
    wire N__11315;
    wire N__11312;
    wire N__11309;
    wire N__11306;
    wire N__11303;
    wire N__11300;
    wire N__11297;
    wire N__11294;
    wire N__11291;
    wire N__11288;
    wire N__11285;
    wire N__11282;
    wire N__11279;
    wire N__11276;
    wire N__11273;
    wire N__11270;
    wire N__11267;
    wire N__11264;
    wire N__11261;
    wire N__11258;
    wire N__11255;
    wire N__11252;
    wire N__11249;
    wire N__11246;
    wire N__11243;
    wire N__11240;
    wire N__11237;
    wire N__11234;
    wire N__11231;
    wire N__11228;
    wire N__11225;
    wire N__11222;
    wire N__11219;
    wire N__11216;
    wire N__11213;
    wire N__11210;
    wire N__11207;
    wire N__11202;
    wire N__11199;
    wire N__11196;
    wire N__11193;
    wire N__11190;
    wire N__11187;
    wire N__11184;
    wire N__11181;
    wire N__11178;
    wire N__11175;
    wire N__11172;
    wire N__11171;
    wire N__11168;
    wire N__11165;
    wire N__11162;
    wire N__11159;
    wire N__11156;
    wire N__11153;
    wire N__11150;
    wire N__11147;
    wire N__11144;
    wire N__11141;
    wire N__11138;
    wire N__11135;
    wire N__11132;
    wire N__11129;
    wire N__11126;
    wire N__11123;
    wire N__11120;
    wire N__11117;
    wire N__11114;
    wire N__11111;
    wire N__11108;
    wire N__11105;
    wire N__11102;
    wire N__11099;
    wire N__11096;
    wire N__11093;
    wire N__11090;
    wire N__11087;
    wire N__11084;
    wire N__11081;
    wire N__11078;
    wire N__11075;
    wire N__11072;
    wire N__11069;
    wire N__11066;
    wire N__11063;
    wire N__11060;
    wire N__11057;
    wire N__11054;
    wire N__11051;
    wire N__11048;
    wire N__11045;
    wire N__11042;
    wire N__11039;
    wire N__11036;
    wire N__11033;
    wire N__11030;
    wire N__11027;
    wire N__11024;
    wire N__11021;
    wire N__11018;
    wire N__11015;
    wire N__11012;
    wire N__11009;
    wire N__11006;
    wire N__11003;
    wire N__11000;
    wire N__10997;
    wire N__10994;
    wire N__10991;
    wire N__10988;
    wire N__10985;
    wire N__10982;
    wire N__10979;
    wire N__10976;
    wire N__10973;
    wire N__10970;
    wire N__10967;
    wire N__10964;
    wire N__10961;
    wire N__10956;
    wire N__10953;
    wire N__10952;
    wire N__10949;
    wire N__10946;
    wire N__10941;
    wire N__10938;
    wire N__10935;
    wire N__10932;
    wire N__10929;
    wire N__10926;
    wire N__10923;
    wire N__10920;
    wire N__10919;
    wire N__10916;
    wire N__10913;
    wire N__10910;
    wire N__10907;
    wire N__10904;
    wire N__10901;
    wire N__10898;
    wire N__10895;
    wire N__10892;
    wire N__10889;
    wire N__10886;
    wire N__10883;
    wire N__10880;
    wire N__10877;
    wire N__10874;
    wire N__10871;
    wire N__10868;
    wire N__10865;
    wire N__10862;
    wire N__10859;
    wire N__10856;
    wire N__10853;
    wire N__10850;
    wire N__10847;
    wire N__10844;
    wire N__10841;
    wire N__10838;
    wire N__10835;
    wire N__10832;
    wire N__10829;
    wire N__10826;
    wire N__10823;
    wire N__10820;
    wire N__10817;
    wire N__10814;
    wire N__10811;
    wire N__10808;
    wire N__10805;
    wire N__10802;
    wire N__10799;
    wire N__10796;
    wire N__10793;
    wire N__10790;
    wire N__10787;
    wire N__10784;
    wire N__10781;
    wire N__10778;
    wire N__10775;
    wire N__10772;
    wire N__10769;
    wire N__10766;
    wire N__10763;
    wire N__10760;
    wire N__10757;
    wire N__10754;
    wire N__10751;
    wire N__10748;
    wire N__10745;
    wire N__10742;
    wire N__10739;
    wire N__10736;
    wire N__10733;
    wire N__10730;
    wire N__10727;
    wire N__10724;
    wire N__10721;
    wire N__10718;
    wire N__10715;
    wire N__10710;
    wire N__10707;
    wire N__10704;
    wire N__10701;
    wire N__10700;
    wire N__10697;
    wire N__10694;
    wire N__10689;
    wire N__10686;
    wire N__10683;
    wire N__10682;
    wire N__10677;
    wire N__10674;
    wire N__10671;
    wire N__10668;
    wire N__10665;
    wire N__10662;
    wire N__10659;
    wire N__10656;
    wire N__10655;
    wire N__10652;
    wire N__10649;
    wire N__10646;
    wire N__10643;
    wire N__10640;
    wire N__10637;
    wire N__10634;
    wire N__10631;
    wire N__10628;
    wire N__10625;
    wire N__10622;
    wire N__10619;
    wire N__10616;
    wire N__10613;
    wire N__10610;
    wire N__10607;
    wire N__10604;
    wire N__10601;
    wire N__10598;
    wire N__10595;
    wire N__10592;
    wire N__10589;
    wire N__10586;
    wire N__10583;
    wire N__10580;
    wire N__10577;
    wire N__10574;
    wire N__10571;
    wire N__10568;
    wire N__10565;
    wire N__10562;
    wire N__10559;
    wire N__10556;
    wire N__10553;
    wire N__10550;
    wire N__10547;
    wire N__10544;
    wire N__10541;
    wire N__10538;
    wire N__10535;
    wire N__10532;
    wire N__10529;
    wire N__10526;
    wire N__10523;
    wire N__10520;
    wire N__10517;
    wire N__10514;
    wire N__10511;
    wire N__10508;
    wire N__10505;
    wire N__10502;
    wire N__10499;
    wire N__10496;
    wire N__10493;
    wire N__10490;
    wire N__10487;
    wire N__10484;
    wire N__10481;
    wire N__10478;
    wire N__10475;
    wire N__10472;
    wire N__10469;
    wire N__10466;
    wire N__10463;
    wire N__10460;
    wire N__10457;
    wire N__10454;
    wire N__10451;
    wire N__10446;
    wire N__10443;
    wire N__10440;
    wire N__10439;
    wire N__10436;
    wire N__10433;
    wire N__10428;
    wire N__10425;
    wire N__10422;
    wire N__10419;
    wire N__10416;
    wire N__10413;
    wire N__10410;
    wire N__10407;
    wire N__10406;
    wire N__10403;
    wire N__10400;
    wire N__10397;
    wire N__10394;
    wire N__10391;
    wire N__10388;
    wire N__10385;
    wire N__10382;
    wire N__10379;
    wire N__10376;
    wire N__10373;
    wire N__10370;
    wire N__10367;
    wire N__10364;
    wire N__10361;
    wire N__10358;
    wire N__10355;
    wire N__10352;
    wire N__10349;
    wire N__10346;
    wire N__10343;
    wire N__10340;
    wire N__10337;
    wire N__10334;
    wire N__10331;
    wire N__10328;
    wire N__10325;
    wire N__10322;
    wire N__10319;
    wire N__10316;
    wire N__10313;
    wire N__10310;
    wire N__10307;
    wire N__10304;
    wire N__10301;
    wire N__10298;
    wire N__10295;
    wire N__10292;
    wire N__10289;
    wire N__10286;
    wire N__10283;
    wire N__10280;
    wire N__10277;
    wire N__10274;
    wire N__10271;
    wire N__10268;
    wire N__10265;
    wire N__10262;
    wire N__10259;
    wire N__10256;
    wire N__10253;
    wire N__10250;
    wire N__10247;
    wire N__10244;
    wire N__10241;
    wire N__10238;
    wire N__10235;
    wire N__10232;
    wire N__10229;
    wire N__10226;
    wire N__10223;
    wire N__10220;
    wire N__10217;
    wire N__10214;
    wire N__10211;
    wire N__10208;
    wire N__10205;
    wire N__10202;
    wire N__10199;
    wire N__10196;
    wire N__10193;
    wire N__10190;
    wire N__10185;
    wire N__10182;
    wire N__10179;
    wire N__10176;
    wire N__10173;
    wire N__10172;
    wire N__10169;
    wire N__10166;
    wire N__10163;
    wire N__10160;
    wire N__10157;
    wire N__10154;
    wire N__10151;
    wire N__10148;
    wire N__10145;
    wire N__10142;
    wire N__10139;
    wire N__10136;
    wire N__10133;
    wire N__10130;
    wire N__10127;
    wire N__10124;
    wire N__10121;
    wire N__10118;
    wire N__10115;
    wire N__10112;
    wire N__10109;
    wire N__10106;
    wire N__10103;
    wire N__10100;
    wire N__10097;
    wire N__10094;
    wire N__10091;
    wire N__10088;
    wire N__10085;
    wire N__10082;
    wire N__10079;
    wire N__10076;
    wire N__10073;
    wire N__10070;
    wire N__10067;
    wire N__10064;
    wire N__10061;
    wire N__10058;
    wire N__10055;
    wire N__10052;
    wire N__10049;
    wire N__10046;
    wire N__10043;
    wire N__10040;
    wire N__10037;
    wire N__10034;
    wire N__10031;
    wire N__10028;
    wire N__10025;
    wire N__10022;
    wire N__10019;
    wire N__10016;
    wire N__10013;
    wire N__10010;
    wire N__10007;
    wire N__10004;
    wire N__10001;
    wire N__9998;
    wire N__9995;
    wire N__9992;
    wire N__9989;
    wire N__9986;
    wire N__9983;
    wire N__9980;
    wire N__9977;
    wire N__9974;
    wire N__9971;
    wire N__9968;
    wire N__9965;
    wire N__9962;
    wire N__9959;
    wire N__9954;
    wire N__9951;
    wire N__9948;
    wire N__9945;
    wire N__9942;
    wire N__9939;
    wire N__9938;
    wire N__9937;
    wire N__9934;
    wire N__9931;
    wire N__9928;
    wire N__9925;
    wire N__9922;
    wire N__9915;
    wire N__9914;
    wire N__9913;
    wire N__9912;
    wire N__9909;
    wire N__9908;
    wire N__9905;
    wire N__9904;
    wire N__9901;
    wire N__9900;
    wire N__9899;
    wire N__9896;
    wire N__9895;
    wire N__9894;
    wire N__9891;
    wire N__9888;
    wire N__9885;
    wire N__9882;
    wire N__9879;
    wire N__9876;
    wire N__9873;
    wire N__9872;
    wire N__9869;
    wire N__9866;
    wire N__9863;
    wire N__9854;
    wire N__9847;
    wire N__9844;
    wire N__9837;
    wire N__9834;
    wire N__9831;
    wire N__9828;
    wire N__9825;
    wire N__9816;
    wire N__9815;
    wire N__9812;
    wire N__9811;
    wire N__9810;
    wire N__9807;
    wire N__9804;
    wire N__9801;
    wire N__9798;
    wire N__9791;
    wire N__9786;
    wire N__9785;
    wire N__9782;
    wire N__9781;
    wire N__9780;
    wire N__9775;
    wire N__9772;
    wire N__9769;
    wire N__9764;
    wire N__9759;
    wire N__9758;
    wire N__9757;
    wire N__9756;
    wire N__9751;
    wire N__9748;
    wire N__9745;
    wire N__9740;
    wire N__9735;
    wire N__9734;
    wire N__9733;
    wire N__9732;
    wire N__9727;
    wire N__9724;
    wire N__9721;
    wire N__9716;
    wire N__9711;
    wire N__9710;
    wire N__9709;
    wire N__9706;
    wire N__9703;
    wire N__9700;
    wire N__9695;
    wire N__9690;
    wire N__9687;
    wire N__9686;
    wire N__9685;
    wire N__9684;
    wire N__9681;
    wire N__9678;
    wire N__9675;
    wire N__9672;
    wire N__9667;
    wire N__9660;
    wire N__9659;
    wire N__9656;
    wire N__9655;
    wire N__9654;
    wire N__9651;
    wire N__9648;
    wire N__9645;
    wire N__9642;
    wire N__9639;
    wire N__9630;
    wire N__9627;
    wire N__9624;
    wire N__9621;
    wire N__9618;
    wire N__9615;
    wire N__9612;
    wire N__9609;
    wire N__9606;
    wire N__9603;
    wire N__9600;
    wire N__9597;
    wire N__9594;
    wire N__9593;
    wire N__9590;
    wire N__9587;
    wire N__9582;
    wire N__9579;
    wire N__9576;
    wire N__9573;
    wire N__9570;
    wire N__9567;
    wire N__9564;
    wire N__9561;
    wire N__9558;
    wire N__9555;
    wire N__9552;
    wire N__9549;
    wire N__9546;
    wire N__9543;
    wire N__9540;
    wire N__9537;
    wire N__9534;
    wire N__9531;
    wire N__9528;
    wire N__9525;
    wire N__9524;
    wire N__9521;
    wire N__9520;
    wire N__9519;
    wire N__9516;
    wire N__9515;
    wire N__9514;
    wire N__9513;
    wire N__9510;
    wire N__9507;
    wire N__9504;
    wire N__9503;
    wire N__9500;
    wire N__9497;
    wire N__9494;
    wire N__9491;
    wire N__9486;
    wire N__9483;
    wire N__9480;
    wire N__9473;
    wire N__9470;
    wire N__9467;
    wire N__9462;
    wire N__9457;
    wire N__9452;
    wire N__9449;
    wire N__9446;
    wire N__9441;
    wire N__9438;
    wire N__9435;
    wire N__9432;
    wire N__9429;
    wire N__9426;
    wire N__9423;
    wire N__9420;
    wire N__9419;
    wire N__9416;
    wire N__9413;
    wire N__9410;
    wire N__9407;
    wire N__9404;
    wire N__9401;
    wire N__9400;
    wire N__9397;
    wire N__9394;
    wire N__9391;
    wire N__9388;
    wire N__9385;
    wire N__9382;
    wire N__9379;
    wire N__9374;
    wire N__9369;
    wire N__9366;
    wire N__9363;
    wire N__9360;
    wire N__9357;
    wire N__9354;
    wire N__9351;
    wire N__9348;
    wire N__9345;
    wire N__9342;
    wire N__9339;
    wire N__9336;
    wire N__9335;
    wire N__9332;
    wire N__9331;
    wire N__9328;
    wire N__9325;
    wire N__9322;
    wire N__9319;
    wire N__9318;
    wire N__9313;
    wire N__9312;
    wire N__9311;
    wire N__9310;
    wire N__9307;
    wire N__9304;
    wire N__9303;
    wire N__9300;
    wire N__9297;
    wire N__9294;
    wire N__9291;
    wire N__9286;
    wire N__9283;
    wire N__9276;
    wire N__9273;
    wire N__9270;
    wire N__9267;
    wire N__9262;
    wire N__9257;
    wire N__9254;
    wire N__9251;
    wire N__9246;
    wire N__9243;
    wire N__9240;
    wire N__9237;
    wire N__9234;
    wire N__9231;
    wire N__9230;
    wire N__9227;
    wire N__9224;
    wire N__9221;
    wire N__9218;
    wire N__9215;
    wire N__9212;
    wire N__9207;
    wire N__9204;
    wire N__9201;
    wire N__9198;
    wire N__9195;
    wire N__9192;
    wire N__9189;
    wire N__9186;
    wire N__9183;
    wire N__9180;
    wire N__9177;
    wire N__9174;
    wire N__9171;
    wire N__9168;
    wire N__9165;
    wire N__9162;
    wire N__9159;
    wire N__9156;
    wire N__9153;
    wire N__9150;
    wire N__9147;
    wire N__9144;
    wire N__9141;
    wire N__9138;
    wire N__9135;
    wire N__9132;
    wire N__9129;
    wire N__9126;
    wire N__9123;
    wire N__9120;
    wire N__9117;
    wire N__9114;
    wire N__9111;
    wire N__9108;
    wire N__9105;
    wire N__9102;
    wire N__9099;
    wire N__9096;
    wire N__9093;
    wire N__9090;
    wire N__9087;
    wire N__9084;
    wire N__9081;
    wire N__9078;
    wire N__9075;
    wire N__9072;
    wire N__9069;
    wire N__9066;
    wire N__9063;
    wire N__9060;
    wire N__9057;
    wire N__9054;
    wire N__9051;
    wire N__9048;
    wire N__9045;
    wire N__9042;
    wire N__9039;
    wire N__9036;
    wire N__9033;
    wire N__9030;
    wire N__9027;
    wire N__9024;
    wire N__9021;
    wire N__9018;
    wire N__9015;
    wire N__9012;
    wire N__9009;
    wire N__9006;
    wire N__9003;
    wire N__9000;
    wire N__8997;
    wire N__8994;
    wire N__8991;
    wire N__8988;
    wire N__8985;
    wire N__8982;
    wire N__8979;
    wire N__8976;
    wire N__8973;
    wire N__8970;
    wire N__8967;
    wire N__8964;
    wire N__8961;
    wire N__8958;
    wire N__8955;
    wire N__8952;
    wire N__8949;
    wire N__8946;
    wire N__8943;
    wire N__8940;
    wire N__8937;
    wire N__8934;
    wire N__8931;
    wire N__8928;
    wire N__8925;
    wire N__8922;
    wire N__8919;
    wire N__8916;
    wire N__8913;
    wire N__8910;
    wire N__8907;
    wire N__8904;
    wire N__8901;
    wire N__8898;
    wire N__8895;
    wire N__8892;
    wire N__8889;
    wire N__8886;
    wire N__8883;
    wire N__8880;
    wire N__8877;
    wire N__8874;
    wire N__8871;
    wire N__8868;
    wire N__8865;
    wire N__8862;
    wire N__8859;
    wire N__8856;
    wire N__8853;
    wire N__8850;
    wire N__8847;
    wire N__8844;
    wire N__8841;
    wire N__8838;
    wire N__8835;
    wire N__8832;
    wire N__8829;
    wire N__8826;
    wire N__8823;
    wire N__8820;
    wire N__8817;
    wire N__8814;
    wire N__8811;
    wire N__8808;
    wire N__8805;
    wire N__8802;
    wire N__8799;
    wire N__8796;
    wire N__8793;
    wire N__8790;
    wire N__8787;
    wire N__8784;
    wire N__8781;
    wire N__8778;
    wire N__8775;
    wire N__8772;
    wire N__8769;
    wire N__8766;
    wire N__8763;
    wire N__8760;
    wire N__8757;
    wire N__8754;
    wire N__8751;
    wire N__8748;
    wire N__8745;
    wire N__8742;
    wire N__8739;
    wire N__8736;
    wire N__8733;
    wire N__8730;
    wire N__8727;
    wire N__8724;
    wire N__8721;
    wire N__8718;
    wire N__8715;
    wire N__8712;
    wire N__8709;
    wire N__8706;
    wire N__8703;
    wire N__8700;
    wire N__8697;
    wire N__8694;
    wire N__8691;
    wire N__8688;
    wire N__8685;
    wire N__8682;
    wire N__8679;
    wire N__8676;
    wire N__8673;
    wire N__8670;
    wire N__8667;
    wire N__8664;
    wire N__8661;
    wire N__8658;
    wire N__8655;
    wire N__8652;
    wire N__8649;
    wire N__8646;
    wire N__8643;
    wire N__8640;
    wire N__8637;
    wire N__8634;
    wire N__8631;
    wire N__8628;
    wire N__8625;
    wire N__8622;
    wire N__8619;
    wire N__8616;
    wire N__8613;
    wire N__8610;
    wire N__8607;
    wire N__8604;
    wire N__8601;
    wire N__8598;
    wire N__8595;
    wire N__8592;
    wire N__8589;
    wire N__8586;
    wire N__8583;
    wire N__8580;
    wire N__8577;
    wire N__8574;
    wire N__8571;
    wire N__8568;
    wire N__8565;
    wire N__8562;
    wire N__8559;
    wire N__8556;
    wire N__8553;
    wire N__8550;
    wire N__8547;
    wire N__8544;
    wire N__8541;
    wire N__8538;
    wire N__8535;
    wire N__8532;
    wire N__8529;
    wire N__8526;
    wire N__8523;
    wire N__8520;
    wire N__8517;
    wire N__8514;
    wire N__8511;
    wire N__8508;
    wire N__8505;
    wire N__8502;
    wire N__8499;
    wire N__8496;
    wire N__8493;
    wire N__8490;
    wire N__8487;
    wire N__8484;
    wire N__8481;
    wire N__8478;
    wire N__8475;
    wire N__8472;
    wire N__8469;
    wire N__8466;
    wire N__8463;
    wire N__8460;
    wire N__8457;
    wire N__8454;
    wire N__8451;
    wire N__8448;
    wire N__8445;
    wire N__8442;
    wire N__8439;
    wire N__8436;
    wire N__8433;
    wire N__8430;
    wire N__8427;
    wire N__8424;
    wire N__8421;
    wire N__8418;
    wire N__8415;
    wire N__8412;
    wire N__8409;
    wire VCCG0;
    wire GNDG0;
    wire \transmit_module.Y_DELTA_PATTERN_38 ;
    wire \transmit_module.Y_DELTA_PATTERN_55 ;
    wire \transmit_module.Y_DELTA_PATTERN_46 ;
    wire \transmit_module.Y_DELTA_PATTERN_58 ;
    wire \transmit_module.Y_DELTA_PATTERN_59 ;
    wire \transmit_module.Y_DELTA_PATTERN_57 ;
    wire \transmit_module.Y_DELTA_PATTERN_56 ;
    wire \transmit_module.Y_DELTA_PATTERN_39 ;
    wire \transmit_module.Y_DELTA_PATTERN_45 ;
    wire \line_buffer.n599 ;
    wire \line_buffer.n591 ;
    wire \line_buffer.n600 ;
    wire \line_buffer.n592 ;
    wire \transmit_module.Y_DELTA_PATTERN_28 ;
    wire \transmit_module.Y_DELTA_PATTERN_27 ;
    wire \transmit_module.Y_DELTA_PATTERN_8 ;
    wire \transmit_module.Y_DELTA_PATTERN_48 ;
    wire \transmit_module.Y_DELTA_PATTERN_47 ;
    wire \transmit_module.Y_DELTA_PATTERN_50 ;
    wire \transmit_module.Y_DELTA_PATTERN_49 ;
    wire \transmit_module.Y_DELTA_PATTERN_54 ;
    wire \transmit_module.Y_DELTA_PATTERN_67 ;
    wire \transmit_module.Y_DELTA_PATTERN_77 ;
    wire \transmit_module.Y_DELTA_PATTERN_69 ;
    wire \transmit_module.Y_DELTA_PATTERN_68 ;
    wire \transmit_module.Y_DELTA_PATTERN_76 ;
    wire \transmit_module.Y_DELTA_PATTERN_66 ;
    wire \transmit_module.Y_DELTA_PATTERN_44 ;
    wire \transmit_module.Y_DELTA_PATTERN_43 ;
    wire \transmit_module.Y_DELTA_PATTERN_42 ;
    wire \transmit_module.Y_DELTA_PATTERN_41 ;
    wire \transmit_module.Y_DELTA_PATTERN_40 ;
    wire \transmit_module.Y_DELTA_PATTERN_60 ;
    wire \transmit_module.Y_DELTA_PATTERN_7 ;
    wire \transmit_module.Y_DELTA_PATTERN_6 ;
    wire \transmit_module.Y_DELTA_PATTERN_5 ;
    wire \transmit_module.Y_DELTA_PATTERN_4 ;
    wire \line_buffer.n466 ;
    wire \line_buffer.n458 ;
    wire \line_buffer.n531 ;
    wire \line_buffer.n523 ;
    wire TVP_VIDEO_c_4;
    wire \transmit_module.Y_DELTA_PATTERN_9 ;
    wire \transmit_module.Y_DELTA_PATTERN_29 ;
    wire \transmit_module.Y_DELTA_PATTERN_30 ;
    wire \transmit_module.Y_DELTA_PATTERN_32 ;
    wire \transmit_module.Y_DELTA_PATTERN_31 ;
    wire \transmit_module.Y_DELTA_PATTERN_33 ;
    wire \transmit_module.Y_DELTA_PATTERN_37 ;
    wire \transmit_module.Y_DELTA_PATTERN_36 ;
    wire \transmit_module.Y_DELTA_PATTERN_35 ;
    wire \transmit_module.Y_DELTA_PATTERN_34 ;
    wire \transmit_module.Y_DELTA_PATTERN_81 ;
    wire \transmit_module.Y_DELTA_PATTERN_82 ;
    wire \transmit_module.Y_DELTA_PATTERN_80 ;
    wire \transmit_module.Y_DELTA_PATTERN_51 ;
    wire \transmit_module.Y_DELTA_PATTERN_70 ;
    wire \transmit_module.Y_DELTA_PATTERN_71 ;
    wire \transmit_module.Y_DELTA_PATTERN_79 ;
    wire \transmit_module.Y_DELTA_PATTERN_78 ;
    wire \transmit_module.Y_DELTA_PATTERN_72 ;
    wire \transmit_module.Y_DELTA_PATTERN_75 ;
    wire \transmit_module.Y_DELTA_PATTERN_53 ;
    wire \transmit_module.Y_DELTA_PATTERN_52 ;
    wire \transmit_module.Y_DELTA_PATTERN_74 ;
    wire \transmit_module.Y_DELTA_PATTERN_73 ;
    wire \transmit_module.Y_DELTA_PATTERN_61 ;
    wire \transmit_module.Y_DELTA_PATTERN_65 ;
    wire \transmit_module.Y_DELTA_PATTERN_64 ;
    wire \transmit_module.Y_DELTA_PATTERN_63 ;
    wire \transmit_module.Y_DELTA_PATTERN_62 ;
    wire \line_buffer.n3569 ;
    wire \line_buffer.n3566 ;
    wire \line_buffer.n3599_cascade_ ;
    wire \line_buffer.n595 ;
    wire \line_buffer.n587 ;
    wire \line_buffer.n3570 ;
    wire TVP_VIDEO_c_3;
    wire \tvp_video_buffer.BUFFER_0_3 ;
    wire \transmit_module.Y_DELTA_PATTERN_12 ;
    wire \transmit_module.Y_DELTA_PATTERN_11 ;
    wire \transmit_module.Y_DELTA_PATTERN_10 ;
    wire \sync_buffer.BUFFER_0_0 ;
    wire \sync_buffer.BUFFER_1_0 ;
    wire RX_TX_SYNC_BUFF;
    wire \transmit_module.video_signal_controller.n3479_cascade_ ;
    wire \transmit_module.video_signal_controller.n3475_cascade_ ;
    wire \transmit_module.video_signal_controller.n55 ;
    wire \line_buffer.n563 ;
    wire \line_buffer.n555 ;
    wire \line_buffer.n3567 ;
    wire bfn_12_16_0_;
    wire \transmit_module.video_signal_controller.n3180 ;
    wire \transmit_module.video_signal_controller.n3181 ;
    wire \transmit_module.video_signal_controller.n3182 ;
    wire \transmit_module.video_signal_controller.n3183 ;
    wire \transmit_module.video_signal_controller.n3184 ;
    wire \transmit_module.video_signal_controller.n3185 ;
    wire \transmit_module.video_signal_controller.n3186 ;
    wire \transmit_module.video_signal_controller.n3187 ;
    wire bfn_12_17_0_;
    wire \transmit_module.video_signal_controller.n3188 ;
    wire \transmit_module.video_signal_controller.n3189 ;
    wire \transmit_module.video_signal_controller.n3190 ;
    wire \transmit_module.Y_DELTA_PATTERN_3 ;
    wire \transmit_module.Y_DELTA_PATTERN_2 ;
    wire \transmit_module.Y_DELTA_PATTERN_1 ;
    wire \line_buffer.n536 ;
    wire \line_buffer.n528 ;
    wire \line_buffer.n3528 ;
    wire \line_buffer.n3527 ;
    wire TX_DATA_2;
    wire n1816;
    wire \line_buffer.n471 ;
    wire \line_buffer.n463 ;
    wire \tvp_video_buffer.BUFFER_1_3 ;
    wire RX_DATA_1;
    wire \tvp_video_buffer.BUFFER_1_7 ;
    wire DEBUG_c_6_c;
    wire \tvp_video_buffer.BUFFER_0_7 ;
    wire \tvp_video_buffer.BUFFER_0_4 ;
    wire \transmit_module.Y_DELTA_PATTERN_17 ;
    wire \transmit_module.Y_DELTA_PATTERN_16 ;
    wire \transmit_module.Y_DELTA_PATTERN_13 ;
    wire \transmit_module.Y_DELTA_PATTERN_15 ;
    wire \transmit_module.Y_DELTA_PATTERN_14 ;
    wire \transmit_module.Y_DELTA_PATTERN_18 ;
    wire \tvp_video_buffer.BUFFER_1_4 ;
    wire RX_DATA_2;
    wire bfn_13_12_0_;
    wire \transmit_module.video_signal_controller.n3191 ;
    wire \transmit_module.video_signal_controller.n3192 ;
    wire \transmit_module.video_signal_controller.n3193 ;
    wire \transmit_module.video_signal_controller.n3194 ;
    wire \transmit_module.video_signal_controller.n3195 ;
    wire \transmit_module.video_signal_controller.n3196 ;
    wire \transmit_module.video_signal_controller.n3197 ;
    wire \transmit_module.video_signal_controller.n3198 ;
    wire bfn_13_13_0_;
    wire \transmit_module.video_signal_controller.n3199 ;
    wire \transmit_module.video_signal_controller.n3200 ;
    wire \transmit_module.video_signal_controller.n3201 ;
    wire \transmit_module.video_signal_controller.n2395 ;
    wire \transmit_module.video_signal_controller.n7 ;
    wire \transmit_module.video_signal_controller.VGA_X_0 ;
    wire \transmit_module.n3680 ;
    wire \transmit_module.video_signal_controller.VGA_X_4 ;
    wire \transmit_module.video_signal_controller.VGA_X_3 ;
    wire \transmit_module.video_signal_controller.VGA_X_5 ;
    wire \transmit_module.video_signal_controller.VGA_X_6 ;
    wire \transmit_module.video_signal_controller.VGA_X_7 ;
    wire \transmit_module.video_signal_controller.n2014_cascade_ ;
    wire \transmit_module.video_signal_controller.VGA_X_2 ;
    wire \transmit_module.video_signal_controller.VGA_X_1 ;
    wire \transmit_module.video_signal_controller.n3676 ;
    wire \transmit_module.n146 ;
    wire \transmit_module.n146_cascade_ ;
    wire n27;
    wire \transmit_module.n107_cascade_ ;
    wire \transmit_module.n145_cascade_ ;
    wire \transmit_module.n115 ;
    wire \transmit_module.n142 ;
    wire \transmit_module.n142_cascade_ ;
    wire n23;
    wire \transmit_module.n111 ;
    wire \transmit_module.n138 ;
    wire \transmit_module.n138_cascade_ ;
    wire \transmit_module.n107 ;
    wire n19;
    wire \transmit_module.n139 ;
    wire \transmit_module.n108 ;
    wire \transmit_module.n139_cascade_ ;
    wire n20;
    wire \transmit_module.ADDR_Y_COMPONENT_10 ;
    wire \transmit_module.n145 ;
    wire n26;
    wire \transmit_module.n114 ;
    wire \transmit_module.n144 ;
    wire \transmit_module.n144_cascade_ ;
    wire n25;
    wire \transmit_module.n113 ;
    wire \transmit_module.ADDR_Y_COMPONENT_2 ;
    wire \transmit_module.ADDR_Y_COMPONENT_3 ;
    wire \line_buffer.n568 ;
    wire \line_buffer.n560 ;
    wire \line_buffer.n3530 ;
    wire \line_buffer.n3531_cascade_ ;
    wire \line_buffer.n3617 ;
    wire TX_DATA_7;
    wire ADV_B_c;
    wire \transmit_module.Y_DELTA_PATTERN_26 ;
    wire \transmit_module.Y_DELTA_PATTERN_25 ;
    wire \transmit_module.Y_DELTA_PATTERN_19 ;
    wire \transmit_module.Y_DELTA_PATTERN_20 ;
    wire \transmit_module.Y_DELTA_PATTERN_21 ;
    wire \transmit_module.Y_DELTA_PATTERN_22 ;
    wire \transmit_module.Y_DELTA_PATTERN_24 ;
    wire \transmit_module.Y_DELTA_PATTERN_23 ;
    wire \transmit_module.X_DELTA_PATTERN_13 ;
    wire \transmit_module.X_DELTA_PATTERN_14 ;
    wire \transmit_module.X_DELTA_PATTERN_6 ;
    wire \transmit_module.X_DELTA_PATTERN_5 ;
    wire \transmit_module.X_DELTA_PATTERN_4 ;
    wire \transmit_module.video_signal_controller.n6_adj_622_cascade_ ;
    wire \transmit_module.video_signal_controller.VGA_Y_3 ;
    wire \transmit_module.video_signal_controller.VGA_Y_4 ;
    wire \transmit_module.video_signal_controller.n3482_cascade_ ;
    wire \transmit_module.video_signal_controller.VGA_Y_6 ;
    wire \transmit_module.video_signal_controller.VGA_Y_5 ;
    wire \transmit_module.video_signal_controller.n6_cascade_ ;
    wire \transmit_module.video_signal_controller.n2016 ;
    wire \transmit_module.video_signal_controller.VGA_Y_8 ;
    wire \transmit_module.video_signal_controller.VGA_Y_7 ;
    wire \transmit_module.video_signal_controller.VGA_Y_2 ;
    wire \transmit_module.video_signal_controller.n3517 ;
    wire \transmit_module.video_signal_controller.VGA_Y_1 ;
    wire \transmit_module.video_signal_controller.VGA_Y_0 ;
    wire \transmit_module.video_signal_controller.n2955 ;
    wire \transmit_module.video_signal_controller.VGA_X_8 ;
    wire \transmit_module.video_signal_controller.n3363 ;
    wire \transmit_module.video_signal_controller.n2014 ;
    wire \transmit_module.video_signal_controller.n2972_cascade_ ;
    wire \transmit_module.video_signal_controller.n2047 ;
    wire \transmit_module.VGA_VISIBLE_Y ;
    wire ADV_HSYNC_c;
    wire \transmit_module.old_VGA_HS ;
    wire \transmit_module.n3675_cascade_ ;
    wire \transmit_module.video_signal_controller.n6_adj_623_cascade_ ;
    wire \transmit_module.video_signal_controller.VGA_VISIBLE_N_588 ;
    wire \transmit_module.video_signal_controller.VGA_X_11 ;
    wire \transmit_module.video_signal_controller.n7_adj_624_cascade_ ;
    wire \transmit_module.video_signal_controller.n3004 ;
    wire \transmit_module.video_signal_controller.VGA_X_10 ;
    wire \transmit_module.video_signal_controller.VGA_X_9 ;
    wire \transmit_module.video_signal_controller.n3014 ;
    wire bfn_14_15_0_;
    wire \transmit_module.n131 ;
    wire \transmit_module.n3159 ;
    wire \transmit_module.TX_ADDR_2 ;
    wire \transmit_module.n130 ;
    wire \transmit_module.n3160 ;
    wire \transmit_module.TX_ADDR_3 ;
    wire \transmit_module.n129 ;
    wire \transmit_module.n3161 ;
    wire \transmit_module.n3162 ;
    wire \transmit_module.n127 ;
    wire \transmit_module.n3163 ;
    wire \transmit_module.n3164 ;
    wire \transmit_module.n3165 ;
    wire \transmit_module.n3166 ;
    wire \transmit_module.n124 ;
    wire bfn_14_16_0_;
    wire \transmit_module.n123 ;
    wire \transmit_module.n3167 ;
    wire \transmit_module.n3168 ;
    wire \transmit_module.n3169 ;
    wire \transmit_module.n3170 ;
    wire \transmit_module.n3171 ;
    wire \transmit_module.TX_ADDR_9 ;
    wire \transmit_module.ADDR_Y_COMPONENT_9 ;
    wire \transmit_module.ADDR_Y_COMPONENT_0 ;
    wire \transmit_module.TX_ADDR_1 ;
    wire \transmit_module.ADDR_Y_COMPONENT_1 ;
    wire \transmit_module.TX_ADDR_8 ;
    wire \transmit_module.ADDR_Y_COMPONENT_8 ;
    wire \transmit_module.TX_ADDR_5 ;
    wire \transmit_module.ADDR_Y_COMPONENT_5 ;
    wire \transmit_module.TX_ADDR_10 ;
    wire \transmit_module.n122 ;
    wire n22;
    wire \transmit_module.n112_cascade_ ;
    wire n24;
    wire \transmit_module.n125 ;
    wire \transmit_module.n140 ;
    wire \transmit_module.n140_cascade_ ;
    wire \transmit_module.n109 ;
    wire n21;
    wire \transmit_module.n106 ;
    wire \transmit_module.n137 ;
    wire n18;
    wire TVP_VIDEO_c_5;
    wire DEBUG_c_1_c;
    wire \tvp_vs_buffer.BUFFER_0_0 ;
    wire \tvp_vs_buffer.BUFFER_1_0 ;
    wire RX_DATA_5;
    wire \receive_module.sync_wd.n6_cascade_ ;
    wire \receive_module.sync_wd.n4_cascade_ ;
    wire \receive_module.sync_wd.old_visible ;
    wire bfn_15_10_0_;
    wire \receive_module.rx_counter.n3207 ;
    wire \receive_module.rx_counter.n3208 ;
    wire \receive_module.rx_counter.n3209 ;
    wire \receive_module.rx_counter.n3210 ;
    wire \receive_module.rx_counter.n3211 ;
    wire \receive_module.rx_counter.n3212 ;
    wire \receive_module.rx_counter.n3213 ;
    wire \receive_module.rx_counter.n3214 ;
    wire bfn_15_11_0_;
    wire \receive_module.rx_counter.n3215 ;
    wire \tvp_vs_buffer.BUFFER_2_0 ;
    wire \transmit_module.video_signal_controller.VGA_Y_11 ;
    wire \transmit_module.video_signal_controller.VGA_Y_10 ;
    wire \transmit_module.video_signal_controller.n3461 ;
    wire \transmit_module.video_signal_controller.n3375 ;
    wire \transmit_module.video_signal_controller.n3673_cascade_ ;
    wire \transmit_module.video_signal_controller.VGA_Y_9 ;
    wire \transmit_module.video_signal_controller.n3379 ;
    wire \transmit_module.X_DELTA_PATTERN_8 ;
    wire \transmit_module.X_DELTA_PATTERN_7 ;
    wire \transmit_module.X_DELTA_PATTERN_3 ;
    wire \transmit_module.X_DELTA_PATTERN_9 ;
    wire \transmit_module.X_DELTA_PATTERN_10 ;
    wire \transmit_module.X_DELTA_PATTERN_12 ;
    wire \transmit_module.X_DELTA_PATTERN_11 ;
    wire \transmit_module.X_DELTA_PATTERN_2 ;
    wire \transmit_module.X_DELTA_PATTERN_1 ;
    wire \transmit_module.n126 ;
    wire \transmit_module.n141 ;
    wire \transmit_module.n141_cascade_ ;
    wire \transmit_module.n110 ;
    wire \transmit_module.n132 ;
    wire \transmit_module.n147_cascade_ ;
    wire n28;
    wire \transmit_module.VGA_VISIBLE ;
    wire \transmit_module.n128 ;
    wire \transmit_module.n143 ;
    wire \transmit_module.n112 ;
    wire \transmit_module.n143_cascade_ ;
    wire \transmit_module.n116 ;
    wire \transmit_module.n147 ;
    wire \transmit_module.TX_ADDR_0 ;
    wire bfn_15_16_0_;
    wire \receive_module.n3146 ;
    wire \receive_module.n3147 ;
    wire \receive_module.n3148 ;
    wire \receive_module.n3149 ;
    wire \receive_module.n3150 ;
    wire \receive_module.n3151 ;
    wire \receive_module.n3152 ;
    wire \receive_module.n3153 ;
    wire bfn_15_17_0_;
    wire \receive_module.n3154 ;
    wire \receive_module.n3155 ;
    wire \receive_module.n3156 ;
    wire \receive_module.n3157 ;
    wire \receive_module.n3158 ;
    wire \transmit_module.TX_ADDR_4 ;
    wire \transmit_module.ADDR_Y_COMPONENT_4 ;
    wire \transmit_module.TX_ADDR_7 ;
    wire \transmit_module.ADDR_Y_COMPONENT_7 ;
    wire \transmit_module.TX_ADDR_6 ;
    wire \transmit_module.ADDR_Y_COMPONENT_6 ;
    wire \transmit_module.n2310 ;
    wire \receive_module.n136 ;
    wire RX_ADDR_1;
    wire \receive_module.n127 ;
    wire RX_ADDR_10;
    wire \receive_module.n137 ;
    wire RX_ADDR_0;
    wire n1818;
    wire \receive_module.n135 ;
    wire RX_ADDR_2;
    wire \tvp_video_buffer.BUFFER_0_5 ;
    wire \receive_module.rx_counter.n3452_cascade_ ;
    wire \tvp_video_buffer.BUFFER_1_5 ;
    wire RX_DATA_3;
    wire \receive_module.rx_counter.n10 ;
    wire \receive_module.rx_counter.n14_cascade_ ;
    wire RX_TX_SYNC;
    wire \receive_module.rx_counter.n4 ;
    wire \receive_module.rx_counter.n5_cascade_ ;
    wire \receive_module.rx_counter.n3450 ;
    wire \receive_module.rx_counter.n3677 ;
    wire \receive_module.rx_counter.n3 ;
    wire \receive_module.rx_counter.X_1 ;
    wire \receive_module.rx_counter.X_2 ;
    wire \receive_module.rx_counter.X_0 ;
    wire bfn_16_12_0_;
    wire \receive_module.rx_counter.n3202 ;
    wire \receive_module.rx_counter.n3203 ;
    wire \receive_module.rx_counter.n3204 ;
    wire \receive_module.rx_counter.n3205 ;
    wire \receive_module.rx_counter.n3206 ;
    wire \receive_module.rx_counter.n6 ;
    wire \receive_module.rx_counter.n7 ;
    wire \receive_module.rx_counter.FRAME_COUNTER_5 ;
    wire \receive_module.rx_counter.FRAME_COUNTER_1 ;
    wire \receive_module.rx_counter.X_3 ;
    wire \receive_module.rx_counter.X_5 ;
    wire \receive_module.rx_counter.X_4 ;
    wire \receive_module.rx_counter.n3222 ;
    wire \receive_module.rx_counter.X_7 ;
    wire \receive_module.rx_counter.n3455_cascade_ ;
    wire \receive_module.rx_counter.X_6 ;
    wire \receive_module.rx_counter.X_8 ;
    wire \receive_module.rx_counter.X_9 ;
    wire \receive_module.rx_counter.n39_cascade_ ;
    wire \receive_module.rx_counter.n3426 ;
    wire \receive_module.rx_counter.n3478 ;
    wire \receive_module.rx_counter.n54_cascade_ ;
    wire \receive_module.rx_counter.n4_adj_612 ;
    wire \line_buffer.n473 ;
    wire \line_buffer.n570 ;
    wire \line_buffer.n571 ;
    wire \transmit_module.ADDR_Y_COMPONENT_11 ;
    wire \transmit_module.n121 ;
    wire \transmit_module.ADDR_Y_COMPONENT_13 ;
    wire \transmit_module.n119 ;
    wire \transmit_module.ADDR_Y_COMPONENT_12 ;
    wire \transmit_module.n3675 ;
    wire \transmit_module.n120 ;
    wire \transmit_module.n2070 ;
    wire \receive_module.n3671 ;
    wire \line_buffer.n603 ;
    wire \line_buffer.n539 ;
    wire \line_buffer.n474 ;
    wire \receive_module.n128 ;
    wire RX_ADDR_9;
    wire \receive_module.n134 ;
    wire RX_ADDR_3;
    wire \receive_module.n133 ;
    wire RX_ADDR_4;
    wire \receive_module.n129 ;
    wire RX_ADDR_8;
    wire \receive_module.n131 ;
    wire RX_ADDR_6;
    wire \receive_module.n130 ;
    wire RX_ADDR_7;
    wire \line_buffer.n564 ;
    wire \line_buffer.n556 ;
    wire \line_buffer.n532 ;
    wire \line_buffer.n524 ;
    wire \line_buffer.n467 ;
    wire \line_buffer.n459 ;
    wire \line_buffer.n3587 ;
    wire \line_buffer.n3590_cascade_ ;
    wire \line_buffer.n3626 ;
    wire TX_DATA_3;
    wire n1815;
    wire \line_buffer.n602 ;
    wire GB_BUFFER_DEBUG_c_3_c_THRU_CO;
    wire DEBUG_c_0;
    wire LED_c;
    wire TVP_VIDEO_c_2;
    wire \tvp_video_buffer.BUFFER_0_2 ;
    wire \receive_module.rx_counter.Y_0 ;
    wire bfn_17_9_0_;
    wire \receive_module.rx_counter.Y_1 ;
    wire \receive_module.rx_counter.n3172 ;
    wire \receive_module.rx_counter.Y_2 ;
    wire \receive_module.rx_counter.n3173 ;
    wire \receive_module.rx_counter.Y_3 ;
    wire \receive_module.rx_counter.n3174 ;
    wire \receive_module.rx_counter.Y_4 ;
    wire \receive_module.rx_counter.n3175 ;
    wire \receive_module.rx_counter.Y_5 ;
    wire \receive_module.rx_counter.n3176 ;
    wire \receive_module.rx_counter.Y_6 ;
    wire \receive_module.rx_counter.n3177 ;
    wire \receive_module.rx_counter.Y_7 ;
    wire \receive_module.rx_counter.n3178 ;
    wire \receive_module.rx_counter.n3179 ;
    wire bfn_17_10_0_;
    wire \receive_module.rx_counter.Y_8 ;
    wire \tvp_video_buffer.BUFFER_1_2 ;
    wire RX_DATA_0;
    wire \receive_module.rx_counter.FRAME_COUNTER_4 ;
    wire \receive_module.rx_counter.FRAME_COUNTER_2 ;
    wire \receive_module.rx_counter.FRAME_COUNTER_0 ;
    wire \receive_module.rx_counter.FRAME_COUNTER_3 ;
    wire \receive_module.rx_counter.n7_adj_619_cascade_ ;
    wire \receive_module.rx_counter.n3519 ;
    wire \receive_module.rx_counter.old_VS ;
    wire \receive_module.rx_counter.n11_cascade_ ;
    wire \receive_module.rx_counter.n2547 ;
    wire \receive_module.rx_counter.n11 ;
    wire PULSE_1HZ;
    wire \receive_module.rx_counter.n3672 ;
    wire RX_ADDR_12;
    wire RX_ADDR_13;
    wire RX_ADDR_11;
    wire \line_buffer.n538 ;
    wire \transmit_module.X_DELTA_PATTERN_0 ;
    wire \transmit_module.X_DELTA_PATTERN_15 ;
    wire \transmit_module.n2084 ;
    wire DEBUG_c_7_c;
    wire RX_DATA_6;
    wire \tvp_video_buffer.BUFFER_0_8 ;
    wire \tvp_video_buffer.BUFFER_1_8 ;
    wire \line_buffer.n598 ;
    wire \line_buffer.n590 ;
    wire \line_buffer.n526 ;
    wire \line_buffer.n534 ;
    wire \line_buffer.n3593_cascade_ ;
    wire \line_buffer.n554 ;
    wire \line_buffer.n562 ;
    wire \receive_module.n132 ;
    wire DEBUG_c_4;
    wire RX_ADDR_5;
    wire \receive_module.n3674 ;
    wire \line_buffer.n596 ;
    wire \line_buffer.n588 ;
    wire \line_buffer.n3623 ;
    wire DEBUG_c_2_c;
    wire \tvp_hs_buffer.BUFFER_0_0 ;
    wire \tvp_hs_buffer.BUFFER_1_0 ;
    wire TVP_VSYNC_buff;
    wire \receive_module.rx_counter.n2078 ;
    wire TVP_HSYNC_buff;
    wire \receive_module.rx_counter.old_HS ;
    wire \transmit_module.Y_DELTA_PATTERN_98 ;
    wire \transmit_module.Y_DELTA_PATTERN_89 ;
    wire \transmit_module.Y_DELTA_PATTERN_92 ;
    wire \transmit_module.Y_DELTA_PATTERN_91 ;
    wire \transmit_module.Y_DELTA_PATTERN_90 ;
    wire \transmit_module.Y_DELTA_PATTERN_0 ;
    wire \transmit_module.Y_DELTA_PATTERN_99 ;
    wire \transmit_module.n3679 ;
    wire \line_buffer.n566 ;
    wire \line_buffer.n558 ;
    wire \line_buffer.n465 ;
    wire \line_buffer.n457 ;
    wire \line_buffer.n3629 ;
    wire \line_buffer.n561 ;
    wire \line_buffer.n553 ;
    wire \line_buffer.n456 ;
    wire \line_buffer.n464 ;
    wire \line_buffer.n3635_cascade_ ;
    wire \line_buffer.n469 ;
    wire \line_buffer.n461 ;
    wire \line_buffer.n3653 ;
    wire \line_buffer.n3656_cascade_ ;
    wire \line_buffer.n3596 ;
    wire \line_buffer.n3638 ;
    wire TX_DATA_0;
    wire \line_buffer.n530 ;
    wire \line_buffer.n522 ;
    wire \line_buffer.n3632 ;
    wire \line_buffer.n3650_cascade_ ;
    wire \line_buffer.n594 ;
    wire \line_buffer.n586 ;
    wire \line_buffer.n3647 ;
    wire \line_buffer.n521 ;
    wire \line_buffer.n529 ;
    wire \line_buffer.n3644 ;
    wire TX_DATA_5;
    wire n1813;
    wire TX_DATA_1;
    wire n1817;
    wire \transmit_module.Y_DELTA_PATTERN_97 ;
    wire \transmit_module.Y_DELTA_PATTERN_96 ;
    wire \transmit_module.Y_DELTA_PATTERN_95 ;
    wire \transmit_module.Y_DELTA_PATTERN_94 ;
    wire \transmit_module.Y_DELTA_PATTERN_93 ;
    wire \transmit_module.Y_DELTA_PATTERN_83 ;
    wire \line_buffer.n593 ;
    wire \line_buffer.n585 ;
    wire \line_buffer.n3641 ;
    wire \line_buffer.n533 ;
    wire \line_buffer.n525 ;
    wire RX_DATA_7;
    wire \line_buffer.n565 ;
    wire \line_buffer.n557 ;
    wire \line_buffer.n3533 ;
    wire \line_buffer.n3549 ;
    wire \line_buffer.n3611_cascade_ ;
    wire RX_DATA_4;
    wire \tvp_video_buffer.BUFFER_1_6 ;
    wire DEBUG_c_5_c;
    wire \tvp_video_buffer.BUFFER_0_6 ;
    wire \line_buffer.n468 ;
    wire \line_buffer.n460 ;
    wire \line_buffer.n3548 ;
    wire \line_buffer.n567 ;
    wire \line_buffer.n559 ;
    wire TX_ADDR_12;
    wire \line_buffer.n3540 ;
    wire \line_buffer.n3573 ;
    wire TX_ADDR_13;
    wire \line_buffer.n3605 ;
    wire TX_DATA_4;
    wire n1814;
    wire TX_DATA_6;
    wire n1812;
    wire \transmit_module.n2385 ;
    wire \line_buffer.n470 ;
    wire \line_buffer.n462 ;
    wire \line_buffer.n3572 ;
    wire CONSTANT_ONE_NET;
    wire TVP_VIDEO_c_9;
    wire \tvp_video_buffer.BUFFER_0_9 ;
    wire \tvp_video_buffer.BUFFER_1_9 ;
    wire DEBUG_c_3_c;
    wire \transmit_module.Y_DELTA_PATTERN_88 ;
    wire \transmit_module.Y_DELTA_PATTERN_84 ;
    wire \transmit_module.Y_DELTA_PATTERN_85 ;
    wire \transmit_module.Y_DELTA_PATTERN_87 ;
    wire \transmit_module.Y_DELTA_PATTERN_86 ;
    wire ADV_CLK_c;
    wire \transmit_module.n2206 ;
    wire ADV_VSYNC_c;
    wire \line_buffer.n589 ;
    wire \line_buffer.n597 ;
    wire \line_buffer.n3534 ;
    wire TX_ADDR_11;
    wire \line_buffer.n535 ;
    wire \line_buffer.n527 ;
    wire \line_buffer.n3539 ;
    wire _gnd_net_;

    defparam \tx_pll.TX_PLL_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \tx_pll.TX_PLL_inst .TEST_MODE=1'b0;
    defparam \tx_pll.TX_PLL_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \tx_pll.TX_PLL_inst .PLLOUT_SELECT="GENCLK";
    defparam \tx_pll.TX_PLL_inst .FILTER_RANGE=3'b010;
    defparam \tx_pll.TX_PLL_inst .FEEDBACK_PATH="SIMPLE";
    defparam \tx_pll.TX_PLL_inst .FDA_RELATIVE=4'b0000;
    defparam \tx_pll.TX_PLL_inst .FDA_FEEDBACK=4'b0000;
    defparam \tx_pll.TX_PLL_inst .ENABLE_ICEGATE=1'b0;
    defparam \tx_pll.TX_PLL_inst .DIVR=4'b0000;
    defparam \tx_pll.TX_PLL_inst .DIVQ=3'b100;
    defparam \tx_pll.TX_PLL_inst .DIVF=7'b0100110;
    defparam \tx_pll.TX_PLL_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \tx_pll.TX_PLL_inst  (
            .EXTFEEDBACK(),
            .LATCHINPUTVALUE(),
            .SCLK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(ADV_CLK_c),
            .REFERENCECLK(N__18215),
            .RESETB(N__22064),
            .BYPASS(GNDG0),
            .SDI(),
            .DYNAMICDELAY({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7}),
            .PLLOUTGLOBAL());
    defparam \line_buffer.mem2_physical .WRITE_MODE=3;
    defparam \line_buffer.mem2_physical .READ_MODE=3;
    defparam \line_buffer.mem2_physical .INIT_F=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem2_physical .INIT_E=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem2_physical .INIT_D=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem2_physical .INIT_C=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem2_physical .INIT_B=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem2_physical .INIT_A=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem2_physical .INIT_9=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem2_physical .INIT_8=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem2_physical .INIT_7=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem2_physical .INIT_6=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem2_physical .INIT_5=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem2_physical .INIT_4=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem2_physical .INIT_3=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem2_physical .INIT_2=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem2_physical .INIT_1=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem2_physical .INIT_0=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    SB_RAM40_4K \line_buffer.mem2_physical  (
            .RDATA({dangling_wire_8,dangling_wire_9,dangling_wire_10,dangling_wire_11,\line_buffer.n471 ,dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,\line_buffer.n470 ,dangling_wire_19,dangling_wire_20,dangling_wire_21}),
            .RADDR({N__12593,N__10277,N__11276,N__12845,N__13319,N__10532,N__13100,N__10796,N__11048,N__10028,N__14129}),
            .WADDR({N__14939,N__17918,N__17168,N__16664,N__16916,N__19397,N__17420,N__17669,N__14402,N__15176,N__14693}),
            .MASK({dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29,dangling_wire_30,dangling_wire_31,dangling_wire_32,dangling_wire_33,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37}),
            .WDATA({dangling_wire_38,dangling_wire_39,dangling_wire_40,dangling_wire_41,N__21057,dangling_wire_42,dangling_wire_43,dangling_wire_44,dangling_wire_45,dangling_wire_46,dangling_wire_47,dangling_wire_48,N__19914,dangling_wire_49,dangling_wire_50,dangling_wire_51}),
            .RCLKE(),
            .RCLK(N__23950),
            .RE(N__22138),
            .WCLKE(),
            .WCLK(N__21988),
            .WE(N__18108));
    defparam \line_buffer.mem14_physical .WRITE_MODE=3;
    defparam \line_buffer.mem14_physical .READ_MODE=3;
    defparam \line_buffer.mem14_physical .INIT_F=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem14_physical .INIT_E=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem14_physical .INIT_D=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem14_physical .INIT_C=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem14_physical .INIT_B=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem14_physical .INIT_A=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem14_physical .INIT_9=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem14_physical .INIT_8=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem14_physical .INIT_7=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem14_physical .INIT_6=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem14_physical .INIT_5=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem14_physical .INIT_4=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem14_physical .INIT_3=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    defparam \line_buffer.mem14_physical .INIT_2=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    defparam \line_buffer.mem14_physical .INIT_1=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    defparam \line_buffer.mem14_physical .INIT_0=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    SB_RAM40_4K \line_buffer.mem14_physical  (
            .RDATA({dangling_wire_52,dangling_wire_53,dangling_wire_54,dangling_wire_55,\line_buffer.n558 ,dangling_wire_56,dangling_wire_57,dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,\line_buffer.n557 ,dangling_wire_63,dangling_wire_64,dangling_wire_65}),
            .RADDR({N__12665,N__10349,N__11348,N__12917,N__13391,N__10604,N__13172,N__10868,N__11120,N__10100,N__14201}),
            .WADDR({N__15011,N__17990,N__17240,N__16736,N__16988,N__19469,N__17492,N__17741,N__14474,N__15248,N__14765}),
            .MASK({dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73,dangling_wire_74,dangling_wire_75,dangling_wire_76,dangling_wire_77,dangling_wire_78,dangling_wire_79,dangling_wire_80,dangling_wire_81}),
            .WDATA({dangling_wire_82,dangling_wire_83,dangling_wire_84,dangling_wire_85,N__13572,dangling_wire_86,dangling_wire_87,dangling_wire_88,dangling_wire_89,dangling_wire_90,dangling_wire_91,dangling_wire_92,N__21727,dangling_wire_93,dangling_wire_94,dangling_wire_95}),
            .RCLKE(),
            .RCLK(N__24336),
            .RE(N__22211),
            .WCLKE(),
            .WCLK(N__21972),
            .WE(N__16466));
    defparam \line_buffer.mem5_physical .WRITE_MODE=3;
    defparam \line_buffer.mem5_physical .READ_MODE=3;
    defparam \line_buffer.mem5_physical .INIT_F=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem5_physical .INIT_E=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem5_physical .INIT_D=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem5_physical .INIT_C=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem5_physical .INIT_B=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem5_physical .INIT_A=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem5_physical .INIT_9=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem5_physical .INIT_8=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem5_physical .INIT_7=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem5_physical .INIT_6=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem5_physical .INIT_5=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem5_physical .INIT_4=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem5_physical .INIT_3=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    defparam \line_buffer.mem5_physical .INIT_2=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    defparam \line_buffer.mem5_physical .INIT_1=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    defparam \line_buffer.mem5_physical .INIT_0=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    SB_RAM40_4K \line_buffer.mem5_physical  (
            .RDATA({dangling_wire_96,dangling_wire_97,dangling_wire_98,dangling_wire_99,\line_buffer.n568 ,dangling_wire_100,dangling_wire_101,dangling_wire_102,dangling_wire_103,dangling_wire_104,dangling_wire_105,dangling_wire_106,\line_buffer.n567 ,dangling_wire_107,dangling_wire_108,dangling_wire_109}),
            .RADDR({N__12596,N__10274,N__11297,N__12848,N__13328,N__10523,N__13103,N__10787,N__11039,N__10043,N__14126}),
            .WADDR({N__14948,N__17927,N__17177,N__16679,N__16931,N__19412,N__17429,N__17672,N__14405,N__15185,N__14702}),
            .MASK({dangling_wire_110,dangling_wire_111,dangling_wire_112,dangling_wire_113,dangling_wire_114,dangling_wire_115,dangling_wire_116,dangling_wire_117,dangling_wire_118,dangling_wire_119,dangling_wire_120,dangling_wire_121,dangling_wire_122,dangling_wire_123,dangling_wire_124,dangling_wire_125}),
            .WDATA({dangling_wire_126,dangling_wire_127,dangling_wire_128,dangling_wire_129,N__21051,dangling_wire_130,dangling_wire_131,dangling_wire_132,dangling_wire_133,dangling_wire_134,dangling_wire_135,dangling_wire_136,N__19909,dangling_wire_137,dangling_wire_138,dangling_wire_139}),
            .RCLKE(),
            .RCLK(N__23616),
            .RE(N__22202),
            .WCLKE(),
            .WCLK(N__21986),
            .WE(N__16427));
    defparam \line_buffer.mem11_physical .WRITE_MODE=3;
    defparam \line_buffer.mem11_physical .READ_MODE=3;
    defparam \line_buffer.mem11_physical .INIT_F=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem11_physical .INIT_E=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem11_physical .INIT_D=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem11_physical .INIT_C=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem11_physical .INIT_B=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem11_physical .INIT_A=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem11_physical .INIT_9=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem11_physical .INIT_8=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem11_physical .INIT_7=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem11_physical .INIT_6=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem11_physical .INIT_5=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem11_physical .INIT_4=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem11_physical .INIT_3=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem11_physical .INIT_2=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem11_physical .INIT_1=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem11_physical .INIT_0=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    SB_RAM40_4K \line_buffer.mem11_physical  (
            .RDATA({dangling_wire_140,dangling_wire_141,dangling_wire_142,dangling_wire_143,\line_buffer.n526 ,dangling_wire_144,dangling_wire_145,dangling_wire_146,dangling_wire_147,dangling_wire_148,dangling_wire_149,dangling_wire_150,\line_buffer.n525 ,dangling_wire_151,dangling_wire_152,dangling_wire_153}),
            .RADDR({N__12701,N__10385,N__11384,N__12953,N__13427,N__10640,N__13208,N__10904,N__11156,N__10136,N__14237}),
            .WADDR({N__15047,N__18026,N__17276,N__16772,N__17024,N__19505,N__17528,N__17777,N__14510,N__15284,N__14801}),
            .MASK({dangling_wire_154,dangling_wire_155,dangling_wire_156,dangling_wire_157,dangling_wire_158,dangling_wire_159,dangling_wire_160,dangling_wire_161,dangling_wire_162,dangling_wire_163,dangling_wire_164,dangling_wire_165,dangling_wire_166,dangling_wire_167,dangling_wire_168,dangling_wire_169}),
            .WDATA({dangling_wire_170,dangling_wire_171,dangling_wire_172,dangling_wire_173,N__13571,dangling_wire_174,dangling_wire_175,dangling_wire_176,dangling_wire_177,dangling_wire_178,dangling_wire_179,dangling_wire_180,N__21738,dangling_wire_181,dangling_wire_182,dangling_wire_183}),
            .RCLKE(),
            .RCLK(N__24138),
            .RE(N__22236),
            .WCLKE(),
            .WCLK(N__21961),
            .WE(N__18725));
    defparam \line_buffer.mem21_physical .WRITE_MODE=3;
    defparam \line_buffer.mem21_physical .READ_MODE=3;
    defparam \line_buffer.mem21_physical .INIT_F=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem21_physical .INIT_E=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem21_physical .INIT_D=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem21_physical .INIT_C=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem21_physical .INIT_B=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem21_physical .INIT_A=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem21_physical .INIT_9=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem21_physical .INIT_8=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem21_physical .INIT_7=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem21_physical .INIT_6=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem21_physical .INIT_5=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem21_physical .INIT_4=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem21_physical .INIT_3=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem21_physical .INIT_2=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem21_physical .INIT_1=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem21_physical .INIT_0=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    SB_RAM40_4K \line_buffer.mem21_physical  (
            .RDATA({dangling_wire_184,dangling_wire_185,dangling_wire_186,dangling_wire_187,\line_buffer.n588 ,dangling_wire_188,dangling_wire_189,dangling_wire_190,dangling_wire_191,dangling_wire_192,dangling_wire_193,dangling_wire_194,\line_buffer.n587 ,dangling_wire_195,dangling_wire_196,dangling_wire_197}),
            .RADDR({N__12569,N__10253,N__11252,N__12821,N__13295,N__10508,N__13076,N__10772,N__11024,N__10004,N__14105}),
            .WADDR({N__14915,N__17894,N__17144,N__16640,N__16892,N__19373,N__17396,N__17645,N__14378,N__15152,N__14669}),
            .MASK({dangling_wire_198,dangling_wire_199,dangling_wire_200,dangling_wire_201,dangling_wire_202,dangling_wire_203,dangling_wire_204,dangling_wire_205,dangling_wire_206,dangling_wire_207,dangling_wire_208,dangling_wire_209,dangling_wire_210,dangling_wire_211,dangling_wire_212,dangling_wire_213}),
            .WDATA({dangling_wire_214,dangling_wire_215,dangling_wire_216,dangling_wire_217,N__15653,dangling_wire_218,dangling_wire_219,dangling_wire_220,dangling_wire_221,dangling_wire_222,dangling_wire_223,dangling_wire_224,N__9524,dangling_wire_225,dangling_wire_226,dangling_wire_227}),
            .RCLKE(),
            .RCLK(N__23811),
            .RE(N__22099),
            .WCLKE(),
            .WCLK(N__21992),
            .WE(N__18271));
    defparam \line_buffer.mem12_physical .WRITE_MODE=3;
    defparam \line_buffer.mem12_physical .READ_MODE=3;
    defparam \line_buffer.mem12_physical .INIT_F=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem12_physical .INIT_E=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem12_physical .INIT_D=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem12_physical .INIT_C=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem12_physical .INIT_B=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem12_physical .INIT_A=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem12_physical .INIT_9=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem12_physical .INIT_8=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem12_physical .INIT_7=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem12_physical .INIT_6=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem12_physical .INIT_5=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem12_physical .INIT_4=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem12_physical .INIT_3=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem12_physical .INIT_2=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem12_physical .INIT_1=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem12_physical .INIT_0=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    SB_RAM40_4K \line_buffer.mem12_physical  (
            .RDATA({dangling_wire_228,dangling_wire_229,dangling_wire_230,dangling_wire_231,\line_buffer.n524 ,dangling_wire_232,dangling_wire_233,dangling_wire_234,dangling_wire_235,dangling_wire_236,dangling_wire_237,dangling_wire_238,\line_buffer.n523 ,dangling_wire_239,dangling_wire_240,dangling_wire_241}),
            .RADDR({N__12689,N__10373,N__11372,N__12941,N__13415,N__10628,N__13196,N__10892,N__11144,N__10124,N__14225}),
            .WADDR({N__15035,N__18014,N__17264,N__16760,N__17012,N__19493,N__17516,N__17765,N__14498,N__15272,N__14789}),
            .MASK({dangling_wire_242,dangling_wire_243,dangling_wire_244,dangling_wire_245,dangling_wire_246,dangling_wire_247,dangling_wire_248,dangling_wire_249,dangling_wire_250,dangling_wire_251,dangling_wire_252,dangling_wire_253,dangling_wire_254,dangling_wire_255,dangling_wire_256,dangling_wire_257}),
            .WDATA({dangling_wire_258,dangling_wire_259,dangling_wire_260,dangling_wire_261,N__15593,dangling_wire_262,dangling_wire_263,dangling_wire_264,dangling_wire_265,dangling_wire_266,dangling_wire_267,dangling_wire_268,N__9513,dangling_wire_269,dangling_wire_270,dangling_wire_271}),
            .RCLKE(),
            .RCLK(N__24001),
            .RE(N__22235),
            .WCLKE(),
            .WCLK(N__21963),
            .WE(N__18718));
    defparam \line_buffer.mem24_physical .WRITE_MODE=3;
    defparam \line_buffer.mem24_physical .READ_MODE=3;
    defparam \line_buffer.mem24_physical .INIT_F=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem24_physical .INIT_E=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem24_physical .INIT_D=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem24_physical .INIT_C=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem24_physical .INIT_B=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem24_physical .INIT_A=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem24_physical .INIT_9=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem24_physical .INIT_8=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem24_physical .INIT_7=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem24_physical .INIT_6=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem24_physical .INIT_5=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem24_physical .INIT_4=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem24_physical .INIT_3=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem24_physical .INIT_2=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem24_physical .INIT_1=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem24_physical .INIT_0=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    SB_RAM40_4K \line_buffer.mem24_physical  (
            .RDATA({dangling_wire_272,dangling_wire_273,dangling_wire_274,dangling_wire_275,\line_buffer.n532 ,dangling_wire_276,dangling_wire_277,dangling_wire_278,dangling_wire_279,dangling_wire_280,dangling_wire_281,dangling_wire_282,\line_buffer.n531 ,dangling_wire_283,dangling_wire_284,dangling_wire_285}),
            .RADDR({N__12716,N__10394,N__11417,N__12968,N__13448,N__10643,N__13223,N__10907,N__11159,N__10163,N__14246}),
            .WADDR({N__15068,N__18047,N__17297,N__16799,N__17051,N__19532,N__17549,N__17792,N__14525,N__15305,N__14822}),
            .MASK({dangling_wire_286,dangling_wire_287,dangling_wire_288,dangling_wire_289,dangling_wire_290,dangling_wire_291,dangling_wire_292,dangling_wire_293,dangling_wire_294,dangling_wire_295,dangling_wire_296,dangling_wire_297,dangling_wire_298,dangling_wire_299,dangling_wire_300,dangling_wire_301}),
            .WDATA({dangling_wire_302,dangling_wire_303,dangling_wire_304,dangling_wire_305,N__15635,dangling_wire_306,dangling_wire_307,dangling_wire_308,dangling_wire_309,dangling_wire_310,dangling_wire_311,dangling_wire_312,N__9519,dangling_wire_313,dangling_wire_314,dangling_wire_315}),
            .RCLKE(),
            .RCLK(N__24362),
            .RE(N__22322),
            .WCLKE(),
            .WCLK(N__21950),
            .WE(N__16103));
    defparam \line_buffer.mem1_physical .WRITE_MODE=3;
    defparam \line_buffer.mem1_physical .READ_MODE=3;
    defparam \line_buffer.mem1_physical .INIT_F=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem1_physical .INIT_E=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem1_physical .INIT_D=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem1_physical .INIT_C=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem1_physical .INIT_B=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem1_physical .INIT_A=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem1_physical .INIT_9=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem1_physical .INIT_8=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem1_physical .INIT_7=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem1_physical .INIT_6=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem1_physical .INIT_5=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem1_physical .INIT_4=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem1_physical .INIT_3=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    defparam \line_buffer.mem1_physical .INIT_2=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    defparam \line_buffer.mem1_physical .INIT_1=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    defparam \line_buffer.mem1_physical .INIT_0=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    SB_RAM40_4K \line_buffer.mem1_physical  (
            .RDATA({dangling_wire_316,dangling_wire_317,dangling_wire_318,dangling_wire_319,\line_buffer.n560 ,dangling_wire_320,dangling_wire_321,dangling_wire_322,dangling_wire_323,dangling_wire_324,dangling_wire_325,dangling_wire_326,\line_buffer.n559 ,dangling_wire_327,dangling_wire_328,dangling_wire_329}),
            .RADDR({N__12725,N__10407,N__11408,N__12977,N__13451,N__10659,N__13232,N__10923,N__11175,N__10160,N__14259}),
            .WADDR({N__15071,N__18050,N__17300,N__16796,N__17048,N__19529,N__17552,N__17801,N__14534,N__15308,N__14825}),
            .MASK({dangling_wire_330,dangling_wire_331,dangling_wire_332,dangling_wire_333,dangling_wire_334,dangling_wire_335,dangling_wire_336,dangling_wire_337,dangling_wire_338,dangling_wire_339,dangling_wire_340,dangling_wire_341,dangling_wire_342,dangling_wire_343,dangling_wire_344,dangling_wire_345}),
            .WDATA({dangling_wire_346,dangling_wire_347,dangling_wire_348,dangling_wire_349,N__21029,dangling_wire_350,dangling_wire_351,dangling_wire_352,dangling_wire_353,dangling_wire_354,dangling_wire_355,dangling_wire_356,N__19922,dangling_wire_357,dangling_wire_358,dangling_wire_359}),
            .RCLKE(),
            .RCLK(N__24248),
            .RE(N__22256),
            .WCLKE(),
            .WCLK(N__21945),
            .WE(N__16473));
    defparam \line_buffer.mem15_physical .WRITE_MODE=3;
    defparam \line_buffer.mem15_physical .READ_MODE=3;
    defparam \line_buffer.mem15_physical .INIT_F=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem15_physical .INIT_E=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem15_physical .INIT_D=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem15_physical .INIT_C=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem15_physical .INIT_B=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem15_physical .INIT_A=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem15_physical .INIT_9=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem15_physical .INIT_8=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem15_physical .INIT_7=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem15_physical .INIT_6=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem15_physical .INIT_5=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem15_physical .INIT_4=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem15_physical .INIT_3=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    defparam \line_buffer.mem15_physical .INIT_2=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    defparam \line_buffer.mem15_physical .INIT_1=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    defparam \line_buffer.mem15_physical .INIT_0=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    SB_RAM40_4K \line_buffer.mem15_physical  (
            .RDATA({dangling_wire_360,dangling_wire_361,dangling_wire_362,dangling_wire_363,\line_buffer.n556 ,dangling_wire_364,dangling_wire_365,dangling_wire_366,dangling_wire_367,dangling_wire_368,dangling_wire_369,dangling_wire_370,\line_buffer.n555 ,dangling_wire_371,dangling_wire_372,dangling_wire_373}),
            .RADDR({N__12653,N__10337,N__11336,N__12905,N__13379,N__10592,N__13160,N__10856,N__11108,N__10088,N__14189}),
            .WADDR({N__14999,N__17978,N__17228,N__16724,N__16976,N__19457,N__17480,N__17729,N__14462,N__15236,N__14753}),
            .MASK({dangling_wire_374,dangling_wire_375,dangling_wire_376,dangling_wire_377,dangling_wire_378,dangling_wire_379,dangling_wire_380,dangling_wire_381,dangling_wire_382,dangling_wire_383,dangling_wire_384,dangling_wire_385,dangling_wire_386,dangling_wire_387,dangling_wire_388,dangling_wire_389}),
            .WDATA({dangling_wire_390,dangling_wire_391,dangling_wire_392,dangling_wire_393,N__15640,dangling_wire_394,dangling_wire_395,dangling_wire_396,dangling_wire_397,dangling_wire_398,dangling_wire_399,dangling_wire_400,N__9514,dangling_wire_401,dangling_wire_402,dangling_wire_403}),
            .RCLKE(),
            .RCLK(N__24114),
            .RE(N__22188),
            .WCLKE(),
            .WCLK(N__21974),
            .WE(N__16464));
    defparam \line_buffer.mem27_physical .WRITE_MODE=3;
    defparam \line_buffer.mem27_physical .READ_MODE=3;
    defparam \line_buffer.mem27_physical .INIT_F=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem27_physical .INIT_E=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem27_physical .INIT_D=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem27_physical .INIT_C=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem27_physical .INIT_B=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem27_physical .INIT_A=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem27_physical .INIT_9=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem27_physical .INIT_8=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem27_physical .INIT_7=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem27_physical .INIT_6=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem27_physical .INIT_5=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem27_physical .INIT_4=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem27_physical .INIT_3=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    defparam \line_buffer.mem27_physical .INIT_2=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    defparam \line_buffer.mem27_physical .INIT_1=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    defparam \line_buffer.mem27_physical .INIT_0=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    SB_RAM40_4K \line_buffer.mem27_physical  (
            .RDATA({dangling_wire_404,dangling_wire_405,dangling_wire_406,dangling_wire_407,\line_buffer.n564 ,dangling_wire_408,dangling_wire_409,dangling_wire_410,dangling_wire_411,dangling_wire_412,dangling_wire_413,dangling_wire_414,\line_buffer.n563 ,dangling_wire_415,dangling_wire_416,dangling_wire_417}),
            .RADDR({N__12680,N__10358,N__11381,N__12932,N__13412,N__10607,N__13187,N__10871,N__11123,N__10127,N__14210}),
            .WADDR({N__15032,N__18011,N__17261,N__16763,N__17015,N__19496,N__17513,N__17756,N__14489,N__15269,N__14786}),
            .MASK({dangling_wire_418,dangling_wire_419,dangling_wire_420,dangling_wire_421,dangling_wire_422,dangling_wire_423,dangling_wire_424,dangling_wire_425,dangling_wire_426,dangling_wire_427,dangling_wire_428,dangling_wire_429,dangling_wire_430,dangling_wire_431,dangling_wire_432,dangling_wire_433}),
            .WDATA({dangling_wire_434,dangling_wire_435,dangling_wire_436,dangling_wire_437,N__15586,dangling_wire_438,dangling_wire_439,dangling_wire_440,dangling_wire_441,dangling_wire_442,dangling_wire_443,dangling_wire_444,N__9503,dangling_wire_445,dangling_wire_446,dangling_wire_447}),
            .RCLKE(),
            .RCLK(N__24337),
            .RE(N__22297),
            .WCLKE(),
            .WCLK(N__21964),
            .WE(N__16423));
    defparam \line_buffer.mem4_physical .WRITE_MODE=3;
    defparam \line_buffer.mem4_physical .READ_MODE=3;
    defparam \line_buffer.mem4_physical .INIT_F=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem4_physical .INIT_E=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem4_physical .INIT_D=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem4_physical .INIT_C=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem4_physical .INIT_B=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem4_physical .INIT_A=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem4_physical .INIT_9=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem4_physical .INIT_8=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem4_physical .INIT_7=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem4_physical .INIT_6=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem4_physical .INIT_5=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem4_physical .INIT_4=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem4_physical .INIT_3=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem4_physical .INIT_2=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem4_physical .INIT_1=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem4_physical .INIT_0=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    SB_RAM40_4K \line_buffer.mem4_physical  (
            .RDATA({dangling_wire_448,dangling_wire_449,dangling_wire_450,dangling_wire_451,\line_buffer.n536 ,dangling_wire_452,dangling_wire_453,dangling_wire_454,dangling_wire_455,dangling_wire_456,dangling_wire_457,dangling_wire_458,\line_buffer.n535 ,dangling_wire_459,dangling_wire_460,dangling_wire_461}),
            .RADDR({N__12608,N__10286,N__11309,N__12860,N__13340,N__10535,N__13115,N__10799,N__11051,N__10055,N__14138}),
            .WADDR({N__14960,N__17939,N__17189,N__16691,N__16943,N__19424,N__17441,N__17684,N__14417,N__15197,N__14714}),
            .MASK({dangling_wire_462,dangling_wire_463,dangling_wire_464,dangling_wire_465,dangling_wire_466,dangling_wire_467,dangling_wire_468,dangling_wire_469,dangling_wire_470,dangling_wire_471,dangling_wire_472,dangling_wire_473,dangling_wire_474,dangling_wire_475,dangling_wire_476,dangling_wire_477}),
            .WDATA({dangling_wire_478,dangling_wire_479,dangling_wire_480,dangling_wire_481,N__21050,dangling_wire_482,dangling_wire_483,dangling_wire_484,dangling_wire_485,dangling_wire_486,dangling_wire_487,dangling_wire_488,N__19891,dangling_wire_489,dangling_wire_490,dangling_wire_491}),
            .RCLKE(),
            .RCLK(N__23948),
            .RE(N__22226),
            .WCLKE(),
            .WCLK(N__21984),
            .WE(N__16087));
    defparam \line_buffer.mem16_physical .WRITE_MODE=3;
    defparam \line_buffer.mem16_physical .READ_MODE=3;
    defparam \line_buffer.mem16_physical .INIT_F=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem16_physical .INIT_E=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem16_physical .INIT_D=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem16_physical .INIT_C=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem16_physical .INIT_B=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem16_physical .INIT_A=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem16_physical .INIT_9=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem16_physical .INIT_8=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem16_physical .INIT_7=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem16_physical .INIT_6=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem16_physical .INIT_5=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem16_physical .INIT_4=256'b0111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011;
    defparam \line_buffer.mem16_physical .INIT_3=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    defparam \line_buffer.mem16_physical .INIT_2=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    defparam \line_buffer.mem16_physical .INIT_1=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    defparam \line_buffer.mem16_physical .INIT_0=256'b0110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011;
    SB_RAM40_4K \line_buffer.mem16_physical  (
            .RDATA({dangling_wire_492,dangling_wire_493,dangling_wire_494,dangling_wire_495,\line_buffer.n554 ,dangling_wire_496,dangling_wire_497,dangling_wire_498,dangling_wire_499,dangling_wire_500,dangling_wire_501,dangling_wire_502,\line_buffer.n553 ,dangling_wire_503,dangling_wire_504,dangling_wire_505}),
            .RADDR({N__12641,N__10325,N__11324,N__12893,N__13367,N__10580,N__13148,N__10844,N__11096,N__10076,N__14177}),
            .WADDR({N__14987,N__17966,N__17216,N__16712,N__16964,N__19445,N__17468,N__17717,N__14450,N__15224,N__14741}),
            .MASK({dangling_wire_506,dangling_wire_507,dangling_wire_508,dangling_wire_509,dangling_wire_510,dangling_wire_511,dangling_wire_512,dangling_wire_513,dangling_wire_514,dangling_wire_515,dangling_wire_516,dangling_wire_517,dangling_wire_518,dangling_wire_519,dangling_wire_520,dangling_wire_521}),
            .WDATA({dangling_wire_522,dangling_wire_523,dangling_wire_524,dangling_wire_525,N__9312,dangling_wire_526,dangling_wire_527,dangling_wire_528,dangling_wire_529,dangling_wire_530,dangling_wire_531,dangling_wire_532,N__19134,dangling_wire_533,dangling_wire_534,dangling_wire_535}),
            .RCLKE(),
            .RCLK(N__24294),
            .RE(N__22187),
            .WCLKE(),
            .WCLK(N__21976),
            .WE(N__16465));
    defparam \line_buffer.mem30_physical .WRITE_MODE=3;
    defparam \line_buffer.mem30_physical .READ_MODE=3;
    defparam \line_buffer.mem30_physical .INIT_F=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem30_physical .INIT_E=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem30_physical .INIT_D=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem30_physical .INIT_C=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem30_physical .INIT_B=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem30_physical .INIT_A=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem30_physical .INIT_9=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem30_physical .INIT_8=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem30_physical .INIT_7=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem30_physical .INIT_6=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem30_physical .INIT_5=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem30_physical .INIT_4=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem30_physical .INIT_3=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    defparam \line_buffer.mem30_physical .INIT_2=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    defparam \line_buffer.mem30_physical .INIT_1=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    defparam \line_buffer.mem30_physical .INIT_0=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    SB_RAM40_4K \line_buffer.mem30_physical  (
            .RDATA({dangling_wire_536,dangling_wire_537,dangling_wire_538,dangling_wire_539,\line_buffer.n596 ,dangling_wire_540,dangling_wire_541,dangling_wire_542,dangling_wire_543,dangling_wire_544,dangling_wire_545,dangling_wire_546,\line_buffer.n595 ,dangling_wire_547,dangling_wire_548,dangling_wire_549}),
            .RADDR({N__12632,N__10310,N__11333,N__12884,N__13364,N__10559,N__13139,N__10823,N__11075,N__10079,N__14162}),
            .WADDR({N__14984,N__17963,N__17213,N__16715,N__16967,N__19448,N__17465,N__17708,N__14441,N__15221,N__14738}),
            .MASK({dangling_wire_550,dangling_wire_551,dangling_wire_552,dangling_wire_553,dangling_wire_554,dangling_wire_555,dangling_wire_556,dangling_wire_557,dangling_wire_558,dangling_wire_559,dangling_wire_560,dangling_wire_561,dangling_wire_562,dangling_wire_563,dangling_wire_564,dangling_wire_565}),
            .WDATA({dangling_wire_566,dangling_wire_567,dangling_wire_568,dangling_wire_569,N__15636,dangling_wire_570,dangling_wire_571,dangling_wire_572,dangling_wire_573,dangling_wire_574,dangling_wire_575,dangling_wire_576,N__9520,dangling_wire_577,dangling_wire_578,dangling_wire_579}),
            .RCLKE(),
            .RCLK(N__24204),
            .RE(N__22260),
            .WCLKE(),
            .WCLK(N__21977),
            .WE(N__16141));
    defparam \line_buffer.mem7_physical .WRITE_MODE=3;
    defparam \line_buffer.mem7_physical .READ_MODE=3;
    defparam \line_buffer.mem7_physical .INIT_F=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem7_physical .INIT_E=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem7_physical .INIT_D=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem7_physical .INIT_C=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem7_physical .INIT_B=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem7_physical .INIT_A=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem7_physical .INIT_9=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem7_physical .INIT_8=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem7_physical .INIT_7=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem7_physical .INIT_6=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem7_physical .INIT_5=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem7_physical .INIT_4=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem7_physical .INIT_3=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem7_physical .INIT_2=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem7_physical .INIT_1=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem7_physical .INIT_0=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    SB_RAM40_4K \line_buffer.mem7_physical  (
            .RDATA({dangling_wire_580,dangling_wire_581,dangling_wire_582,dangling_wire_583,\line_buffer.n463 ,dangling_wire_584,dangling_wire_585,dangling_wire_586,dangling_wire_587,dangling_wire_588,dangling_wire_589,dangling_wire_590,\line_buffer.n462 ,dangling_wire_591,dangling_wire_592,dangling_wire_593}),
            .RADDR({N__12572,N__10250,N__11273,N__12824,N__13304,N__10499,N__13079,N__10763,N__11015,N__10019,N__14102}),
            .WADDR({N__14924,N__17903,N__17153,N__16655,N__16907,N__19388,N__17405,N__17648,N__14381,N__15161,N__14678}),
            .MASK({dangling_wire_594,dangling_wire_595,dangling_wire_596,dangling_wire_597,dangling_wire_598,dangling_wire_599,dangling_wire_600,dangling_wire_601,dangling_wire_602,dangling_wire_603,dangling_wire_604,dangling_wire_605,dangling_wire_606,dangling_wire_607,dangling_wire_608,dangling_wire_609}),
            .WDATA({dangling_wire_610,dangling_wire_611,dangling_wire_612,dangling_wire_613,N__21053,dangling_wire_614,dangling_wire_615,dangling_wire_616,dangling_wire_617,dangling_wire_618,dangling_wire_619,dangling_wire_620,N__19921,dangling_wire_621,dangling_wire_622,dangling_wire_623}),
            .RCLKE(),
            .RCLK(N__23807),
            .RE(N__22154),
            .WCLKE(),
            .WCLK(N__21991),
            .WE(N__16528));
    defparam \line_buffer.mem20_physical .WRITE_MODE=3;
    defparam \line_buffer.mem20_physical .READ_MODE=3;
    defparam \line_buffer.mem20_physical .INIT_F=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem20_physical .INIT_E=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem20_physical .INIT_D=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem20_physical .INIT_C=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem20_physical .INIT_B=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem20_physical .INIT_A=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem20_physical .INIT_9=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem20_physical .INIT_8=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem20_physical .INIT_7=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem20_physical .INIT_6=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem20_physical .INIT_5=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem20_physical .INIT_4=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem20_physical .INIT_3=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem20_physical .INIT_2=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem20_physical .INIT_1=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem20_physical .INIT_0=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    SB_RAM40_4K \line_buffer.mem20_physical  (
            .RDATA({dangling_wire_624,dangling_wire_625,dangling_wire_626,dangling_wire_627,\line_buffer.n590 ,dangling_wire_628,dangling_wire_629,dangling_wire_630,dangling_wire_631,dangling_wire_632,dangling_wire_633,dangling_wire_634,\line_buffer.n589 ,dangling_wire_635,dangling_wire_636,dangling_wire_637}),
            .RADDR({N__12581,N__10265,N__11264,N__12833,N__13307,N__10520,N__13088,N__10784,N__11036,N__10016,N__14117}),
            .WADDR({N__14927,N__17906,N__17156,N__16652,N__16904,N__19385,N__17408,N__17657,N__14390,N__15164,N__14681}),
            .MASK({dangling_wire_638,dangling_wire_639,dangling_wire_640,dangling_wire_641,dangling_wire_642,dangling_wire_643,dangling_wire_644,dangling_wire_645,dangling_wire_646,dangling_wire_647,dangling_wire_648,dangling_wire_649,dangling_wire_650,dangling_wire_651,dangling_wire_652,dangling_wire_653}),
            .WDATA({dangling_wire_654,dangling_wire_655,dangling_wire_656,dangling_wire_657,N__13580,dangling_wire_658,dangling_wire_659,dangling_wire_660,dangling_wire_661,dangling_wire_662,dangling_wire_663,dangling_wire_664,N__21737,dangling_wire_665,dangling_wire_666,dangling_wire_667}),
            .RCLKE(),
            .RCLK(N__23909),
            .RE(N__22112),
            .WCLKE(),
            .WCLK(N__21990),
            .WE(N__18270));
    defparam \line_buffer.mem13_physical .WRITE_MODE=3;
    defparam \line_buffer.mem13_physical .READ_MODE=3;
    defparam \line_buffer.mem13_physical .INIT_F=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem13_physical .INIT_E=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem13_physical .INIT_D=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem13_physical .INIT_C=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem13_physical .INIT_B=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem13_physical .INIT_A=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem13_physical .INIT_9=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem13_physical .INIT_8=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem13_physical .INIT_7=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem13_physical .INIT_6=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem13_physical .INIT_5=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem13_physical .INIT_4=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem13_physical .INIT_3=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem13_physical .INIT_2=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem13_physical .INIT_1=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem13_physical .INIT_0=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    SB_RAM40_4K \line_buffer.mem13_physical  (
            .RDATA({dangling_wire_668,dangling_wire_669,dangling_wire_670,dangling_wire_671,\line_buffer.n522 ,dangling_wire_672,dangling_wire_673,dangling_wire_674,dangling_wire_675,dangling_wire_676,dangling_wire_677,dangling_wire_678,\line_buffer.n521 ,dangling_wire_679,dangling_wire_680,dangling_wire_681}),
            .RADDR({N__12677,N__10361,N__11360,N__12929,N__13403,N__10616,N__13184,N__10880,N__11132,N__10112,N__14213}),
            .WADDR({N__15023,N__18002,N__17252,N__16748,N__17000,N__19481,N__17504,N__17753,N__14486,N__15260,N__14777}),
            .MASK({dangling_wire_682,dangling_wire_683,dangling_wire_684,dangling_wire_685,dangling_wire_686,dangling_wire_687,dangling_wire_688,dangling_wire_689,dangling_wire_690,dangling_wire_691,dangling_wire_692,dangling_wire_693,dangling_wire_694,dangling_wire_695,dangling_wire_696,dangling_wire_697}),
            .WDATA({dangling_wire_698,dangling_wire_699,dangling_wire_700,dangling_wire_701,N__9311,dangling_wire_702,dangling_wire_703,dangling_wire_704,dangling_wire_705,dangling_wire_706,dangling_wire_707,dangling_wire_708,N__19119,dangling_wire_709,dangling_wire_710,dangling_wire_711}),
            .RCLKE(),
            .RCLK(N__23869),
            .RE(N__22212),
            .WCLKE(),
            .WCLK(N__21967),
            .WE(N__18717));
    defparam \line_buffer.mem19_physical .WRITE_MODE=3;
    defparam \line_buffer.mem19_physical .READ_MODE=3;
    defparam \line_buffer.mem19_physical .INIT_F=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem19_physical .INIT_E=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem19_physical .INIT_D=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem19_physical .INIT_C=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem19_physical .INIT_B=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem19_physical .INIT_A=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem19_physical .INIT_9=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem19_physical .INIT_8=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem19_physical .INIT_7=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem19_physical .INIT_6=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem19_physical .INIT_5=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem19_physical .INIT_4=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem19_physical .INIT_3=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem19_physical .INIT_2=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem19_physical .INIT_1=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem19_physical .INIT_0=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    SB_RAM40_4K \line_buffer.mem19_physical  (
            .RDATA({dangling_wire_712,dangling_wire_713,dangling_wire_714,dangling_wire_715,\line_buffer.n465 ,dangling_wire_716,dangling_wire_717,dangling_wire_718,dangling_wire_719,dangling_wire_720,dangling_wire_721,dangling_wire_722,\line_buffer.n464 ,dangling_wire_723,dangling_wire_724,dangling_wire_725}),
            .RADDR({N__12605,N__10289,N__11288,N__12857,N__13331,N__10544,N__13112,N__10808,N__11060,N__10040,N__14141}),
            .WADDR({N__14951,N__17930,N__17180,N__16676,N__16928,N__19409,N__17432,N__17681,N__14414,N__15188,N__14705}),
            .MASK({dangling_wire_726,dangling_wire_727,dangling_wire_728,dangling_wire_729,dangling_wire_730,dangling_wire_731,dangling_wire_732,dangling_wire_733,dangling_wire_734,dangling_wire_735,dangling_wire_736,dangling_wire_737,dangling_wire_738,dangling_wire_739,dangling_wire_740,dangling_wire_741}),
            .WDATA({dangling_wire_742,dangling_wire_743,dangling_wire_744,dangling_wire_745,N__9331,dangling_wire_746,dangling_wire_747,dangling_wire_748,dangling_wire_749,dangling_wire_750,dangling_wire_751,dangling_wire_752,N__19148,dangling_wire_753,dangling_wire_754,dangling_wire_755}),
            .RCLKE(),
            .RCLK(N__23735),
            .RE(N__22139),
            .WCLKE(),
            .WCLK(N__21985),
            .WE(N__18097));
    defparam \line_buffer.mem23_physical .WRITE_MODE=3;
    defparam \line_buffer.mem23_physical .READ_MODE=3;
    defparam \line_buffer.mem23_physical .INIT_F=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem23_physical .INIT_E=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem23_physical .INIT_D=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem23_physical .INIT_C=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem23_physical .INIT_B=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem23_physical .INIT_A=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem23_physical .INIT_9=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem23_physical .INIT_8=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem23_physical .INIT_7=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem23_physical .INIT_6=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem23_physical .INIT_5=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem23_physical .INIT_4=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem23_physical .INIT_3=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem23_physical .INIT_2=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem23_physical .INIT_1=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem23_physical .INIT_0=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    SB_RAM40_4K \line_buffer.mem23_physical  (
            .RDATA({dangling_wire_756,dangling_wire_757,dangling_wire_758,dangling_wire_759,\line_buffer.n534 ,dangling_wire_760,dangling_wire_761,dangling_wire_762,dangling_wire_763,dangling_wire_764,dangling_wire_765,dangling_wire_766,\line_buffer.n533 ,dangling_wire_767,dangling_wire_768,dangling_wire_769}),
            .RADDR({N__12728,N__10406,N__11424,N__12980,N__13460,N__10655,N__13235,N__10919,N__11171,N__10173,N__14258}),
            .WADDR({N__15080,N__18059,N__17309,N__16809,N__17061,N__19542,N__17561,N__17804,N__14537,N__15317,N__14834}),
            .MASK({dangling_wire_770,dangling_wire_771,dangling_wire_772,dangling_wire_773,dangling_wire_774,dangling_wire_775,dangling_wire_776,dangling_wire_777,dangling_wire_778,dangling_wire_779,dangling_wire_780,dangling_wire_781,dangling_wire_782,dangling_wire_783,dangling_wire_784,dangling_wire_785}),
            .WDATA({dangling_wire_786,dangling_wire_787,dangling_wire_788,dangling_wire_789,N__13553,dangling_wire_790,dangling_wire_791,dangling_wire_792,dangling_wire_793,dangling_wire_794,dangling_wire_795,dangling_wire_796,N__21726,dangling_wire_797,dangling_wire_798,dangling_wire_799}),
            .RCLKE(),
            .RCLK(N__24363),
            .RE(N__22326),
            .WCLKE(),
            .WCLK(N__21939),
            .WE(N__16104));
    defparam \line_buffer.mem0_physical .WRITE_MODE=3;
    defparam \line_buffer.mem0_physical .READ_MODE=3;
    defparam \line_buffer.mem0_physical .INIT_F=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem0_physical .INIT_E=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem0_physical .INIT_D=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem0_physical .INIT_C=256'b1100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110;
    defparam \line_buffer.mem0_physical .INIT_B=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem0_physical .INIT_A=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem0_physical .INIT_9=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem0_physical .INIT_8=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem0_physical .INIT_7=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem0_physical .INIT_6=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem0_physical .INIT_5=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem0_physical .INIT_4=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem0_physical .INIT_3=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem0_physical .INIT_2=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem0_physical .INIT_1=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem0_physical .INIT_0=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    SB_RAM40_4K \line_buffer.mem0_physical  (
            .RDATA({dangling_wire_800,dangling_wire_801,dangling_wire_802,dangling_wire_803,\line_buffer.n528 ,dangling_wire_804,dangling_wire_805,dangling_wire_806,dangling_wire_807,dangling_wire_808,dangling_wire_809,dangling_wire_810,\line_buffer.n527 ,dangling_wire_811,dangling_wire_812,dangling_wire_813}),
            .RADDR({N__12732,N__10413,N__11420,N__12984,N__13461,N__10665,N__13239,N__10929,N__11181,N__10172,N__14265}),
            .WADDR({N__15081,N__18060,N__17310,N__16808,N__17060,N__19541,N__17562,N__17808,N__14541,N__15318,N__14835}),
            .MASK({dangling_wire_814,dangling_wire_815,dangling_wire_816,dangling_wire_817,dangling_wire_818,dangling_wire_819,dangling_wire_820,dangling_wire_821,dangling_wire_822,dangling_wire_823,dangling_wire_824,dangling_wire_825,dangling_wire_826,dangling_wire_827,dangling_wire_828,dangling_wire_829}),
            .WDATA({dangling_wire_830,dangling_wire_831,dangling_wire_832,dangling_wire_833,N__21049,dangling_wire_834,dangling_wire_835,dangling_wire_836,dangling_wire_837,dangling_wire_838,dangling_wire_839,dangling_wire_840,N__19926,dangling_wire_841,dangling_wire_842,dangling_wire_843}),
            .RCLKE(),
            .RCLK(N__24249),
            .RE(N__22269),
            .WCLKE(),
            .WCLK(N__21934),
            .WE(N__18729));
    defparam \line_buffer.mem26_physical .WRITE_MODE=3;
    defparam \line_buffer.mem26_physical .READ_MODE=3;
    defparam \line_buffer.mem26_physical .INIT_F=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem26_physical .INIT_E=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem26_physical .INIT_D=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem26_physical .INIT_C=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem26_physical .INIT_B=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem26_physical .INIT_A=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem26_physical .INIT_9=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem26_physical .INIT_8=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem26_physical .INIT_7=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem26_physical .INIT_6=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem26_physical .INIT_5=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem26_physical .INIT_4=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem26_physical .INIT_3=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    defparam \line_buffer.mem26_physical .INIT_2=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    defparam \line_buffer.mem26_physical .INIT_1=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    defparam \line_buffer.mem26_physical .INIT_0=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    SB_RAM40_4K \line_buffer.mem26_physical  (
            .RDATA({dangling_wire_844,dangling_wire_845,dangling_wire_846,dangling_wire_847,\line_buffer.n566 ,dangling_wire_848,dangling_wire_849,dangling_wire_850,dangling_wire_851,dangling_wire_852,dangling_wire_853,dangling_wire_854,\line_buffer.n565 ,dangling_wire_855,dangling_wire_856,dangling_wire_857}),
            .RADDR({N__12692,N__10370,N__11393,N__12944,N__13424,N__10619,N__13199,N__10883,N__11135,N__10139,N__14222}),
            .WADDR({N__15044,N__18023,N__17273,N__16775,N__17027,N__19508,N__17525,N__17768,N__14501,N__15281,N__14798}),
            .MASK({dangling_wire_858,dangling_wire_859,dangling_wire_860,dangling_wire_861,dangling_wire_862,dangling_wire_863,dangling_wire_864,dangling_wire_865,dangling_wire_866,dangling_wire_867,dangling_wire_868,dangling_wire_869,dangling_wire_870,dangling_wire_871,dangling_wire_872,dangling_wire_873}),
            .WDATA({dangling_wire_874,dangling_wire_875,dangling_wire_876,dangling_wire_877,N__13570,dangling_wire_878,dangling_wire_879,dangling_wire_880,dangling_wire_881,dangling_wire_882,dangling_wire_883,dangling_wire_884,N__21724,dangling_wire_885,dangling_wire_886,dangling_wire_887}),
            .RCLKE(),
            .RCLK(N__24354),
            .RE(N__22306),
            .WCLKE(),
            .WCLK(N__21962),
            .WE(N__16428));
    defparam \line_buffer.mem3_physical .WRITE_MODE=3;
    defparam \line_buffer.mem3_physical .READ_MODE=3;
    defparam \line_buffer.mem3_physical .INIT_F=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem3_physical .INIT_E=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem3_physical .INIT_D=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem3_physical .INIT_C=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem3_physical .INIT_B=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem3_physical .INIT_A=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem3_physical .INIT_9=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem3_physical .INIT_8=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem3_physical .INIT_7=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem3_physical .INIT_6=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem3_physical .INIT_5=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem3_physical .INIT_4=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem3_physical .INIT_3=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem3_physical .INIT_2=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem3_physical .INIT_1=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem3_physical .INIT_0=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    SB_RAM40_4K \line_buffer.mem3_physical  (
            .RDATA({dangling_wire_888,dangling_wire_889,dangling_wire_890,dangling_wire_891,\line_buffer.n592 ,dangling_wire_892,dangling_wire_893,dangling_wire_894,dangling_wire_895,dangling_wire_896,dangling_wire_897,dangling_wire_898,\line_buffer.n591 ,dangling_wire_899,dangling_wire_900,dangling_wire_901}),
            .RADDR({N__12644,N__10322,N__11345,N__12896,N__13376,N__10571,N__13151,N__10835,N__11087,N__10091,N__14174}),
            .WADDR({N__14996,N__17975,N__17225,N__16727,N__16979,N__19460,N__17477,N__17720,N__14453,N__15233,N__14750}),
            .MASK({dangling_wire_902,dangling_wire_903,dangling_wire_904,dangling_wire_905,dangling_wire_906,dangling_wire_907,dangling_wire_908,dangling_wire_909,dangling_wire_910,dangling_wire_911,dangling_wire_912,dangling_wire_913,dangling_wire_914,dangling_wire_915,dangling_wire_916,dangling_wire_917}),
            .WDATA({dangling_wire_918,dangling_wire_919,dangling_wire_920,dangling_wire_921,N__21033,dangling_wire_922,dangling_wire_923,dangling_wire_924,dangling_wire_925,dangling_wire_926,dangling_wire_927,dangling_wire_928,N__19874,dangling_wire_929,dangling_wire_930,dangling_wire_931}),
            .RCLKE(),
            .RCLK(N__24293),
            .RE(N__22270),
            .WCLKE(),
            .WCLK(N__21975),
            .WE(N__18275));
    defparam \line_buffer.mem17_physical .WRITE_MODE=3;
    defparam \line_buffer.mem17_physical .READ_MODE=3;
    defparam \line_buffer.mem17_physical .INIT_F=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem17_physical .INIT_E=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem17_physical .INIT_D=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem17_physical .INIT_C=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem17_physical .INIT_B=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem17_physical .INIT_A=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem17_physical .INIT_9=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem17_physical .INIT_8=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem17_physical .INIT_7=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem17_physical .INIT_6=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem17_physical .INIT_5=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem17_physical .INIT_4=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem17_physical .INIT_3=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem17_physical .INIT_2=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem17_physical .INIT_1=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem17_physical .INIT_0=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    SB_RAM40_4K \line_buffer.mem17_physical  (
            .RDATA({dangling_wire_932,dangling_wire_933,dangling_wire_934,dangling_wire_935,\line_buffer.n469 ,dangling_wire_936,dangling_wire_937,dangling_wire_938,dangling_wire_939,dangling_wire_940,dangling_wire_941,dangling_wire_942,\line_buffer.n468 ,dangling_wire_943,dangling_wire_944,dangling_wire_945}),
            .RADDR({N__12629,N__10313,N__11312,N__12881,N__13355,N__10568,N__13136,N__10832,N__11084,N__10064,N__14165}),
            .WADDR({N__14975,N__17954,N__17204,N__16700,N__16952,N__19433,N__17456,N__17705,N__14438,N__15212,N__14729}),
            .MASK({dangling_wire_946,dangling_wire_947,dangling_wire_948,dangling_wire_949,dangling_wire_950,dangling_wire_951,dangling_wire_952,dangling_wire_953,dangling_wire_954,dangling_wire_955,dangling_wire_956,dangling_wire_957,dangling_wire_958,dangling_wire_959,dangling_wire_960,dangling_wire_961}),
            .WDATA({dangling_wire_962,dangling_wire_963,dangling_wire_964,dangling_wire_965,N__13573,dangling_wire_966,dangling_wire_967,dangling_wire_968,dangling_wire_969,dangling_wire_970,dangling_wire_971,dangling_wire_972,N__21714,dangling_wire_973,dangling_wire_974,dangling_wire_975}),
            .RCLKE(),
            .RCLK(N__23980),
            .RE(N__22164),
            .WCLKE(),
            .WCLK(N__21981),
            .WE(N__18091));
    defparam \line_buffer.mem31_physical .WRITE_MODE=3;
    defparam \line_buffer.mem31_physical .READ_MODE=3;
    defparam \line_buffer.mem31_physical .INIT_F=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem31_physical .INIT_E=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem31_physical .INIT_D=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem31_physical .INIT_C=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem31_physical .INIT_B=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem31_physical .INIT_A=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem31_physical .INIT_9=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem31_physical .INIT_8=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem31_physical .INIT_7=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem31_physical .INIT_6=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem31_physical .INIT_5=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem31_physical .INIT_4=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem31_physical .INIT_3=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    defparam \line_buffer.mem31_physical .INIT_2=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    defparam \line_buffer.mem31_physical .INIT_1=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    defparam \line_buffer.mem31_physical .INIT_0=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    SB_RAM40_4K \line_buffer.mem31_physical  (
            .RDATA({dangling_wire_976,dangling_wire_977,dangling_wire_978,dangling_wire_979,\line_buffer.n594 ,dangling_wire_980,dangling_wire_981,dangling_wire_982,dangling_wire_983,dangling_wire_984,dangling_wire_985,dangling_wire_986,\line_buffer.n593 ,dangling_wire_987,dangling_wire_988,dangling_wire_989}),
            .RADDR({N__12620,N__10298,N__11321,N__12872,N__13352,N__10547,N__13127,N__10811,N__11063,N__10067,N__14150}),
            .WADDR({N__14972,N__17951,N__17201,N__16703,N__16955,N__19436,N__17453,N__17696,N__14429,N__15209,N__14726}),
            .MASK({dangling_wire_990,dangling_wire_991,dangling_wire_992,dangling_wire_993,dangling_wire_994,dangling_wire_995,dangling_wire_996,dangling_wire_997,dangling_wire_998,dangling_wire_999,dangling_wire_1000,dangling_wire_1001,dangling_wire_1002,dangling_wire_1003,dangling_wire_1004,dangling_wire_1005}),
            .WDATA({dangling_wire_1006,dangling_wire_1007,dangling_wire_1008,dangling_wire_1009,N__9335,dangling_wire_1010,dangling_wire_1011,dangling_wire_1012,dangling_wire_1013,dangling_wire_1014,dangling_wire_1015,dangling_wire_1016,N__19133,dangling_wire_1017,dangling_wire_1018,dangling_wire_1019}),
            .RCLKE(),
            .RCLK(N__23979),
            .RE(N__22246),
            .WCLKE(),
            .WCLK(N__21982),
            .WE(N__16148));
    defparam \line_buffer.mem9_physical .INIT_0=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem9_physical .WRITE_MODE=3;
    defparam \line_buffer.mem9_physical .READ_MODE=3;
    defparam \line_buffer.mem9_physical .INIT_F=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem9_physical .INIT_E=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem9_physical .INIT_D=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem9_physical .INIT_C=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem9_physical .INIT_B=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem9_physical .INIT_A=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem9_physical .INIT_9=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem9_physical .INIT_8=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem9_physical .INIT_7=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem9_physical .INIT_6=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem9_physical .INIT_5=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem9_physical .INIT_4=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem9_physical .INIT_3=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem9_physical .INIT_2=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem9_physical .INIT_1=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    SB_RAM40_4K \line_buffer.mem9_physical  (
            .RDATA({dangling_wire_1020,dangling_wire_1021,dangling_wire_1022,dangling_wire_1023,\line_buffer.n459 ,dangling_wire_1024,dangling_wire_1025,dangling_wire_1026,dangling_wire_1027,dangling_wire_1028,dangling_wire_1029,dangling_wire_1030,\line_buffer.n458 ,dangling_wire_1031,dangling_wire_1032,dangling_wire_1033}),
            .RADDR({N__12548,N__10226,N__11249,N__12800,N__13280,N__10475,N__13055,N__10739,N__10991,N__9995,N__14078}),
            .WADDR({N__14900,N__17879,N__17129,N__16631,N__16883,N__19364,N__17381,N__17624,N__14357,N__15137,N__14654}),
            .MASK({dangling_wire_1034,dangling_wire_1035,dangling_wire_1036,dangling_wire_1037,dangling_wire_1038,dangling_wire_1039,dangling_wire_1040,dangling_wire_1041,dangling_wire_1042,dangling_wire_1043,dangling_wire_1044,dangling_wire_1045,dangling_wire_1046,dangling_wire_1047,dangling_wire_1048,dangling_wire_1049}),
            .WDATA({dangling_wire_1050,dangling_wire_1051,dangling_wire_1052,dangling_wire_1053,N__15657,dangling_wire_1054,dangling_wire_1055,dangling_wire_1056,dangling_wire_1057,dangling_wire_1058,dangling_wire_1059,dangling_wire_1060,N__9534,dangling_wire_1061,dangling_wire_1062,dangling_wire_1063}),
            .RCLKE(),
            .RCLK(N__23643),
            .RE(N__22153),
            .WCLKE(),
            .WCLK(N__21995),
            .WE(N__16532));
    defparam \line_buffer.mem29_physical .WRITE_MODE=3;
    defparam \line_buffer.mem29_physical .READ_MODE=3;
    defparam \line_buffer.mem29_physical .INIT_F=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem29_physical .INIT_E=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem29_physical .INIT_D=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem29_physical .INIT_C=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem29_physical .INIT_B=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem29_physical .INIT_A=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem29_physical .INIT_9=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem29_physical .INIT_8=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem29_physical .INIT_7=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem29_physical .INIT_6=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem29_physical .INIT_5=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem29_physical .INIT_4=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem29_physical .INIT_3=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    defparam \line_buffer.mem29_physical .INIT_2=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    defparam \line_buffer.mem29_physical .INIT_1=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    defparam \line_buffer.mem29_physical .INIT_0=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    SB_RAM40_4K \line_buffer.mem29_physical  (
            .RDATA({dangling_wire_1064,dangling_wire_1065,dangling_wire_1066,dangling_wire_1067,\line_buffer.n598 ,dangling_wire_1068,dangling_wire_1069,dangling_wire_1070,dangling_wire_1071,dangling_wire_1072,dangling_wire_1073,dangling_wire_1074,\line_buffer.n597 ,dangling_wire_1075,dangling_wire_1076,dangling_wire_1077}),
            .RADDR({N__12656,N__10334,N__11357,N__12908,N__13388,N__10583,N__13163,N__10847,N__11099,N__10103,N__14186}),
            .WADDR({N__15008,N__17987,N__17237,N__16739,N__16991,N__19472,N__17489,N__17732,N__14465,N__15245,N__14762}),
            .MASK({dangling_wire_1078,dangling_wire_1079,dangling_wire_1080,dangling_wire_1081,dangling_wire_1082,dangling_wire_1083,dangling_wire_1084,dangling_wire_1085,dangling_wire_1086,dangling_wire_1087,dangling_wire_1088,dangling_wire_1089,dangling_wire_1090,dangling_wire_1091,dangling_wire_1092,dangling_wire_1093}),
            .WDATA({dangling_wire_1094,dangling_wire_1095,dangling_wire_1096,dangling_wire_1097,N__13554,dangling_wire_1098,dangling_wire_1099,dangling_wire_1100,dangling_wire_1101,dangling_wire_1102,dangling_wire_1103,dangling_wire_1104,N__21704,dangling_wire_1105,dangling_wire_1106,dangling_wire_1107}),
            .RCLKE(),
            .RCLK(N__24313),
            .RE(N__22279),
            .WCLKE(),
            .WCLK(N__21973),
            .WE(N__16140));
    defparam \line_buffer.mem6_physical .WRITE_MODE=3;
    defparam \line_buffer.mem6_physical .READ_MODE=3;
    defparam \line_buffer.mem6_physical .INIT_F=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem6_physical .INIT_E=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem6_physical .INIT_D=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem6_physical .INIT_C=256'b1111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011111100110111001111110011011100111111001101110011;
    defparam \line_buffer.mem6_physical .INIT_B=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem6_physical .INIT_A=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem6_physical .INIT_9=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem6_physical .INIT_8=256'b1110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011111000110110001111100011011000111110001101100011;
    defparam \line_buffer.mem6_physical .INIT_7=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem6_physical .INIT_6=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem6_physical .INIT_5=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem6_physical .INIT_4=256'b1110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111111001110110011111100111011001111110011101100111;
    defparam \line_buffer.mem6_physical .INIT_3=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    defparam \line_buffer.mem6_physical .INIT_2=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    defparam \line_buffer.mem6_physical .INIT_1=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    defparam \line_buffer.mem6_physical .INIT_0=256'b1110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110111001100110011011100110011001101110011001100110;
    SB_RAM40_4K \line_buffer.mem6_physical  (
            .RDATA({dangling_wire_1108,dangling_wire_1109,dangling_wire_1110,dangling_wire_1111,\line_buffer.n600 ,dangling_wire_1112,dangling_wire_1113,dangling_wire_1114,dangling_wire_1115,dangling_wire_1116,dangling_wire_1117,dangling_wire_1118,\line_buffer.n599 ,dangling_wire_1119,dangling_wire_1120,dangling_wire_1121}),
            .RADDR({N__12584,N__10262,N__11285,N__12836,N__13316,N__10511,N__13091,N__10775,N__11027,N__10031,N__14114}),
            .WADDR({N__14936,N__17915,N__17165,N__16667,N__16919,N__19400,N__17417,N__17660,N__14393,N__15173,N__14690}),
            .MASK({dangling_wire_1122,dangling_wire_1123,dangling_wire_1124,dangling_wire_1125,dangling_wire_1126,dangling_wire_1127,dangling_wire_1128,dangling_wire_1129,dangling_wire_1130,dangling_wire_1131,dangling_wire_1132,dangling_wire_1133,dangling_wire_1134,dangling_wire_1135,dangling_wire_1136,dangling_wire_1137}),
            .WDATA({dangling_wire_1138,dangling_wire_1139,dangling_wire_1140,dangling_wire_1141,N__21052,dangling_wire_1142,dangling_wire_1143,dangling_wire_1144,dangling_wire_1145,dangling_wire_1146,dangling_wire_1147,dangling_wire_1148,N__19910,dangling_wire_1149,dangling_wire_1150,dangling_wire_1151}),
            .RCLKE(),
            .RCLK(N__23949),
            .RE(N__22178),
            .WCLKE(),
            .WCLK(N__21989),
            .WE(N__16152));
    defparam \line_buffer.mem10_physical .WRITE_MODE=3;
    defparam \line_buffer.mem10_physical .READ_MODE=3;
    defparam \line_buffer.mem10_physical .INIT_F=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem10_physical .INIT_E=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem10_physical .INIT_D=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem10_physical .INIT_C=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem10_physical .INIT_B=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem10_physical .INIT_A=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem10_physical .INIT_9=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem10_physical .INIT_8=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem10_physical .INIT_7=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem10_physical .INIT_6=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem10_physical .INIT_5=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem10_physical .INIT_4=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem10_physical .INIT_3=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem10_physical .INIT_2=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem10_physical .INIT_1=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem10_physical .INIT_0=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    SB_RAM40_4K \line_buffer.mem10_physical  (
            .RDATA({dangling_wire_1152,dangling_wire_1153,dangling_wire_1154,dangling_wire_1155,\line_buffer.n457 ,dangling_wire_1156,dangling_wire_1157,dangling_wire_1158,dangling_wire_1159,dangling_wire_1160,dangling_wire_1161,dangling_wire_1162,\line_buffer.n456 ,dangling_wire_1163,dangling_wire_1164,dangling_wire_1165}),
            .RADDR({N__12713,N__10397,N__11396,N__12965,N__13439,N__10652,N__13220,N__10916,N__11168,N__10148,N__14249}),
            .WADDR({N__15059,N__18038,N__17288,N__16784,N__17036,N__19517,N__17540,N__17789,N__14522,N__15296,N__14813}),
            .MASK({dangling_wire_1166,dangling_wire_1167,dangling_wire_1168,dangling_wire_1169,dangling_wire_1170,dangling_wire_1171,dangling_wire_1172,dangling_wire_1173,dangling_wire_1174,dangling_wire_1175,dangling_wire_1176,dangling_wire_1177,dangling_wire_1178,dangling_wire_1179,dangling_wire_1180,dangling_wire_1181}),
            .WDATA({dangling_wire_1182,dangling_wire_1183,dangling_wire_1184,dangling_wire_1185,N__9310,dangling_wire_1186,dangling_wire_1187,dangling_wire_1188,dangling_wire_1189,dangling_wire_1190,dangling_wire_1191,dangling_wire_1192,N__19140,dangling_wire_1193,dangling_wire_1194,dangling_wire_1195}),
            .RCLKE(),
            .RCLK(N__24139),
            .RE(N__22255),
            .WCLKE(),
            .WCLK(N__21954),
            .WE(N__16533));
    defparam \line_buffer.mem22_physical .INIT_0=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem22_physical .WRITE_MODE=3;
    defparam \line_buffer.mem22_physical .READ_MODE=3;
    defparam \line_buffer.mem22_physical .INIT_F=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem22_physical .INIT_E=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem22_physical .INIT_D=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem22_physical .INIT_C=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem22_physical .INIT_B=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem22_physical .INIT_A=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem22_physical .INIT_9=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem22_physical .INIT_8=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem22_physical .INIT_7=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem22_physical .INIT_6=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem22_physical .INIT_5=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem22_physical .INIT_4=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem22_physical .INIT_3=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem22_physical .INIT_2=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    defparam \line_buffer.mem22_physical .INIT_1=256'b0011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011;
    SB_RAM40_4K \line_buffer.mem22_physical  (
            .RDATA({dangling_wire_1196,dangling_wire_1197,dangling_wire_1198,dangling_wire_1199,\line_buffer.n586 ,dangling_wire_1200,dangling_wire_1201,dangling_wire_1202,dangling_wire_1203,dangling_wire_1204,dangling_wire_1205,dangling_wire_1206,\line_buffer.n585 ,dangling_wire_1207,dangling_wire_1208,dangling_wire_1209}),
            .RADDR({N__12557,N__10241,N__11240,N__12809,N__13283,N__10496,N__13064,N__10760,N__11012,N__9992,N__14093}),
            .WADDR({N__14903,N__17882,N__17132,N__16628,N__16880,N__19361,N__17384,N__17633,N__14366,N__15140,N__14657}),
            .MASK({dangling_wire_1210,dangling_wire_1211,dangling_wire_1212,dangling_wire_1213,dangling_wire_1214,dangling_wire_1215,dangling_wire_1216,dangling_wire_1217,dangling_wire_1218,dangling_wire_1219,dangling_wire_1220,dangling_wire_1221,dangling_wire_1222,dangling_wire_1223,dangling_wire_1224,dangling_wire_1225}),
            .WDATA({dangling_wire_1226,dangling_wire_1227,dangling_wire_1228,dangling_wire_1229,N__9339,dangling_wire_1230,dangling_wire_1231,dangling_wire_1232,dangling_wire_1233,dangling_wire_1234,dangling_wire_1235,dangling_wire_1236,N__19155,dangling_wire_1237,dangling_wire_1238,dangling_wire_1239}),
            .RCLKE(),
            .RCLK(N__23764),
            .RE(N__22111),
            .WCLKE(),
            .WCLK(N__21994),
            .WE(N__18276));
    defparam \line_buffer.mem25_physical .WRITE_MODE=3;
    defparam \line_buffer.mem25_physical .READ_MODE=3;
    defparam \line_buffer.mem25_physical .INIT_F=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem25_physical .INIT_E=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem25_physical .INIT_D=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem25_physical .INIT_C=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem25_physical .INIT_B=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem25_physical .INIT_A=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem25_physical .INIT_9=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem25_physical .INIT_8=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem25_physical .INIT_7=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem25_physical .INIT_6=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem25_physical .INIT_5=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem25_physical .INIT_4=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem25_physical .INIT_3=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem25_physical .INIT_2=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem25_physical .INIT_1=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem25_physical .INIT_0=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    SB_RAM40_4K \line_buffer.mem25_physical  (
            .RDATA({dangling_wire_1240,dangling_wire_1241,dangling_wire_1242,dangling_wire_1243,\line_buffer.n530 ,dangling_wire_1244,dangling_wire_1245,dangling_wire_1246,dangling_wire_1247,dangling_wire_1248,dangling_wire_1249,dangling_wire_1250,\line_buffer.n529 ,dangling_wire_1251,dangling_wire_1252,dangling_wire_1253}),
            .RADDR({N__12704,N__10382,N__11405,N__12956,N__13436,N__10631,N__13211,N__10895,N__11147,N__10151,N__14234}),
            .WADDR({N__15056,N__18035,N__17285,N__16787,N__17039,N__19520,N__17537,N__17780,N__14513,N__15293,N__14810}),
            .MASK({dangling_wire_1254,dangling_wire_1255,dangling_wire_1256,dangling_wire_1257,dangling_wire_1258,dangling_wire_1259,dangling_wire_1260,dangling_wire_1261,dangling_wire_1262,dangling_wire_1263,dangling_wire_1264,dangling_wire_1265,dangling_wire_1266,dangling_wire_1267,dangling_wire_1268,dangling_wire_1269}),
            .WDATA({dangling_wire_1270,dangling_wire_1271,dangling_wire_1272,dangling_wire_1273,N__9303,dangling_wire_1274,dangling_wire_1275,dangling_wire_1276,dangling_wire_1277,dangling_wire_1278,dangling_wire_1279,dangling_wire_1280,N__19141,dangling_wire_1281,dangling_wire_1282,dangling_wire_1283}),
            .RCLKE(),
            .RCLK(N__24355),
            .RE(N__22315),
            .WCLKE(),
            .WCLK(N__21956),
            .WE(N__16096));
    defparam \line_buffer.mem8_physical .WRITE_MODE=3;
    defparam \line_buffer.mem8_physical .READ_MODE=3;
    defparam \line_buffer.mem8_physical .INIT_F=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem8_physical .INIT_E=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem8_physical .INIT_D=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem8_physical .INIT_C=256'b1100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100;
    defparam \line_buffer.mem8_physical .INIT_B=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem8_physical .INIT_A=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem8_physical .INIT_9=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem8_physical .INIT_8=256'b1000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100;
    defparam \line_buffer.mem8_physical .INIT_7=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem8_physical .INIT_6=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem8_physical .INIT_5=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem8_physical .INIT_4=256'b1001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100;
    defparam \line_buffer.mem8_physical .INIT_3=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem8_physical .INIT_2=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem8_physical .INIT_1=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    defparam \line_buffer.mem8_physical .INIT_0=256'b1001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000;
    SB_RAM40_4K \line_buffer.mem8_physical  (
            .RDATA({dangling_wire_1284,dangling_wire_1285,dangling_wire_1286,dangling_wire_1287,\line_buffer.n461 ,dangling_wire_1288,dangling_wire_1289,dangling_wire_1290,dangling_wire_1291,dangling_wire_1292,dangling_wire_1293,dangling_wire_1294,\line_buffer.n460 ,dangling_wire_1295,dangling_wire_1296,dangling_wire_1297}),
            .RADDR({N__12560,N__10238,N__11261,N__12812,N__13292,N__10487,N__13067,N__10751,N__11003,N__10007,N__14090}),
            .WADDR({N__14912,N__17891,N__17141,N__16643,N__16895,N__19376,N__17393,N__17636,N__14369,N__15149,N__14666}),
            .MASK({dangling_wire_1298,dangling_wire_1299,dangling_wire_1300,dangling_wire_1301,dangling_wire_1302,dangling_wire_1303,dangling_wire_1304,dangling_wire_1305,dangling_wire_1306,dangling_wire_1307,dangling_wire_1308,dangling_wire_1309,dangling_wire_1310,dangling_wire_1311,dangling_wire_1312,dangling_wire_1313}),
            .WDATA({dangling_wire_1314,dangling_wire_1315,dangling_wire_1316,dangling_wire_1317,N__13581,dangling_wire_1318,dangling_wire_1319,dangling_wire_1320,dangling_wire_1321,dangling_wire_1322,dangling_wire_1323,dangling_wire_1324,N__21725,dangling_wire_1325,dangling_wire_1326,dangling_wire_1327}),
            .RCLKE(),
            .RCLK(N__23681),
            .RE(N__22126),
            .WCLKE(),
            .WCLK(N__21993),
            .WE(N__16527));
    defparam \line_buffer.mem28_physical .WRITE_MODE=3;
    defparam \line_buffer.mem28_physical .READ_MODE=3;
    defparam \line_buffer.mem28_physical .INIT_F=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem28_physical .INIT_E=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem28_physical .INIT_D=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem28_physical .INIT_C=256'b0110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111011001110110011101100111;
    defparam \line_buffer.mem28_physical .INIT_B=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem28_physical .INIT_A=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem28_physical .INIT_9=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem28_physical .INIT_8=256'b0110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110;
    defparam \line_buffer.mem28_physical .INIT_7=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem28_physical .INIT_6=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem28_physical .INIT_5=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem28_physical .INIT_4=256'b1110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110111001101110011011100110;
    defparam \line_buffer.mem28_physical .INIT_3=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    defparam \line_buffer.mem28_physical .INIT_2=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    defparam \line_buffer.mem28_physical .INIT_1=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    defparam \line_buffer.mem28_physical .INIT_0=256'b1100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110110001101100011011000110;
    SB_RAM40_4K \line_buffer.mem28_physical  (
            .RDATA({dangling_wire_1328,dangling_wire_1329,dangling_wire_1330,dangling_wire_1331,\line_buffer.n562 ,dangling_wire_1332,dangling_wire_1333,dangling_wire_1334,dangling_wire_1335,dangling_wire_1336,dangling_wire_1337,dangling_wire_1338,\line_buffer.n561 ,dangling_wire_1339,dangling_wire_1340,dangling_wire_1341}),
            .RADDR({N__12668,N__10346,N__11369,N__12920,N__13400,N__10595,N__13175,N__10859,N__11111,N__10115,N__14198}),
            .WADDR({N__15020,N__17999,N__17249,N__16751,N__17003,N__19484,N__17501,N__17744,N__14477,N__15257,N__14774}),
            .MASK({dangling_wire_1342,dangling_wire_1343,dangling_wire_1344,dangling_wire_1345,dangling_wire_1346,dangling_wire_1347,dangling_wire_1348,dangling_wire_1349,dangling_wire_1350,dangling_wire_1351,dangling_wire_1352,dangling_wire_1353,dangling_wire_1354,dangling_wire_1355,dangling_wire_1356,dangling_wire_1357}),
            .WDATA({dangling_wire_1358,dangling_wire_1359,dangling_wire_1360,dangling_wire_1361,N__9318,dangling_wire_1362,dangling_wire_1363,dangling_wire_1364,dangling_wire_1365,dangling_wire_1366,dangling_wire_1367,dangling_wire_1368,N__19129,dangling_wire_1369,dangling_wire_1370,dangling_wire_1371}),
            .RCLKE(),
            .RCLK(N__23745),
            .RE(N__22288),
            .WCLKE(),
            .WCLK(N__21970),
            .WE(N__16413));
    defparam \line_buffer.mem18_physical .WRITE_MODE=3;
    defparam \line_buffer.mem18_physical .READ_MODE=3;
    defparam \line_buffer.mem18_physical .INIT_F=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem18_physical .INIT_E=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem18_physical .INIT_D=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem18_physical .INIT_C=256'b1001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011001;
    defparam \line_buffer.mem18_physical .INIT_B=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem18_physical .INIT_A=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem18_physical .INIT_9=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem18_physical .INIT_8=256'b0001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001000110010001100100011001;
    defparam \line_buffer.mem18_physical .INIT_7=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem18_physical .INIT_6=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem18_physical .INIT_5=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem18_physical .INIT_4=256'b0011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001001110010011100100111001;
    defparam \line_buffer.mem18_physical .INIT_3=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem18_physical .INIT_2=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem18_physical .INIT_1=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    defparam \line_buffer.mem18_physical .INIT_0=256'b0011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001001100010011000100110001;
    SB_RAM40_4K \line_buffer.mem18_physical  (
            .RDATA({dangling_wire_1372,dangling_wire_1373,dangling_wire_1374,dangling_wire_1375,\line_buffer.n467 ,dangling_wire_1376,dangling_wire_1377,dangling_wire_1378,dangling_wire_1379,dangling_wire_1380,dangling_wire_1381,dangling_wire_1382,\line_buffer.n466 ,dangling_wire_1383,dangling_wire_1384,dangling_wire_1385}),
            .RADDR({N__12617,N__10301,N__11300,N__12869,N__13343,N__10556,N__13124,N__10820,N__11072,N__10052,N__14153}),
            .WADDR({N__14963,N__17942,N__17192,N__16688,N__16940,N__19421,N__17444,N__17693,N__14426,N__15200,N__14717}),
            .MASK({dangling_wire_1386,dangling_wire_1387,dangling_wire_1388,dangling_wire_1389,dangling_wire_1390,dangling_wire_1391,dangling_wire_1392,dangling_wire_1393,dangling_wire_1394,dangling_wire_1395,dangling_wire_1396,dangling_wire_1397,dangling_wire_1398,dangling_wire_1399,dangling_wire_1400,dangling_wire_1401}),
            .WDATA({dangling_wire_1402,dangling_wire_1403,dangling_wire_1404,dangling_wire_1405,N__15631,dangling_wire_1406,dangling_wire_1407,dangling_wire_1408,dangling_wire_1409,dangling_wire_1410,dangling_wire_1411,dangling_wire_1412,N__9515,dangling_wire_1413,dangling_wire_1414,dangling_wire_1415}),
            .RCLKE(),
            .RCLK(N__24065),
            .RE(N__22163),
            .WCLKE(),
            .WCLK(N__21983),
            .WE(N__18104));
    PRE_IO_GBUF DEBUG_c_3_pad_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__24832),
            .GLOBALBUFFEROUTPUT(DEBUG_c_3_c));
    defparam DEBUG_c_3_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_c_3_pad_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_c_3_pad_iopad (
            .OE(N__24834),
            .DIN(N__24833),
            .DOUT(N__24832),
            .PACKAGEPIN(TVP_CLK));
    defparam DEBUG_c_3_pad_preio.PIN_TYPE=6'b000001;
    defparam DEBUG_c_3_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_c_3_pad_preio (
            .PADOEN(N__24834),
            .PADOUT(N__24833),
            .PADIN(N__24832),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_CLK_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_CLK_pad_iopad.PULLUP=1'b0;
    IO_PAD ADV_CLK_pad_iopad (
            .OE(N__24823),
            .DIN(N__24822),
            .DOUT(N__24821),
            .PACKAGEPIN(ADV_CLK));
    defparam ADV_CLK_pad_preio.PIN_TYPE=6'b011001;
    defparam ADV_CLK_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_CLK_pad_preio (
            .PADOEN(N__24823),
            .PADOUT(N__24822),
            .PADIN(N__24821),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__24064),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_c_2_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_c_2_pad_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_c_2_pad_iopad (
            .OE(N__24814),
            .DIN(N__24813),
            .DOUT(N__24812),
            .PACKAGEPIN(TVP_HSYNC));
    defparam DEBUG_c_2_pad_preio.PIN_TYPE=6'b000001;
    defparam DEBUG_c_2_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_c_2_pad_preio (
            .PADOEN(N__24814),
            .PADOUT(N__24813),
            .PADIN(N__24812),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DEBUG_c_2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_3_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_3_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_3_iopad (
            .OE(N__24805),
            .DIN(N__24804),
            .DOUT(N__24803),
            .PACKAGEPIN(DEBUG[3]));
    defparam DEBUG_pad_3_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_3_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_3_preio (
            .PADOEN(N__24805),
            .PADOUT(N__24804),
            .PADIN(N__24803),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__18225),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_VIDEO_pad_2_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_VIDEO_pad_2_iopad.PULLUP=1'b1;
    IO_PAD TVP_VIDEO_pad_2_iopad (
            .OE(N__24796),
            .DIN(N__24795),
            .DOUT(N__24794),
            .PACKAGEPIN(TVP_VIDEO[2]));
    defparam TVP_VIDEO_pad_2_preio.PIN_TYPE=6'b000001;
    defparam TVP_VIDEO_pad_2_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_VIDEO_pad_2_preio (
            .PADOEN(N__24796),
            .PADOUT(N__24795),
            .PADIN(N__24794),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_VIDEO_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_5_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_5_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_5_iopad (
            .OE(N__24787),
            .DIN(N__24786),
            .DOUT(N__24785),
            .PACKAGEPIN(ADV_G[5]));
    defparam ADV_G_pad_5_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_5_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_5_preio (
            .PADOEN(N__24787),
            .PADOUT(N__24786),
            .PADIN(N__24785),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__20762),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_3_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_3_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_3_iopad (
            .OE(N__24778),
            .DIN(N__24777),
            .DOUT(N__24776),
            .PACKAGEPIN(ADV_R[3]));
    defparam ADV_R_pad_3_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_3_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_3_preio (
            .PADOEN(N__24778),
            .PADOUT(N__24777),
            .PADIN(N__24776),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__18337),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_0_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_0_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_0_iopad (
            .OE(N__24769),
            .DIN(N__24768),
            .DOUT(N__24767),
            .PACKAGEPIN(ADV_R[0]));
    defparam ADV_R_pad_0_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_0_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_0_preio (
            .PADOEN(N__24769),
            .PADOUT(N__24768),
            .PADIN(N__24767),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__14598),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_2_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_2_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_2_iopad (
            .OE(N__24760),
            .DIN(N__24759),
            .DOUT(N__24758),
            .PACKAGEPIN(DEBUG[2]));
    defparam DEBUG_pad_2_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_2_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_2_preio (
            .PADOEN(N__24760),
            .PADOUT(N__24759),
            .PADIN(N__24758),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__20181),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_VIDEO_pad_3_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_VIDEO_pad_3_iopad.PULLUP=1'b1;
    IO_PAD TVP_VIDEO_pad_3_iopad (
            .OE(N__24751),
            .DIN(N__24750),
            .DOUT(N__24749),
            .PACKAGEPIN(TVP_VIDEO[3]));
    defparam TVP_VIDEO_pad_3_preio.PIN_TYPE=6'b000001;
    defparam TVP_VIDEO_pad_3_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_VIDEO_pad_3_preio (
            .PADOEN(N__24751),
            .PADOUT(N__24750),
            .PADIN(N__24749),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_VIDEO_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_4_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_4_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_4_iopad (
            .OE(N__24742),
            .DIN(N__24741),
            .DOUT(N__24740),
            .PACKAGEPIN(ADV_G[4]));
    defparam ADV_G_pad_4_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_4_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_4_preio (
            .PADOEN(N__24742),
            .PADOUT(N__24741),
            .PADIN(N__24740),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__22548),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_5_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_5_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_5_iopad (
            .OE(N__24733),
            .DIN(N__24732),
            .DOUT(N__24731),
            .PACKAGEPIN(ADV_R[5]));
    defparam ADV_R_pad_5_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_5_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_5_preio (
            .PADOEN(N__24733),
            .PADOUT(N__24732),
            .PADIN(N__24731),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__20766),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_VIDEO_pad_9_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_VIDEO_pad_9_iopad.PULLUP=1'b1;
    IO_PAD TVP_VIDEO_pad_9_iopad (
            .OE(N__24724),
            .DIN(N__24723),
            .DOUT(N__24722),
            .PACKAGEPIN(TVP_VIDEO[9]));
    defparam TVP_VIDEO_pad_9_preio.PIN_TYPE=6'b000001;
    defparam TVP_VIDEO_pad_9_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_VIDEO_pad_9_preio (
            .PADOEN(N__24724),
            .PADOUT(N__24723),
            .PADIN(N__24722),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_VIDEO_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_1_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_1_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_1_iopad (
            .OE(N__24715),
            .DIN(N__24714),
            .DOUT(N__24713),
            .PACKAGEPIN(DEBUG[1]));
    defparam DEBUG_pad_1_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_1_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_1_preio (
            .PADOEN(N__24715),
            .PADOUT(N__24714),
            .PADIN(N__24713),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__13623),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_c_6_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_c_6_pad_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_c_6_pad_iopad (
            .OE(N__24706),
            .DIN(N__24705),
            .DOUT(N__24704),
            .PACKAGEPIN(TVP_VIDEO[7]));
    defparam DEBUG_c_6_pad_preio.PIN_TYPE=6'b000001;
    defparam DEBUG_c_6_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_c_6_pad_preio (
            .PADOEN(N__24706),
            .PADOUT(N__24705),
            .PADIN(N__24704),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DEBUG_c_6_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_1_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_1_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_1_iopad (
            .OE(N__24697),
            .DIN(N__24696),
            .DOUT(N__24695),
            .PACKAGEPIN(ADV_B[1]));
    defparam ADV_B_pad_1_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_1_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_1_preio (
            .PADOEN(N__24697),
            .PADOUT(N__24696),
            .PADIN(N__24695),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__20678),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_SYNC_N_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_SYNC_N_pad_iopad.PULLUP=1'b1;
    IO_PAD ADV_SYNC_N_pad_iopad (
            .OE(N__24688),
            .DIN(N__24687),
            .DOUT(N__24686),
            .PACKAGEPIN(ADV_SYNC_N));
    defparam ADV_SYNC_N_pad_preio.PIN_TYPE=6'b011001;
    defparam ADV_SYNC_N_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_SYNC_N_pad_preio (
            .PADOEN(N__24688),
            .PADOUT(N__24687),
            .PADIN(N__24686),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_6_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_6_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_6_iopad (
            .OE(N__24679),
            .DIN(N__24678),
            .DOUT(N__24677),
            .PACKAGEPIN(ADV_B[6]));
    defparam ADV_B_pad_6_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_6_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_6_preio (
            .PADOEN(N__24679),
            .PADOUT(N__24678),
            .PADIN(N__24677),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__22481),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_6_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_6_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_6_iopad (
            .OE(N__24670),
            .DIN(N__24669),
            .DOUT(N__24668),
            .PACKAGEPIN(DEBUG[6]));
    defparam DEBUG_pad_6_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_6_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_6_preio (
            .PADOEN(N__24670),
            .PADOUT(N__24669),
            .PADIN(N__24668),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9240),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_0_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_0_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_0_iopad (
            .OE(N__24661),
            .DIN(N__24660),
            .DOUT(N__24659),
            .PACKAGEPIN(ADV_G[0]));
    defparam ADV_G_pad_0_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_0_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_0_preio (
            .PADOEN(N__24661),
            .PADOUT(N__24660),
            .PADIN(N__24659),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__14597),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_1_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_1_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_1_iopad (
            .OE(N__24652),
            .DIN(N__24651),
            .DOUT(N__24650),
            .PACKAGEPIN(ADV_R[1]));
    defparam ADV_R_pad_1_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_1_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_1_preio (
            .PADOEN(N__24652),
            .PADOUT(N__24651),
            .PADIN(N__24650),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__20696),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_5_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_5_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_5_iopad (
            .OE(N__24643),
            .DIN(N__24642),
            .DOUT(N__24641),
            .PACKAGEPIN(DEBUG[5]));
    defparam DEBUG_pad_5_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_5_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_5_preio (
            .PADOEN(N__24643),
            .PADOUT(N__24642),
            .PADIN(N__24641),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__21627),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_7_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_7_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_7_iopad (
            .OE(N__24634),
            .DIN(N__24633),
            .DOUT(N__24632),
            .PACKAGEPIN(ADV_G[7]));
    defparam ADV_G_pad_7_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_7_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_7_preio (
            .PADOEN(N__24634),
            .PADOUT(N__24633),
            .PADIN(N__24632),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11519),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_6_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_6_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_6_iopad (
            .OE(N__24625),
            .DIN(N__24624),
            .DOUT(N__24623),
            .PACKAGEPIN(ADV_R[6]));
    defparam ADV_R_pad_6_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_6_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_6_preio (
            .PADOEN(N__24625),
            .PADOUT(N__24624),
            .PADIN(N__24623),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__22488),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_BLANK_N_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_BLANK_N_pad_iopad.PULLUP=1'b1;
    IO_PAD ADV_BLANK_N_pad_iopad (
            .OE(N__24616),
            .DIN(N__24615),
            .DOUT(N__24614),
            .PACKAGEPIN(ADV_BLANK_N));
    defparam ADV_BLANK_N_pad_preio.PIN_TYPE=6'b011001;
    defparam ADV_BLANK_N_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_BLANK_N_pad_preio (
            .PADOEN(N__24616),
            .PADOUT(N__24615),
            .PADIN(N__24614),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__22060),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_0_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_0_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_0_iopad (
            .OE(N__24607),
            .DIN(N__24606),
            .DOUT(N__24605),
            .PACKAGEPIN(DEBUG[0]));
    defparam DEBUG_pad_0_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_0_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_0_preio (
            .PADOEN(N__24607),
            .PADOUT(N__24606),
            .PADIN(N__24605),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__18186),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_2_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_2_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_2_iopad (
            .OE(N__24598),
            .DIN(N__24597),
            .DOUT(N__24596),
            .PACKAGEPIN(ADV_B[2]));
    defparam ADV_B_pad_2_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_2_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_2_preio (
            .PADOEN(N__24598),
            .PADOUT(N__24597),
            .PADIN(N__24596),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9419),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_c_7_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_c_7_pad_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_c_7_pad_iopad (
            .OE(N__24589),
            .DIN(N__24588),
            .DOUT(N__24587),
            .PACKAGEPIN(TVP_VIDEO[8]));
    defparam DEBUG_c_7_pad_preio.PIN_TYPE=6'b000001;
    defparam DEBUG_c_7_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_c_7_pad_preio (
            .PADOEN(N__24589),
            .PADOUT(N__24588),
            .PADIN(N__24587),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DEBUG_c_7_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_c_1_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_c_1_pad_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_c_1_pad_iopad (
            .OE(N__24580),
            .DIN(N__24579),
            .DOUT(N__24578),
            .PACKAGEPIN(TVP_VSYNC));
    defparam DEBUG_c_1_pad_preio.PIN_TYPE=6'b000001;
    defparam DEBUG_c_1_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_c_1_pad_preio (
            .PADOEN(N__24580),
            .PADOUT(N__24579),
            .PADIN(N__24578),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DEBUG_c_1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_c_5_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_c_5_pad_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_c_5_pad_iopad (
            .OE(N__24571),
            .DIN(N__24570),
            .DOUT(N__24569),
            .PACKAGEPIN(TVP_VIDEO[6]));
    defparam DEBUG_c_5_pad_preio.PIN_TYPE=6'b000001;
    defparam DEBUG_c_5_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_c_5_pad_preio (
            .PADOEN(N__24571),
            .PADOUT(N__24570),
            .PADIN(N__24569),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(DEBUG_c_5_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_7_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_7_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_7_iopad (
            .OE(N__24562),
            .DIN(N__24561),
            .DOUT(N__24560),
            .PACKAGEPIN(ADV_B[7]));
    defparam ADV_B_pad_7_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_7_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_7_preio (
            .PADOEN(N__24562),
            .PADOUT(N__24561),
            .PADIN(N__24560),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11518),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam LED_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam LED_pad_iopad.PULLUP=1'b1;
    IO_PAD LED_pad_iopad (
            .OE(N__24553),
            .DIN(N__24552),
            .DOUT(N__24551),
            .PACKAGEPIN(LED));
    defparam LED_pad_preio.PIN_TYPE=6'b011001;
    defparam LED_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO LED_pad_preio (
            .PADOEN(N__24553),
            .PADOUT(N__24552),
            .PADIN(N__24551),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__18147),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_VIDEO_pad_4_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_VIDEO_pad_4_iopad.PULLUP=1'b1;
    IO_PAD TVP_VIDEO_pad_4_iopad (
            .OE(N__24544),
            .DIN(N__24543),
            .DOUT(N__24542),
            .PACKAGEPIN(TVP_VIDEO[4]));
    defparam TVP_VIDEO_pad_4_preio.PIN_TYPE=6'b000001;
    defparam TVP_VIDEO_pad_4_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_VIDEO_pad_4_preio (
            .PADOEN(N__24544),
            .PADOUT(N__24543),
            .PADIN(N__24542),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_VIDEO_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_3_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_3_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_3_iopad (
            .OE(N__24535),
            .DIN(N__24534),
            .DOUT(N__24533),
            .PACKAGEPIN(ADV_G[3]));
    defparam ADV_G_pad_3_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_3_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_3_preio (
            .PADOEN(N__24535),
            .PADOUT(N__24534),
            .PADIN(N__24533),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__18339),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_HSYNC_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_HSYNC_pad_iopad.PULLUP=1'b0;
    IO_PAD ADV_HSYNC_pad_iopad (
            .OE(N__24526),
            .DIN(N__24525),
            .DOUT(N__24524),
            .PACKAGEPIN(ADV_HSYNC));
    defparam ADV_HSYNC_pad_preio.PIN_TYPE=6'b011001;
    defparam ADV_HSYNC_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_HSYNC_pad_preio (
            .PADOEN(N__24526),
            .PADOUT(N__24525),
            .PADIN(N__24524),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11832),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_2_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_2_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_2_iopad (
            .OE(N__24517),
            .DIN(N__24516),
            .DOUT(N__24515),
            .PACKAGEPIN(ADV_R[2]));
    defparam ADV_R_pad_2_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_2_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_2_preio (
            .PADOEN(N__24517),
            .PADOUT(N__24516),
            .PADIN(N__24515),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9400),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_4_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_4_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_4_iopad (
            .OE(N__24508),
            .DIN(N__24507),
            .DOUT(N__24506),
            .PACKAGEPIN(ADV_B[4]));
    defparam ADV_B_pad_4_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_4_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_4_preio (
            .PADOEN(N__24508),
            .PADOUT(N__24507),
            .PADIN(N__24506),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__22531),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_4_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_4_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_4_iopad (
            .OE(N__24499),
            .DIN(N__24498),
            .DOUT(N__24497),
            .PACKAGEPIN(DEBUG[4]));
    defparam DEBUG_pad_4_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_4_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_4_preio (
            .PADOEN(N__24499),
            .PADOUT(N__24498),
            .PADIN(N__24497),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__19701),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_6_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_6_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_6_iopad (
            .OE(N__24490),
            .DIN(N__24489),
            .DOUT(N__24488),
            .PACKAGEPIN(ADV_G[6]));
    defparam ADV_G_pad_6_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_6_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_6_preio (
            .PADOEN(N__24490),
            .PADOUT(N__24489),
            .PADIN(N__24488),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__22477),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_7_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_7_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_7_iopad (
            .OE(N__24481),
            .DIN(N__24480),
            .DOUT(N__24479),
            .PACKAGEPIN(ADV_R[7]));
    defparam ADV_R_pad_7_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_7_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_7_preio (
            .PADOEN(N__24481),
            .PADOUT(N__24480),
            .PADIN(N__24479),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__11520),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_3_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_3_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_3_iopad (
            .OE(N__24472),
            .DIN(N__24471),
            .DOUT(N__24470),
            .PACKAGEPIN(ADV_B[3]));
    defparam ADV_B_pad_3_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_3_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_3_preio (
            .PADOEN(N__24472),
            .PADOUT(N__24471),
            .PADIN(N__24470),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__18338),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_4_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_4_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_4_iopad (
            .OE(N__24463),
            .DIN(N__24462),
            .DOUT(N__24461),
            .PACKAGEPIN(ADV_R[4]));
    defparam ADV_R_pad_4_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_4_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_4_preio (
            .PADOEN(N__24463),
            .PADOUT(N__24462),
            .PADIN(N__24461),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__22538),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_0_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_0_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_0_iopad (
            .OE(N__24454),
            .DIN(N__24453),
            .DOUT(N__24452),
            .PACKAGEPIN(ADV_B[0]));
    defparam ADV_B_pad_0_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_0_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_0_preio (
            .PADOEN(N__24454),
            .PADOUT(N__24453),
            .PADIN(N__24452),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__14593),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_VIDEO_pad_5_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_VIDEO_pad_5_iopad.PULLUP=1'b1;
    IO_PAD TVP_VIDEO_pad_5_iopad (
            .OE(N__24445),
            .DIN(N__24444),
            .DOUT(N__24443),
            .PACKAGEPIN(TVP_VIDEO[5]));
    defparam TVP_VIDEO_pad_5_preio.PIN_TYPE=6'b000001;
    defparam TVP_VIDEO_pad_5_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_VIDEO_pad_5_preio (
            .PADOEN(N__24445),
            .PADOUT(N__24444),
            .PADIN(N__24443),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_VIDEO_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_2_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_2_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_2_iopad (
            .OE(N__24436),
            .DIN(N__24435),
            .DOUT(N__24434),
            .PACKAGEPIN(ADV_G[2]));
    defparam ADV_G_pad_2_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_2_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_2_preio (
            .PADOEN(N__24436),
            .PADOUT(N__24435),
            .PADIN(N__24434),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9420),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_VSYNC_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_VSYNC_pad_iopad.PULLUP=1'b0;
    IO_PAD ADV_VSYNC_pad_iopad (
            .OE(N__24427),
            .DIN(N__24426),
            .DOUT(N__24425),
            .PACKAGEPIN(ADV_VSYNC));
    defparam ADV_VSYNC_pad_preio.PIN_TYPE=6'b011001;
    defparam ADV_VSYNC_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_VSYNC_pad_preio (
            .PADOEN(N__24427),
            .PADOUT(N__24426),
            .PADIN(N__24425),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__23346),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_5_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_5_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_5_iopad (
            .OE(N__24418),
            .DIN(N__24417),
            .DOUT(N__24416),
            .PACKAGEPIN(ADV_B[5]));
    defparam ADV_B_pad_5_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_5_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_5_preio (
            .PADOEN(N__24418),
            .PADOUT(N__24417),
            .PADIN(N__24416),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__20743),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_7_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_7_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_7_iopad (
            .OE(N__24409),
            .DIN(N__24408),
            .DOUT(N__24407),
            .PACKAGEPIN(DEBUG[7]));
    defparam DEBUG_pad_7_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_7_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_7_preio (
            .PADOEN(N__24409),
            .PADOUT(N__24408),
            .PADIN(N__24407),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__19965),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_1_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_1_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_1_iopad (
            .OE(N__24400),
            .DIN(N__24399),
            .DOUT(N__24398),
            .PACKAGEPIN(ADV_G[1]));
    defparam ADV_G_pad_1_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_1_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_1_preio (
            .PADOEN(N__24400),
            .PADOUT(N__24399),
            .PADIN(N__24398),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__20700),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__5856 (
            .O(N__24381),
            .I(N__24378));
    LocalMux I__5855 (
            .O(N__24378),
            .I(\transmit_module.Y_DELTA_PATTERN_85 ));
    InMux I__5854 (
            .O(N__24375),
            .I(N__24372));
    LocalMux I__5853 (
            .O(N__24372),
            .I(\transmit_module.Y_DELTA_PATTERN_87 ));
    InMux I__5852 (
            .O(N__24369),
            .I(N__24366));
    LocalMux I__5851 (
            .O(N__24366),
            .I(\transmit_module.Y_DELTA_PATTERN_86 ));
    ClkMux I__5850 (
            .O(N__24363),
            .I(N__24359));
    ClkMux I__5849 (
            .O(N__24362),
            .I(N__24356));
    LocalMux I__5848 (
            .O(N__24359),
            .I(N__24344));
    LocalMux I__5847 (
            .O(N__24356),
            .I(N__24344));
    ClkMux I__5846 (
            .O(N__24355),
            .I(N__24341));
    ClkMux I__5845 (
            .O(N__24354),
            .I(N__24338));
    ClkMux I__5844 (
            .O(N__24353),
            .I(N__24328));
    ClkMux I__5843 (
            .O(N__24352),
            .I(N__24325));
    ClkMux I__5842 (
            .O(N__24351),
            .I(N__24322));
    ClkMux I__5841 (
            .O(N__24350),
            .I(N__24319));
    ClkMux I__5840 (
            .O(N__24349),
            .I(N__24316));
    Span4Mux_s2_v I__5839 (
            .O(N__24344),
            .I(N__24305));
    LocalMux I__5838 (
            .O(N__24341),
            .I(N__24305));
    LocalMux I__5837 (
            .O(N__24338),
            .I(N__24305));
    ClkMux I__5836 (
            .O(N__24337),
            .I(N__24302));
    ClkMux I__5835 (
            .O(N__24336),
            .I(N__24296));
    ClkMux I__5834 (
            .O(N__24335),
            .I(N__24288));
    ClkMux I__5833 (
            .O(N__24334),
            .I(N__24284));
    ClkMux I__5832 (
            .O(N__24333),
            .I(N__24280));
    ClkMux I__5831 (
            .O(N__24332),
            .I(N__24277));
    ClkMux I__5830 (
            .O(N__24331),
            .I(N__24274));
    LocalMux I__5829 (
            .O(N__24328),
            .I(N__24267));
    LocalMux I__5828 (
            .O(N__24325),
            .I(N__24258));
    LocalMux I__5827 (
            .O(N__24322),
            .I(N__24258));
    LocalMux I__5826 (
            .O(N__24319),
            .I(N__24258));
    LocalMux I__5825 (
            .O(N__24316),
            .I(N__24258));
    ClkMux I__5824 (
            .O(N__24315),
            .I(N__24255));
    ClkMux I__5823 (
            .O(N__24314),
            .I(N__24252));
    ClkMux I__5822 (
            .O(N__24313),
            .I(N__24245));
    ClkMux I__5821 (
            .O(N__24312),
            .I(N__24242));
    Span4Mux_v I__5820 (
            .O(N__24305),
            .I(N__24236));
    LocalMux I__5819 (
            .O(N__24302),
            .I(N__24236));
    ClkMux I__5818 (
            .O(N__24301),
            .I(N__24233));
    ClkMux I__5817 (
            .O(N__24300),
            .I(N__24230));
    ClkMux I__5816 (
            .O(N__24299),
            .I(N__24224));
    LocalMux I__5815 (
            .O(N__24296),
            .I(N__24217));
    ClkMux I__5814 (
            .O(N__24295),
            .I(N__24214));
    ClkMux I__5813 (
            .O(N__24294),
            .I(N__24210));
    ClkMux I__5812 (
            .O(N__24293),
            .I(N__24205));
    ClkMux I__5811 (
            .O(N__24292),
            .I(N__24201));
    ClkMux I__5810 (
            .O(N__24291),
            .I(N__24198));
    LocalMux I__5809 (
            .O(N__24288),
            .I(N__24194));
    ClkMux I__5808 (
            .O(N__24287),
            .I(N__24191));
    LocalMux I__5807 (
            .O(N__24284),
            .I(N__24188));
    ClkMux I__5806 (
            .O(N__24283),
            .I(N__24185));
    LocalMux I__5805 (
            .O(N__24280),
            .I(N__24181));
    LocalMux I__5804 (
            .O(N__24277),
            .I(N__24176));
    LocalMux I__5803 (
            .O(N__24274),
            .I(N__24176));
    ClkMux I__5802 (
            .O(N__24273),
            .I(N__24173));
    ClkMux I__5801 (
            .O(N__24272),
            .I(N__24170));
    ClkMux I__5800 (
            .O(N__24271),
            .I(N__24167));
    ClkMux I__5799 (
            .O(N__24270),
            .I(N__24164));
    Span4Mux_v I__5798 (
            .O(N__24267),
            .I(N__24159));
    Span4Mux_v I__5797 (
            .O(N__24258),
            .I(N__24159));
    LocalMux I__5796 (
            .O(N__24255),
            .I(N__24156));
    LocalMux I__5795 (
            .O(N__24252),
            .I(N__24153));
    ClkMux I__5794 (
            .O(N__24251),
            .I(N__24150));
    ClkMux I__5793 (
            .O(N__24250),
            .I(N__24147));
    ClkMux I__5792 (
            .O(N__24249),
            .I(N__24143));
    ClkMux I__5791 (
            .O(N__24248),
            .I(N__24140));
    LocalMux I__5790 (
            .O(N__24245),
            .I(N__24133));
    LocalMux I__5789 (
            .O(N__24242),
            .I(N__24133));
    ClkMux I__5788 (
            .O(N__24241),
            .I(N__24130));
    Span4Mux_v I__5787 (
            .O(N__24236),
            .I(N__24125));
    LocalMux I__5786 (
            .O(N__24233),
            .I(N__24125));
    LocalMux I__5785 (
            .O(N__24230),
            .I(N__24122));
    ClkMux I__5784 (
            .O(N__24229),
            .I(N__24119));
    ClkMux I__5783 (
            .O(N__24228),
            .I(N__24116));
    ClkMux I__5782 (
            .O(N__24227),
            .I(N__24109));
    LocalMux I__5781 (
            .O(N__24224),
            .I(N__24106));
    ClkMux I__5780 (
            .O(N__24223),
            .I(N__24103));
    ClkMux I__5779 (
            .O(N__24222),
            .I(N__24099));
    ClkMux I__5778 (
            .O(N__24221),
            .I(N__24096));
    ClkMux I__5777 (
            .O(N__24220),
            .I(N__24093));
    Span4Mux_h I__5776 (
            .O(N__24217),
            .I(N__24087));
    LocalMux I__5775 (
            .O(N__24214),
            .I(N__24087));
    ClkMux I__5774 (
            .O(N__24213),
            .I(N__24084));
    LocalMux I__5773 (
            .O(N__24210),
            .I(N__24081));
    ClkMux I__5772 (
            .O(N__24209),
            .I(N__24078));
    ClkMux I__5771 (
            .O(N__24208),
            .I(N__24075));
    LocalMux I__5770 (
            .O(N__24205),
            .I(N__24071));
    ClkMux I__5769 (
            .O(N__24204),
            .I(N__24068));
    LocalMux I__5768 (
            .O(N__24201),
            .I(N__24061));
    LocalMux I__5767 (
            .O(N__24198),
            .I(N__24058));
    ClkMux I__5766 (
            .O(N__24197),
            .I(N__24055));
    Span4Mux_v I__5765 (
            .O(N__24194),
            .I(N__24050));
    LocalMux I__5764 (
            .O(N__24191),
            .I(N__24050));
    Span4Mux_h I__5763 (
            .O(N__24188),
            .I(N__24045));
    LocalMux I__5762 (
            .O(N__24185),
            .I(N__24045));
    ClkMux I__5761 (
            .O(N__24184),
            .I(N__24042));
    Span4Mux_v I__5760 (
            .O(N__24181),
            .I(N__24033));
    Span4Mux_h I__5759 (
            .O(N__24176),
            .I(N__24033));
    LocalMux I__5758 (
            .O(N__24173),
            .I(N__24033));
    LocalMux I__5757 (
            .O(N__24170),
            .I(N__24033));
    LocalMux I__5756 (
            .O(N__24167),
            .I(N__24028));
    LocalMux I__5755 (
            .O(N__24164),
            .I(N__24028));
    Span4Mux_h I__5754 (
            .O(N__24159),
            .I(N__24017));
    Span4Mux_h I__5753 (
            .O(N__24156),
            .I(N__24017));
    Span4Mux_v I__5752 (
            .O(N__24153),
            .I(N__24017));
    LocalMux I__5751 (
            .O(N__24150),
            .I(N__24017));
    LocalMux I__5750 (
            .O(N__24147),
            .I(N__24017));
    ClkMux I__5749 (
            .O(N__24146),
            .I(N__24014));
    LocalMux I__5748 (
            .O(N__24143),
            .I(N__24011));
    LocalMux I__5747 (
            .O(N__24140),
            .I(N__24008));
    ClkMux I__5746 (
            .O(N__24139),
            .I(N__24005));
    ClkMux I__5745 (
            .O(N__24138),
            .I(N__24002));
    Span4Mux_v I__5744 (
            .O(N__24133),
            .I(N__23996));
    LocalMux I__5743 (
            .O(N__24130),
            .I(N__23996));
    Span4Mux_h I__5742 (
            .O(N__24125),
            .I(N__23987));
    Span4Mux_v I__5741 (
            .O(N__24122),
            .I(N__23987));
    LocalMux I__5740 (
            .O(N__24119),
            .I(N__23987));
    LocalMux I__5739 (
            .O(N__24116),
            .I(N__23987));
    ClkMux I__5738 (
            .O(N__24115),
            .I(N__23984));
    ClkMux I__5737 (
            .O(N__24114),
            .I(N__23981));
    ClkMux I__5736 (
            .O(N__24113),
            .I(N__23974));
    ClkMux I__5735 (
            .O(N__24112),
            .I(N__23969));
    LocalMux I__5734 (
            .O(N__24109),
            .I(N__23966));
    Span4Mux_h I__5733 (
            .O(N__24106),
            .I(N__23961));
    LocalMux I__5732 (
            .O(N__24103),
            .I(N__23961));
    ClkMux I__5731 (
            .O(N__24102),
            .I(N__23958));
    LocalMux I__5730 (
            .O(N__24099),
            .I(N__23952));
    LocalMux I__5729 (
            .O(N__24096),
            .I(N__23952));
    LocalMux I__5728 (
            .O(N__24093),
            .I(N__23945));
    ClkMux I__5727 (
            .O(N__24092),
            .I(N__23942));
    Span4Mux_h I__5726 (
            .O(N__24087),
            .I(N__23937));
    LocalMux I__5725 (
            .O(N__24084),
            .I(N__23937));
    Span4Mux_h I__5724 (
            .O(N__24081),
            .I(N__23934));
    LocalMux I__5723 (
            .O(N__24078),
            .I(N__23931));
    LocalMux I__5722 (
            .O(N__24075),
            .I(N__23928));
    ClkMux I__5721 (
            .O(N__24074),
            .I(N__23925));
    Span4Mux_v I__5720 (
            .O(N__24071),
            .I(N__23920));
    LocalMux I__5719 (
            .O(N__24068),
            .I(N__23920));
    ClkMux I__5718 (
            .O(N__24067),
            .I(N__23917));
    ClkMux I__5717 (
            .O(N__24066),
            .I(N__23914));
    ClkMux I__5716 (
            .O(N__24065),
            .I(N__23911));
    IoInMux I__5715 (
            .O(N__24064),
            .I(N__23906));
    Span4Mux_v I__5714 (
            .O(N__24061),
            .I(N__23899));
    Span4Mux_v I__5713 (
            .O(N__24058),
            .I(N__23899));
    LocalMux I__5712 (
            .O(N__24055),
            .I(N__23899));
    Span4Mux_h I__5711 (
            .O(N__24050),
            .I(N__23892));
    Span4Mux_v I__5710 (
            .O(N__24045),
            .I(N__23892));
    LocalMux I__5709 (
            .O(N__24042),
            .I(N__23892));
    Span4Mux_v I__5708 (
            .O(N__24033),
            .I(N__23883));
    Span4Mux_h I__5707 (
            .O(N__24028),
            .I(N__23883));
    Span4Mux_h I__5706 (
            .O(N__24017),
            .I(N__23883));
    LocalMux I__5705 (
            .O(N__24014),
            .I(N__23883));
    Span4Mux_s2_v I__5704 (
            .O(N__24011),
            .I(N__23876));
    Span4Mux_h I__5703 (
            .O(N__24008),
            .I(N__23876));
    LocalMux I__5702 (
            .O(N__24005),
            .I(N__23876));
    LocalMux I__5701 (
            .O(N__24002),
            .I(N__23873));
    ClkMux I__5700 (
            .O(N__24001),
            .I(N__23870));
    Span4Mux_h I__5699 (
            .O(N__23996),
            .I(N__23862));
    Span4Mux_v I__5698 (
            .O(N__23987),
            .I(N__23862));
    LocalMux I__5697 (
            .O(N__23984),
            .I(N__23862));
    LocalMux I__5696 (
            .O(N__23981),
            .I(N__23859));
    ClkMux I__5695 (
            .O(N__23980),
            .I(N__23856));
    ClkMux I__5694 (
            .O(N__23979),
            .I(N__23853));
    ClkMux I__5693 (
            .O(N__23978),
            .I(N__23849));
    ClkMux I__5692 (
            .O(N__23977),
            .I(N__23846));
    LocalMux I__5691 (
            .O(N__23974),
            .I(N__23842));
    ClkMux I__5690 (
            .O(N__23973),
            .I(N__23839));
    ClkMux I__5689 (
            .O(N__23972),
            .I(N__23836));
    LocalMux I__5688 (
            .O(N__23969),
            .I(N__23832));
    Span4Mux_h I__5687 (
            .O(N__23966),
            .I(N__23825));
    Span4Mux_h I__5686 (
            .O(N__23961),
            .I(N__23825));
    LocalMux I__5685 (
            .O(N__23958),
            .I(N__23825));
    ClkMux I__5684 (
            .O(N__23957),
            .I(N__23822));
    Span4Mux_v I__5683 (
            .O(N__23952),
            .I(N__23819));
    ClkMux I__5682 (
            .O(N__23951),
            .I(N__23816));
    ClkMux I__5681 (
            .O(N__23950),
            .I(N__23812));
    ClkMux I__5680 (
            .O(N__23949),
            .I(N__23808));
    ClkMux I__5679 (
            .O(N__23948),
            .I(N__23804));
    Span4Mux_h I__5678 (
            .O(N__23945),
            .I(N__23799));
    LocalMux I__5677 (
            .O(N__23942),
            .I(N__23799));
    Span4Mux_h I__5676 (
            .O(N__23937),
            .I(N__23795));
    Span4Mux_h I__5675 (
            .O(N__23934),
            .I(N__23786));
    Span4Mux_v I__5674 (
            .O(N__23931),
            .I(N__23786));
    Span4Mux_h I__5673 (
            .O(N__23928),
            .I(N__23786));
    LocalMux I__5672 (
            .O(N__23925),
            .I(N__23786));
    Span4Mux_h I__5671 (
            .O(N__23920),
            .I(N__23779));
    LocalMux I__5670 (
            .O(N__23917),
            .I(N__23779));
    LocalMux I__5669 (
            .O(N__23914),
            .I(N__23779));
    LocalMux I__5668 (
            .O(N__23911),
            .I(N__23776));
    ClkMux I__5667 (
            .O(N__23910),
            .I(N__23773));
    ClkMux I__5666 (
            .O(N__23909),
            .I(N__23768));
    LocalMux I__5665 (
            .O(N__23906),
            .I(N__23765));
    Span4Mux_h I__5664 (
            .O(N__23899),
            .I(N__23759));
    Span4Mux_v I__5663 (
            .O(N__23892),
            .I(N__23759));
    Span4Mux_v I__5662 (
            .O(N__23883),
            .I(N__23756));
    Span4Mux_v I__5661 (
            .O(N__23876),
            .I(N__23749));
    Span4Mux_h I__5660 (
            .O(N__23873),
            .I(N__23749));
    LocalMux I__5659 (
            .O(N__23870),
            .I(N__23749));
    ClkMux I__5658 (
            .O(N__23869),
            .I(N__23746));
    Span4Mux_h I__5657 (
            .O(N__23862),
            .I(N__23742));
    Span4Mux_h I__5656 (
            .O(N__23859),
            .I(N__23739));
    LocalMux I__5655 (
            .O(N__23856),
            .I(N__23736));
    LocalMux I__5654 (
            .O(N__23853),
            .I(N__23732));
    ClkMux I__5653 (
            .O(N__23852),
            .I(N__23729));
    LocalMux I__5652 (
            .O(N__23849),
            .I(N__23726));
    LocalMux I__5651 (
            .O(N__23846),
            .I(N__23723));
    ClkMux I__5650 (
            .O(N__23845),
            .I(N__23720));
    Span4Mux_v I__5649 (
            .O(N__23842),
            .I(N__23713));
    LocalMux I__5648 (
            .O(N__23839),
            .I(N__23713));
    LocalMux I__5647 (
            .O(N__23836),
            .I(N__23713));
    ClkMux I__5646 (
            .O(N__23835),
            .I(N__23710));
    Span4Mux_h I__5645 (
            .O(N__23832),
            .I(N__23705));
    Span4Mux_v I__5644 (
            .O(N__23825),
            .I(N__23705));
    LocalMux I__5643 (
            .O(N__23822),
            .I(N__23702));
    Span4Mux_v I__5642 (
            .O(N__23819),
            .I(N__23697));
    LocalMux I__5641 (
            .O(N__23816),
            .I(N__23697));
    ClkMux I__5640 (
            .O(N__23815),
            .I(N__23694));
    LocalMux I__5639 (
            .O(N__23812),
            .I(N__23691));
    ClkMux I__5638 (
            .O(N__23811),
            .I(N__23688));
    LocalMux I__5637 (
            .O(N__23808),
            .I(N__23685));
    ClkMux I__5636 (
            .O(N__23807),
            .I(N__23682));
    LocalMux I__5635 (
            .O(N__23804),
            .I(N__23678));
    Span4Mux_v I__5634 (
            .O(N__23799),
            .I(N__23675));
    ClkMux I__5633 (
            .O(N__23798),
            .I(N__23672));
    Span4Mux_v I__5632 (
            .O(N__23795),
            .I(N__23665));
    Span4Mux_h I__5631 (
            .O(N__23786),
            .I(N__23665));
    Span4Mux_h I__5630 (
            .O(N__23779),
            .I(N__23665));
    Span4Mux_h I__5629 (
            .O(N__23776),
            .I(N__23660));
    LocalMux I__5628 (
            .O(N__23773),
            .I(N__23660));
    ClkMux I__5627 (
            .O(N__23772),
            .I(N__23657));
    ClkMux I__5626 (
            .O(N__23771),
            .I(N__23654));
    LocalMux I__5625 (
            .O(N__23768),
            .I(N__23650));
    IoSpan4Mux I__5624 (
            .O(N__23765),
            .I(N__23647));
    ClkMux I__5623 (
            .O(N__23764),
            .I(N__23644));
    Span4Mux_v I__5622 (
            .O(N__23759),
            .I(N__23640));
    Span4Mux_v I__5621 (
            .O(N__23756),
            .I(N__23637));
    Span4Mux_v I__5620 (
            .O(N__23749),
            .I(N__23634));
    LocalMux I__5619 (
            .O(N__23746),
            .I(N__23631));
    ClkMux I__5618 (
            .O(N__23745),
            .I(N__23628));
    Span4Mux_v I__5617 (
            .O(N__23742),
            .I(N__23625));
    Span4Mux_v I__5616 (
            .O(N__23739),
            .I(N__23620));
    Span4Mux_h I__5615 (
            .O(N__23736),
            .I(N__23620));
    ClkMux I__5614 (
            .O(N__23735),
            .I(N__23617));
    Span4Mux_h I__5613 (
            .O(N__23732),
            .I(N__23611));
    LocalMux I__5612 (
            .O(N__23729),
            .I(N__23611));
    Span4Mux_h I__5611 (
            .O(N__23726),
            .I(N__23604));
    Span4Mux_v I__5610 (
            .O(N__23723),
            .I(N__23604));
    LocalMux I__5609 (
            .O(N__23720),
            .I(N__23604));
    Span4Mux_v I__5608 (
            .O(N__23713),
            .I(N__23599));
    LocalMux I__5607 (
            .O(N__23710),
            .I(N__23599));
    Span4Mux_v I__5606 (
            .O(N__23705),
            .I(N__23590));
    Span4Mux_h I__5605 (
            .O(N__23702),
            .I(N__23590));
    Span4Mux_h I__5604 (
            .O(N__23697),
            .I(N__23590));
    LocalMux I__5603 (
            .O(N__23694),
            .I(N__23590));
    Span4Mux_h I__5602 (
            .O(N__23691),
            .I(N__23587));
    LocalMux I__5601 (
            .O(N__23688),
            .I(N__23584));
    Span4Mux_h I__5600 (
            .O(N__23685),
            .I(N__23579));
    LocalMux I__5599 (
            .O(N__23682),
            .I(N__23579));
    ClkMux I__5598 (
            .O(N__23681),
            .I(N__23576));
    Span4Mux_h I__5597 (
            .O(N__23678),
            .I(N__23573));
    Span4Mux_v I__5596 (
            .O(N__23675),
            .I(N__23568));
    LocalMux I__5595 (
            .O(N__23672),
            .I(N__23568));
    Span4Mux_v I__5594 (
            .O(N__23665),
            .I(N__23559));
    Span4Mux_h I__5593 (
            .O(N__23660),
            .I(N__23559));
    LocalMux I__5592 (
            .O(N__23657),
            .I(N__23559));
    LocalMux I__5591 (
            .O(N__23654),
            .I(N__23559));
    ClkMux I__5590 (
            .O(N__23653),
            .I(N__23556));
    Span4Mux_h I__5589 (
            .O(N__23650),
            .I(N__23553));
    Span4Mux_s1_v I__5588 (
            .O(N__23647),
            .I(N__23550));
    LocalMux I__5587 (
            .O(N__23644),
            .I(N__23547));
    ClkMux I__5586 (
            .O(N__23643),
            .I(N__23544));
    Span4Mux_v I__5585 (
            .O(N__23640),
            .I(N__23541));
    Span4Mux_v I__5584 (
            .O(N__23637),
            .I(N__23538));
    Sp12to4 I__5583 (
            .O(N__23634),
            .I(N__23533));
    Sp12to4 I__5582 (
            .O(N__23631),
            .I(N__23533));
    LocalMux I__5581 (
            .O(N__23628),
            .I(N__23530));
    Span4Mux_v I__5580 (
            .O(N__23625),
            .I(N__23527));
    Span4Mux_v I__5579 (
            .O(N__23620),
            .I(N__23522));
    LocalMux I__5578 (
            .O(N__23617),
            .I(N__23522));
    ClkMux I__5577 (
            .O(N__23616),
            .I(N__23519));
    Span4Mux_h I__5576 (
            .O(N__23611),
            .I(N__23516));
    Span4Mux_v I__5575 (
            .O(N__23604),
            .I(N__23509));
    Span4Mux_h I__5574 (
            .O(N__23599),
            .I(N__23509));
    Span4Mux_h I__5573 (
            .O(N__23590),
            .I(N__23509));
    Span4Mux_v I__5572 (
            .O(N__23587),
            .I(N__23504));
    Span4Mux_h I__5571 (
            .O(N__23584),
            .I(N__23504));
    Span4Mux_v I__5570 (
            .O(N__23579),
            .I(N__23499));
    LocalMux I__5569 (
            .O(N__23576),
            .I(N__23499));
    Span4Mux_h I__5568 (
            .O(N__23573),
            .I(N__23490));
    Span4Mux_h I__5567 (
            .O(N__23568),
            .I(N__23490));
    Span4Mux_h I__5566 (
            .O(N__23559),
            .I(N__23490));
    LocalMux I__5565 (
            .O(N__23556),
            .I(N__23490));
    Span4Mux_v I__5564 (
            .O(N__23553),
            .I(N__23483));
    Span4Mux_h I__5563 (
            .O(N__23550),
            .I(N__23483));
    Span4Mux_h I__5562 (
            .O(N__23547),
            .I(N__23483));
    LocalMux I__5561 (
            .O(N__23544),
            .I(N__23480));
    Span4Mux_v I__5560 (
            .O(N__23541),
            .I(N__23477));
    Span4Mux_v I__5559 (
            .O(N__23538),
            .I(N__23474));
    Span12Mux_h I__5558 (
            .O(N__23533),
            .I(N__23469));
    Span12Mux_h I__5557 (
            .O(N__23530),
            .I(N__23469));
    Sp12to4 I__5556 (
            .O(N__23527),
            .I(N__23464));
    Sp12to4 I__5555 (
            .O(N__23522),
            .I(N__23464));
    LocalMux I__5554 (
            .O(N__23519),
            .I(N__23461));
    Span4Mux_v I__5553 (
            .O(N__23516),
            .I(N__23458));
    Span4Mux_v I__5552 (
            .O(N__23509),
            .I(N__23455));
    Span4Mux_h I__5551 (
            .O(N__23504),
            .I(N__23452));
    Span4Mux_h I__5550 (
            .O(N__23499),
            .I(N__23449));
    Span4Mux_v I__5549 (
            .O(N__23490),
            .I(N__23446));
    Span4Mux_h I__5548 (
            .O(N__23483),
            .I(N__23443));
    Span4Mux_h I__5547 (
            .O(N__23480),
            .I(N__23440));
    IoSpan4Mux I__5546 (
            .O(N__23477),
            .I(N__23437));
    IoSpan4Mux I__5545 (
            .O(N__23474),
            .I(N__23434));
    Span12Mux_v I__5544 (
            .O(N__23469),
            .I(N__23425));
    Span12Mux_h I__5543 (
            .O(N__23464),
            .I(N__23425));
    Span12Mux_h I__5542 (
            .O(N__23461),
            .I(N__23425));
    Sp12to4 I__5541 (
            .O(N__23458),
            .I(N__23425));
    Span4Mux_v I__5540 (
            .O(N__23455),
            .I(N__23422));
    Span4Mux_h I__5539 (
            .O(N__23452),
            .I(N__23415));
    Span4Mux_h I__5538 (
            .O(N__23449),
            .I(N__23415));
    Span4Mux_v I__5537 (
            .O(N__23446),
            .I(N__23415));
    Span4Mux_h I__5536 (
            .O(N__23443),
            .I(N__23410));
    Span4Mux_h I__5535 (
            .O(N__23440),
            .I(N__23410));
    Odrv4 I__5534 (
            .O(N__23437),
            .I(ADV_CLK_c));
    Odrv4 I__5533 (
            .O(N__23434),
            .I(ADV_CLK_c));
    Odrv12 I__5532 (
            .O(N__23425),
            .I(ADV_CLK_c));
    Odrv4 I__5531 (
            .O(N__23422),
            .I(ADV_CLK_c));
    Odrv4 I__5530 (
            .O(N__23415),
            .I(ADV_CLK_c));
    Odrv4 I__5529 (
            .O(N__23410),
            .I(ADV_CLK_c));
    CEMux I__5528 (
            .O(N__23397),
            .I(N__23392));
    CEMux I__5527 (
            .O(N__23396),
            .I(N__23388));
    CEMux I__5526 (
            .O(N__23395),
            .I(N__23384));
    LocalMux I__5525 (
            .O(N__23392),
            .I(N__23381));
    CEMux I__5524 (
            .O(N__23391),
            .I(N__23378));
    LocalMux I__5523 (
            .O(N__23388),
            .I(N__23375));
    CEMux I__5522 (
            .O(N__23387),
            .I(N__23372));
    LocalMux I__5521 (
            .O(N__23384),
            .I(N__23369));
    Span4Mux_v I__5520 (
            .O(N__23381),
            .I(N__23364));
    LocalMux I__5519 (
            .O(N__23378),
            .I(N__23364));
    Span4Mux_h I__5518 (
            .O(N__23375),
            .I(N__23359));
    LocalMux I__5517 (
            .O(N__23372),
            .I(N__23359));
    Span4Mux_h I__5516 (
            .O(N__23369),
            .I(N__23356));
    Span4Mux_h I__5515 (
            .O(N__23364),
            .I(N__23351));
    Span4Mux_h I__5514 (
            .O(N__23359),
            .I(N__23351));
    Odrv4 I__5513 (
            .O(N__23356),
            .I(\transmit_module.n2206 ));
    Odrv4 I__5512 (
            .O(N__23351),
            .I(\transmit_module.n2206 ));
    IoInMux I__5511 (
            .O(N__23346),
            .I(N__23343));
    LocalMux I__5510 (
            .O(N__23343),
            .I(N__23340));
    IoSpan4Mux I__5509 (
            .O(N__23340),
            .I(N__23337));
    Span4Mux_s1_h I__5508 (
            .O(N__23337),
            .I(N__23328));
    SRMux I__5507 (
            .O(N__23336),
            .I(N__23320));
    SRMux I__5506 (
            .O(N__23335),
            .I(N__23317));
    SRMux I__5505 (
            .O(N__23334),
            .I(N__23314));
    SRMux I__5504 (
            .O(N__23333),
            .I(N__23311));
    SRMux I__5503 (
            .O(N__23332),
            .I(N__23307));
    SRMux I__5502 (
            .O(N__23331),
            .I(N__23304));
    Span4Mux_h I__5501 (
            .O(N__23328),
            .I(N__23293));
    SRMux I__5500 (
            .O(N__23327),
            .I(N__23290));
    SRMux I__5499 (
            .O(N__23326),
            .I(N__23287));
    SRMux I__5498 (
            .O(N__23325),
            .I(N__23277));
    SRMux I__5497 (
            .O(N__23324),
            .I(N__23271));
    SRMux I__5496 (
            .O(N__23323),
            .I(N__23268));
    LocalMux I__5495 (
            .O(N__23320),
            .I(N__23265));
    LocalMux I__5494 (
            .O(N__23317),
            .I(N__23262));
    LocalMux I__5493 (
            .O(N__23314),
            .I(N__23257));
    LocalMux I__5492 (
            .O(N__23311),
            .I(N__23257));
    SRMux I__5491 (
            .O(N__23310),
            .I(N__23254));
    LocalMux I__5490 (
            .O(N__23307),
            .I(N__23247));
    LocalMux I__5489 (
            .O(N__23304),
            .I(N__23247));
    SRMux I__5488 (
            .O(N__23303),
            .I(N__23244));
    CascadeMux I__5487 (
            .O(N__23302),
            .I(N__23235));
    CascadeMux I__5486 (
            .O(N__23301),
            .I(N__23230));
    SRMux I__5485 (
            .O(N__23300),
            .I(N__23225));
    CascadeMux I__5484 (
            .O(N__23299),
            .I(N__23220));
    CascadeMux I__5483 (
            .O(N__23298),
            .I(N__23217));
    CascadeMux I__5482 (
            .O(N__23297),
            .I(N__23214));
    SRMux I__5481 (
            .O(N__23296),
            .I(N__23209));
    Span4Mux_h I__5480 (
            .O(N__23293),
            .I(N__23202));
    LocalMux I__5479 (
            .O(N__23290),
            .I(N__23202));
    LocalMux I__5478 (
            .O(N__23287),
            .I(N__23202));
    InMux I__5477 (
            .O(N__23286),
            .I(N__23199));
    SRMux I__5476 (
            .O(N__23285),
            .I(N__23193));
    SRMux I__5475 (
            .O(N__23284),
            .I(N__23190));
    SRMux I__5474 (
            .O(N__23283),
            .I(N__23187));
    SRMux I__5473 (
            .O(N__23282),
            .I(N__23184));
    SRMux I__5472 (
            .O(N__23281),
            .I(N__23181));
    SRMux I__5471 (
            .O(N__23280),
            .I(N__23178));
    LocalMux I__5470 (
            .O(N__23277),
            .I(N__23175));
    SRMux I__5469 (
            .O(N__23276),
            .I(N__23171));
    SRMux I__5468 (
            .O(N__23275),
            .I(N__23168));
    SRMux I__5467 (
            .O(N__23274),
            .I(N__23165));
    LocalMux I__5466 (
            .O(N__23271),
            .I(N__23158));
    LocalMux I__5465 (
            .O(N__23268),
            .I(N__23158));
    Span4Mux_v I__5464 (
            .O(N__23265),
            .I(N__23158));
    Span4Mux_h I__5463 (
            .O(N__23262),
            .I(N__23151));
    Span4Mux_v I__5462 (
            .O(N__23257),
            .I(N__23151));
    LocalMux I__5461 (
            .O(N__23254),
            .I(N__23151));
    InMux I__5460 (
            .O(N__23253),
            .I(N__23148));
    SRMux I__5459 (
            .O(N__23252),
            .I(N__23145));
    Span4Mux_v I__5458 (
            .O(N__23247),
            .I(N__23135));
    LocalMux I__5457 (
            .O(N__23244),
            .I(N__23135));
    SRMux I__5456 (
            .O(N__23243),
            .I(N__23132));
    CascadeMux I__5455 (
            .O(N__23242),
            .I(N__23129));
    CascadeMux I__5454 (
            .O(N__23241),
            .I(N__23126));
    CascadeMux I__5453 (
            .O(N__23240),
            .I(N__23122));
    SRMux I__5452 (
            .O(N__23239),
            .I(N__23116));
    SRMux I__5451 (
            .O(N__23238),
            .I(N__23111));
    InMux I__5450 (
            .O(N__23235),
            .I(N__23111));
    InMux I__5449 (
            .O(N__23234),
            .I(N__23108));
    InMux I__5448 (
            .O(N__23233),
            .I(N__23101));
    InMux I__5447 (
            .O(N__23230),
            .I(N__23101));
    InMux I__5446 (
            .O(N__23229),
            .I(N__23101));
    SRMux I__5445 (
            .O(N__23228),
            .I(N__23098));
    LocalMux I__5444 (
            .O(N__23225),
            .I(N__23095));
    SRMux I__5443 (
            .O(N__23224),
            .I(N__23092));
    CascadeMux I__5442 (
            .O(N__23223),
            .I(N__23088));
    InMux I__5441 (
            .O(N__23220),
            .I(N__23083));
    InMux I__5440 (
            .O(N__23217),
            .I(N__23083));
    InMux I__5439 (
            .O(N__23214),
            .I(N__23080));
    InMux I__5438 (
            .O(N__23213),
            .I(N__23075));
    InMux I__5437 (
            .O(N__23212),
            .I(N__23075));
    LocalMux I__5436 (
            .O(N__23209),
            .I(N__23068));
    Span4Mux_v I__5435 (
            .O(N__23202),
            .I(N__23068));
    LocalMux I__5434 (
            .O(N__23199),
            .I(N__23068));
    SRMux I__5433 (
            .O(N__23198),
            .I(N__23065));
    SRMux I__5432 (
            .O(N__23197),
            .I(N__23062));
    SRMux I__5431 (
            .O(N__23196),
            .I(N__23059));
    LocalMux I__5430 (
            .O(N__23193),
            .I(N__23056));
    LocalMux I__5429 (
            .O(N__23190),
            .I(N__23053));
    LocalMux I__5428 (
            .O(N__23187),
            .I(N__23050));
    LocalMux I__5427 (
            .O(N__23184),
            .I(N__23047));
    LocalMux I__5426 (
            .O(N__23181),
            .I(N__23040));
    LocalMux I__5425 (
            .O(N__23178),
            .I(N__23040));
    Span4Mux_v I__5424 (
            .O(N__23175),
            .I(N__23040));
    CascadeMux I__5423 (
            .O(N__23174),
            .I(N__23037));
    LocalMux I__5422 (
            .O(N__23171),
            .I(N__23034));
    LocalMux I__5421 (
            .O(N__23168),
            .I(N__23031));
    LocalMux I__5420 (
            .O(N__23165),
            .I(N__23026));
    Span4Mux_v I__5419 (
            .O(N__23158),
            .I(N__23026));
    Span4Mux_v I__5418 (
            .O(N__23151),
            .I(N__23019));
    LocalMux I__5417 (
            .O(N__23148),
            .I(N__23019));
    LocalMux I__5416 (
            .O(N__23145),
            .I(N__23016));
    InMux I__5415 (
            .O(N__23144),
            .I(N__23007));
    InMux I__5414 (
            .O(N__23143),
            .I(N__23007));
    InMux I__5413 (
            .O(N__23142),
            .I(N__23007));
    InMux I__5412 (
            .O(N__23141),
            .I(N__23007));
    SRMux I__5411 (
            .O(N__23140),
            .I(N__23004));
    Span4Mux_v I__5410 (
            .O(N__23135),
            .I(N__23001));
    LocalMux I__5409 (
            .O(N__23132),
            .I(N__22998));
    InMux I__5408 (
            .O(N__23129),
            .I(N__22991));
    InMux I__5407 (
            .O(N__23126),
            .I(N__22991));
    InMux I__5406 (
            .O(N__23125),
            .I(N__22991));
    InMux I__5405 (
            .O(N__23122),
            .I(N__22982));
    InMux I__5404 (
            .O(N__23121),
            .I(N__22982));
    InMux I__5403 (
            .O(N__23120),
            .I(N__22982));
    InMux I__5402 (
            .O(N__23119),
            .I(N__22982));
    LocalMux I__5401 (
            .O(N__23116),
            .I(N__22973));
    LocalMux I__5400 (
            .O(N__23111),
            .I(N__22973));
    LocalMux I__5399 (
            .O(N__23108),
            .I(N__22973));
    LocalMux I__5398 (
            .O(N__23101),
            .I(N__22973));
    LocalMux I__5397 (
            .O(N__23098),
            .I(N__22970));
    Span4Mux_h I__5396 (
            .O(N__23095),
            .I(N__22965));
    LocalMux I__5395 (
            .O(N__23092),
            .I(N__22965));
    InMux I__5394 (
            .O(N__23091),
            .I(N__22960));
    InMux I__5393 (
            .O(N__23088),
            .I(N__22960));
    LocalMux I__5392 (
            .O(N__23083),
            .I(N__22951));
    LocalMux I__5391 (
            .O(N__23080),
            .I(N__22951));
    LocalMux I__5390 (
            .O(N__23075),
            .I(N__22951));
    Span4Mux_h I__5389 (
            .O(N__23068),
            .I(N__22951));
    LocalMux I__5388 (
            .O(N__23065),
            .I(N__22946));
    LocalMux I__5387 (
            .O(N__23062),
            .I(N__22946));
    LocalMux I__5386 (
            .O(N__23059),
            .I(N__22941));
    Span4Mux_h I__5385 (
            .O(N__23056),
            .I(N__22941));
    Span4Mux_h I__5384 (
            .O(N__23053),
            .I(N__22932));
    Span4Mux_v I__5383 (
            .O(N__23050),
            .I(N__22932));
    Span4Mux_v I__5382 (
            .O(N__23047),
            .I(N__22932));
    Span4Mux_h I__5381 (
            .O(N__23040),
            .I(N__22932));
    InMux I__5380 (
            .O(N__23037),
            .I(N__22929));
    Span4Mux_v I__5379 (
            .O(N__23034),
            .I(N__22922));
    Span4Mux_v I__5378 (
            .O(N__23031),
            .I(N__22922));
    Span4Mux_h I__5377 (
            .O(N__23026),
            .I(N__22922));
    InMux I__5376 (
            .O(N__23025),
            .I(N__22917));
    InMux I__5375 (
            .O(N__23024),
            .I(N__22917));
    Span4Mux_h I__5374 (
            .O(N__23019),
            .I(N__22910));
    Span4Mux_v I__5373 (
            .O(N__23016),
            .I(N__22910));
    LocalMux I__5372 (
            .O(N__23007),
            .I(N__22910));
    LocalMux I__5371 (
            .O(N__23004),
            .I(N__22897));
    Span4Mux_h I__5370 (
            .O(N__23001),
            .I(N__22897));
    Span4Mux_h I__5369 (
            .O(N__22998),
            .I(N__22897));
    LocalMux I__5368 (
            .O(N__22991),
            .I(N__22897));
    LocalMux I__5367 (
            .O(N__22982),
            .I(N__22897));
    Span4Mux_v I__5366 (
            .O(N__22973),
            .I(N__22897));
    Span4Mux_h I__5365 (
            .O(N__22970),
            .I(N__22888));
    Span4Mux_h I__5364 (
            .O(N__22965),
            .I(N__22888));
    LocalMux I__5363 (
            .O(N__22960),
            .I(N__22888));
    Span4Mux_v I__5362 (
            .O(N__22951),
            .I(N__22888));
    Odrv4 I__5361 (
            .O(N__22946),
            .I(ADV_VSYNC_c));
    Odrv4 I__5360 (
            .O(N__22941),
            .I(ADV_VSYNC_c));
    Odrv4 I__5359 (
            .O(N__22932),
            .I(ADV_VSYNC_c));
    LocalMux I__5358 (
            .O(N__22929),
            .I(ADV_VSYNC_c));
    Odrv4 I__5357 (
            .O(N__22922),
            .I(ADV_VSYNC_c));
    LocalMux I__5356 (
            .O(N__22917),
            .I(ADV_VSYNC_c));
    Odrv4 I__5355 (
            .O(N__22910),
            .I(ADV_VSYNC_c));
    Odrv4 I__5354 (
            .O(N__22897),
            .I(ADV_VSYNC_c));
    Odrv4 I__5353 (
            .O(N__22888),
            .I(ADV_VSYNC_c));
    InMux I__5352 (
            .O(N__22869),
            .I(N__22866));
    LocalMux I__5351 (
            .O(N__22866),
            .I(N__22863));
    Span12Mux_h I__5350 (
            .O(N__22863),
            .I(N__22860));
    Span12Mux_v I__5349 (
            .O(N__22860),
            .I(N__22857));
    Odrv12 I__5348 (
            .O(N__22857),
            .I(\line_buffer.n589 ));
    InMux I__5347 (
            .O(N__22854),
            .I(N__22851));
    LocalMux I__5346 (
            .O(N__22851),
            .I(N__22848));
    Span4Mux_v I__5345 (
            .O(N__22848),
            .I(N__22845));
    Sp12to4 I__5344 (
            .O(N__22845),
            .I(N__22842));
    Odrv12 I__5343 (
            .O(N__22842),
            .I(\line_buffer.n597 ));
    InMux I__5342 (
            .O(N__22839),
            .I(N__22836));
    LocalMux I__5341 (
            .O(N__22836),
            .I(\line_buffer.n3534 ));
    InMux I__5340 (
            .O(N__22833),
            .I(N__22822));
    InMux I__5339 (
            .O(N__22832),
            .I(N__22818));
    InMux I__5338 (
            .O(N__22831),
            .I(N__22815));
    InMux I__5337 (
            .O(N__22830),
            .I(N__22812));
    InMux I__5336 (
            .O(N__22829),
            .I(N__22809));
    InMux I__5335 (
            .O(N__22828),
            .I(N__22804));
    InMux I__5334 (
            .O(N__22827),
            .I(N__22799));
    InMux I__5333 (
            .O(N__22826),
            .I(N__22799));
    InMux I__5332 (
            .O(N__22825),
            .I(N__22795));
    LocalMux I__5331 (
            .O(N__22822),
            .I(N__22792));
    InMux I__5330 (
            .O(N__22821),
            .I(N__22789));
    LocalMux I__5329 (
            .O(N__22818),
            .I(N__22786));
    LocalMux I__5328 (
            .O(N__22815),
            .I(N__22783));
    LocalMux I__5327 (
            .O(N__22812),
            .I(N__22778));
    LocalMux I__5326 (
            .O(N__22809),
            .I(N__22778));
    InMux I__5325 (
            .O(N__22808),
            .I(N__22775));
    InMux I__5324 (
            .O(N__22807),
            .I(N__22772));
    LocalMux I__5323 (
            .O(N__22804),
            .I(N__22764));
    LocalMux I__5322 (
            .O(N__22799),
            .I(N__22760));
    InMux I__5321 (
            .O(N__22798),
            .I(N__22756));
    LocalMux I__5320 (
            .O(N__22795),
            .I(N__22748));
    Span4Mux_v I__5319 (
            .O(N__22792),
            .I(N__22748));
    LocalMux I__5318 (
            .O(N__22789),
            .I(N__22745));
    Span4Mux_h I__5317 (
            .O(N__22786),
            .I(N__22736));
    Span4Mux_h I__5316 (
            .O(N__22783),
            .I(N__22736));
    Span4Mux_v I__5315 (
            .O(N__22778),
            .I(N__22736));
    LocalMux I__5314 (
            .O(N__22775),
            .I(N__22736));
    LocalMux I__5313 (
            .O(N__22772),
            .I(N__22733));
    InMux I__5312 (
            .O(N__22771),
            .I(N__22730));
    InMux I__5311 (
            .O(N__22770),
            .I(N__22727));
    InMux I__5310 (
            .O(N__22769),
            .I(N__22724));
    InMux I__5309 (
            .O(N__22768),
            .I(N__22720));
    InMux I__5308 (
            .O(N__22767),
            .I(N__22717));
    Span4Mux_v I__5307 (
            .O(N__22764),
            .I(N__22714));
    InMux I__5306 (
            .O(N__22763),
            .I(N__22711));
    Span4Mux_h I__5305 (
            .O(N__22760),
            .I(N__22708));
    InMux I__5304 (
            .O(N__22759),
            .I(N__22704));
    LocalMux I__5303 (
            .O(N__22756),
            .I(N__22701));
    InMux I__5302 (
            .O(N__22755),
            .I(N__22698));
    InMux I__5301 (
            .O(N__22754),
            .I(N__22695));
    InMux I__5300 (
            .O(N__22753),
            .I(N__22692));
    Span4Mux_v I__5299 (
            .O(N__22748),
            .I(N__22689));
    Span4Mux_v I__5298 (
            .O(N__22745),
            .I(N__22684));
    Span4Mux_v I__5297 (
            .O(N__22736),
            .I(N__22684));
    Span4Mux_v I__5296 (
            .O(N__22733),
            .I(N__22675));
    LocalMux I__5295 (
            .O(N__22730),
            .I(N__22675));
    LocalMux I__5294 (
            .O(N__22727),
            .I(N__22675));
    LocalMux I__5293 (
            .O(N__22724),
            .I(N__22675));
    InMux I__5292 (
            .O(N__22723),
            .I(N__22672));
    LocalMux I__5291 (
            .O(N__22720),
            .I(N__22669));
    LocalMux I__5290 (
            .O(N__22717),
            .I(N__22662));
    Span4Mux_v I__5289 (
            .O(N__22714),
            .I(N__22662));
    LocalMux I__5288 (
            .O(N__22711),
            .I(N__22662));
    Span4Mux_h I__5287 (
            .O(N__22708),
            .I(N__22659));
    InMux I__5286 (
            .O(N__22707),
            .I(N__22656));
    LocalMux I__5285 (
            .O(N__22704),
            .I(N__22651));
    Span4Mux_h I__5284 (
            .O(N__22701),
            .I(N__22651));
    LocalMux I__5283 (
            .O(N__22698),
            .I(N__22648));
    LocalMux I__5282 (
            .O(N__22695),
            .I(N__22643));
    LocalMux I__5281 (
            .O(N__22692),
            .I(N__22643));
    Span4Mux_v I__5280 (
            .O(N__22689),
            .I(N__22634));
    Span4Mux_h I__5279 (
            .O(N__22684),
            .I(N__22634));
    Span4Mux_v I__5278 (
            .O(N__22675),
            .I(N__22634));
    LocalMux I__5277 (
            .O(N__22672),
            .I(N__22634));
    Span4Mux_h I__5276 (
            .O(N__22669),
            .I(N__22620));
    Span4Mux_h I__5275 (
            .O(N__22662),
            .I(N__22620));
    Span4Mux_v I__5274 (
            .O(N__22659),
            .I(N__22620));
    LocalMux I__5273 (
            .O(N__22656),
            .I(N__22620));
    Span4Mux_v I__5272 (
            .O(N__22651),
            .I(N__22620));
    Span4Mux_v I__5271 (
            .O(N__22648),
            .I(N__22620));
    Span4Mux_v I__5270 (
            .O(N__22643),
            .I(N__22617));
    Span4Mux_h I__5269 (
            .O(N__22634),
            .I(N__22614));
    InMux I__5268 (
            .O(N__22633),
            .I(N__22611));
    Odrv4 I__5267 (
            .O(N__22620),
            .I(TX_ADDR_11));
    Odrv4 I__5266 (
            .O(N__22617),
            .I(TX_ADDR_11));
    Odrv4 I__5265 (
            .O(N__22614),
            .I(TX_ADDR_11));
    LocalMux I__5264 (
            .O(N__22611),
            .I(TX_ADDR_11));
    InMux I__5263 (
            .O(N__22602),
            .I(N__22599));
    LocalMux I__5262 (
            .O(N__22599),
            .I(N__22596));
    Span4Mux_v I__5261 (
            .O(N__22596),
            .I(N__22593));
    Sp12to4 I__5260 (
            .O(N__22593),
            .I(N__22590));
    Odrv12 I__5259 (
            .O(N__22590),
            .I(\line_buffer.n535 ));
    InMux I__5258 (
            .O(N__22587),
            .I(N__22584));
    LocalMux I__5257 (
            .O(N__22584),
            .I(N__22581));
    Span4Mux_h I__5256 (
            .O(N__22581),
            .I(N__22578));
    Span4Mux_v I__5255 (
            .O(N__22578),
            .I(N__22575));
    Sp12to4 I__5254 (
            .O(N__22575),
            .I(N__22572));
    Span12Mux_v I__5253 (
            .O(N__22572),
            .I(N__22569));
    Odrv12 I__5252 (
            .O(N__22569),
            .I(\line_buffer.n527 ));
    InMux I__5251 (
            .O(N__22566),
            .I(N__22563));
    LocalMux I__5250 (
            .O(N__22563),
            .I(\line_buffer.n3539 ));
    InMux I__5249 (
            .O(N__22560),
            .I(N__22557));
    LocalMux I__5248 (
            .O(N__22557),
            .I(N__22554));
    Span4Mux_v I__5247 (
            .O(N__22554),
            .I(N__22551));
    Odrv4 I__5246 (
            .O(N__22551),
            .I(TX_DATA_4));
    IoInMux I__5245 (
            .O(N__22548),
            .I(N__22545));
    LocalMux I__5244 (
            .O(N__22545),
            .I(N__22542));
    IoSpan4Mux I__5243 (
            .O(N__22542),
            .I(N__22539));
    IoSpan4Mux I__5242 (
            .O(N__22539),
            .I(N__22535));
    IoInMux I__5241 (
            .O(N__22538),
            .I(N__22532));
    IoSpan4Mux I__5240 (
            .O(N__22535),
            .I(N__22526));
    LocalMux I__5239 (
            .O(N__22532),
            .I(N__22526));
    IoInMux I__5238 (
            .O(N__22531),
            .I(N__22523));
    IoSpan4Mux I__5237 (
            .O(N__22526),
            .I(N__22520));
    LocalMux I__5236 (
            .O(N__22523),
            .I(N__22517));
    Span4Mux_s2_h I__5235 (
            .O(N__22520),
            .I(N__22514));
    Span4Mux_s1_v I__5234 (
            .O(N__22517),
            .I(N__22511));
    Sp12to4 I__5233 (
            .O(N__22514),
            .I(N__22508));
    Sp12to4 I__5232 (
            .O(N__22511),
            .I(N__22505));
    Span12Mux_h I__5231 (
            .O(N__22508),
            .I(N__22502));
    Span12Mux_h I__5230 (
            .O(N__22505),
            .I(N__22499));
    Odrv12 I__5229 (
            .O(N__22502),
            .I(n1814));
    Odrv12 I__5228 (
            .O(N__22499),
            .I(n1814));
    InMux I__5227 (
            .O(N__22494),
            .I(N__22491));
    LocalMux I__5226 (
            .O(N__22491),
            .I(TX_DATA_6));
    IoInMux I__5225 (
            .O(N__22488),
            .I(N__22485));
    LocalMux I__5224 (
            .O(N__22485),
            .I(N__22482));
    IoSpan4Mux I__5223 (
            .O(N__22482),
            .I(N__22478));
    IoInMux I__5222 (
            .O(N__22481),
            .I(N__22474));
    Span4Mux_s1_h I__5221 (
            .O(N__22478),
            .I(N__22471));
    IoInMux I__5220 (
            .O(N__22477),
            .I(N__22468));
    LocalMux I__5219 (
            .O(N__22474),
            .I(N__22465));
    Span4Mux_h I__5218 (
            .O(N__22471),
            .I(N__22462));
    LocalMux I__5217 (
            .O(N__22468),
            .I(N__22459));
    Span4Mux_s3_v I__5216 (
            .O(N__22465),
            .I(N__22456));
    Span4Mux_h I__5215 (
            .O(N__22462),
            .I(N__22451));
    Span4Mux_s3_v I__5214 (
            .O(N__22459),
            .I(N__22451));
    Span4Mux_v I__5213 (
            .O(N__22456),
            .I(N__22448));
    Span4Mux_v I__5212 (
            .O(N__22451),
            .I(N__22445));
    Sp12to4 I__5211 (
            .O(N__22448),
            .I(N__22442));
    Sp12to4 I__5210 (
            .O(N__22445),
            .I(N__22439));
    Span12Mux_h I__5209 (
            .O(N__22442),
            .I(N__22434));
    Span12Mux_h I__5208 (
            .O(N__22439),
            .I(N__22434));
    Odrv12 I__5207 (
            .O(N__22434),
            .I(n1812));
    SRMux I__5206 (
            .O(N__22431),
            .I(N__22428));
    LocalMux I__5205 (
            .O(N__22428),
            .I(N__22421));
    SRMux I__5204 (
            .O(N__22427),
            .I(N__22418));
    SRMux I__5203 (
            .O(N__22426),
            .I(N__22415));
    SRMux I__5202 (
            .O(N__22425),
            .I(N__22411));
    SRMux I__5201 (
            .O(N__22424),
            .I(N__22408));
    Span4Mux_h I__5200 (
            .O(N__22421),
            .I(N__22401));
    LocalMux I__5199 (
            .O(N__22418),
            .I(N__22401));
    LocalMux I__5198 (
            .O(N__22415),
            .I(N__22401));
    SRMux I__5197 (
            .O(N__22414),
            .I(N__22398));
    LocalMux I__5196 (
            .O(N__22411),
            .I(N__22394));
    LocalMux I__5195 (
            .O(N__22408),
            .I(N__22391));
    Span4Mux_h I__5194 (
            .O(N__22401),
            .I(N__22386));
    LocalMux I__5193 (
            .O(N__22398),
            .I(N__22386));
    SRMux I__5192 (
            .O(N__22397),
            .I(N__22383));
    Span4Mux_h I__5191 (
            .O(N__22394),
            .I(N__22380));
    Span4Mux_v I__5190 (
            .O(N__22391),
            .I(N__22377));
    Span4Mux_h I__5189 (
            .O(N__22386),
            .I(N__22374));
    LocalMux I__5188 (
            .O(N__22383),
            .I(N__22371));
    Odrv4 I__5187 (
            .O(N__22380),
            .I(\transmit_module.n2385 ));
    Odrv4 I__5186 (
            .O(N__22377),
            .I(\transmit_module.n2385 ));
    Odrv4 I__5185 (
            .O(N__22374),
            .I(\transmit_module.n2385 ));
    Odrv12 I__5184 (
            .O(N__22371),
            .I(\transmit_module.n2385 ));
    InMux I__5183 (
            .O(N__22362),
            .I(N__22359));
    LocalMux I__5182 (
            .O(N__22359),
            .I(N__22356));
    Span4Mux_h I__5181 (
            .O(N__22356),
            .I(N__22353));
    Span4Mux_h I__5180 (
            .O(N__22353),
            .I(N__22350));
    Odrv4 I__5179 (
            .O(N__22350),
            .I(\line_buffer.n470 ));
    InMux I__5178 (
            .O(N__22347),
            .I(N__22344));
    LocalMux I__5177 (
            .O(N__22344),
            .I(N__22341));
    Span12Mux_v I__5176 (
            .O(N__22341),
            .I(N__22338));
    Odrv12 I__5175 (
            .O(N__22338),
            .I(\line_buffer.n462 ));
    InMux I__5174 (
            .O(N__22335),
            .I(N__22332));
    LocalMux I__5173 (
            .O(N__22332),
            .I(N__22329));
    Odrv4 I__5172 (
            .O(N__22329),
            .I(\line_buffer.n3572 ));
    SRMux I__5171 (
            .O(N__22326),
            .I(N__22323));
    LocalMux I__5170 (
            .O(N__22323),
            .I(N__22319));
    SRMux I__5169 (
            .O(N__22322),
            .I(N__22316));
    Span4Mux_h I__5168 (
            .O(N__22319),
            .I(N__22310));
    LocalMux I__5167 (
            .O(N__22316),
            .I(N__22310));
    SRMux I__5166 (
            .O(N__22315),
            .I(N__22307));
    Span4Mux_v I__5165 (
            .O(N__22310),
            .I(N__22301));
    LocalMux I__5164 (
            .O(N__22307),
            .I(N__22301));
    SRMux I__5163 (
            .O(N__22306),
            .I(N__22298));
    Span4Mux_h I__5162 (
            .O(N__22301),
            .I(N__22292));
    LocalMux I__5161 (
            .O(N__22298),
            .I(N__22292));
    SRMux I__5160 (
            .O(N__22297),
            .I(N__22289));
    Span4Mux_v I__5159 (
            .O(N__22292),
            .I(N__22283));
    LocalMux I__5158 (
            .O(N__22289),
            .I(N__22283));
    SRMux I__5157 (
            .O(N__22288),
            .I(N__22280));
    Span4Mux_h I__5156 (
            .O(N__22283),
            .I(N__22274));
    LocalMux I__5155 (
            .O(N__22280),
            .I(N__22274));
    SRMux I__5154 (
            .O(N__22279),
            .I(N__22271));
    Span4Mux_v I__5153 (
            .O(N__22274),
            .I(N__22264));
    LocalMux I__5152 (
            .O(N__22271),
            .I(N__22264));
    SRMux I__5151 (
            .O(N__22270),
            .I(N__22261));
    SRMux I__5150 (
            .O(N__22269),
            .I(N__22257));
    Span4Mux_h I__5149 (
            .O(N__22264),
            .I(N__22250));
    LocalMux I__5148 (
            .O(N__22261),
            .I(N__22250));
    SRMux I__5147 (
            .O(N__22260),
            .I(N__22247));
    LocalMux I__5146 (
            .O(N__22257),
            .I(N__22243));
    SRMux I__5145 (
            .O(N__22256),
            .I(N__22240));
    SRMux I__5144 (
            .O(N__22255),
            .I(N__22237));
    Span4Mux_v I__5143 (
            .O(N__22250),
            .I(N__22230));
    LocalMux I__5142 (
            .O(N__22247),
            .I(N__22230));
    SRMux I__5141 (
            .O(N__22246),
            .I(N__22227));
    Span4Mux_s1_v I__5140 (
            .O(N__22243),
            .I(N__22219));
    LocalMux I__5139 (
            .O(N__22240),
            .I(N__22219));
    LocalMux I__5138 (
            .O(N__22237),
            .I(N__22219));
    SRMux I__5137 (
            .O(N__22236),
            .I(N__22216));
    SRMux I__5136 (
            .O(N__22235),
            .I(N__22213));
    Span4Mux_h I__5135 (
            .O(N__22230),
            .I(N__22206));
    LocalMux I__5134 (
            .O(N__22227),
            .I(N__22206));
    SRMux I__5133 (
            .O(N__22226),
            .I(N__22203));
    Span4Mux_v I__5132 (
            .O(N__22219),
            .I(N__22195));
    LocalMux I__5131 (
            .O(N__22216),
            .I(N__22195));
    LocalMux I__5130 (
            .O(N__22213),
            .I(N__22195));
    SRMux I__5129 (
            .O(N__22212),
            .I(N__22192));
    SRMux I__5128 (
            .O(N__22211),
            .I(N__22189));
    Span4Mux_v I__5127 (
            .O(N__22206),
            .I(N__22182));
    LocalMux I__5126 (
            .O(N__22203),
            .I(N__22182));
    SRMux I__5125 (
            .O(N__22202),
            .I(N__22179));
    Span4Mux_v I__5124 (
            .O(N__22195),
            .I(N__22171));
    LocalMux I__5123 (
            .O(N__22192),
            .I(N__22171));
    LocalMux I__5122 (
            .O(N__22189),
            .I(N__22171));
    SRMux I__5121 (
            .O(N__22188),
            .I(N__22168));
    SRMux I__5120 (
            .O(N__22187),
            .I(N__22165));
    Span4Mux_h I__5119 (
            .O(N__22182),
            .I(N__22158));
    LocalMux I__5118 (
            .O(N__22179),
            .I(N__22158));
    SRMux I__5117 (
            .O(N__22178),
            .I(N__22155));
    Span4Mux_v I__5116 (
            .O(N__22171),
            .I(N__22146));
    LocalMux I__5115 (
            .O(N__22168),
            .I(N__22146));
    LocalMux I__5114 (
            .O(N__22165),
            .I(N__22146));
    SRMux I__5113 (
            .O(N__22164),
            .I(N__22143));
    SRMux I__5112 (
            .O(N__22163),
            .I(N__22140));
    Span4Mux_v I__5111 (
            .O(N__22158),
            .I(N__22133));
    LocalMux I__5110 (
            .O(N__22155),
            .I(N__22133));
    SRMux I__5109 (
            .O(N__22154),
            .I(N__22130));
    SRMux I__5108 (
            .O(N__22153),
            .I(N__22127));
    Span4Mux_v I__5107 (
            .O(N__22146),
            .I(N__22119));
    LocalMux I__5106 (
            .O(N__22143),
            .I(N__22119));
    LocalMux I__5105 (
            .O(N__22140),
            .I(N__22119));
    SRMux I__5104 (
            .O(N__22139),
            .I(N__22116));
    SRMux I__5103 (
            .O(N__22138),
            .I(N__22113));
    Span4Mux_h I__5102 (
            .O(N__22133),
            .I(N__22106));
    LocalMux I__5101 (
            .O(N__22130),
            .I(N__22106));
    LocalMux I__5100 (
            .O(N__22127),
            .I(N__22103));
    SRMux I__5099 (
            .O(N__22126),
            .I(N__22100));
    Span4Mux_v I__5098 (
            .O(N__22119),
            .I(N__22092));
    LocalMux I__5097 (
            .O(N__22116),
            .I(N__22092));
    LocalMux I__5096 (
            .O(N__22113),
            .I(N__22092));
    SRMux I__5095 (
            .O(N__22112),
            .I(N__22089));
    SRMux I__5094 (
            .O(N__22111),
            .I(N__22086));
    Span4Mux_v I__5093 (
            .O(N__22106),
            .I(N__22079));
    Span4Mux_s3_v I__5092 (
            .O(N__22103),
            .I(N__22079));
    LocalMux I__5091 (
            .O(N__22100),
            .I(N__22079));
    SRMux I__5090 (
            .O(N__22099),
            .I(N__22076));
    Span4Mux_v I__5089 (
            .O(N__22092),
            .I(N__22071));
    LocalMux I__5088 (
            .O(N__22089),
            .I(N__22071));
    LocalMux I__5087 (
            .O(N__22086),
            .I(N__22068));
    Span4Mux_h I__5086 (
            .O(N__22079),
            .I(N__22065));
    LocalMux I__5085 (
            .O(N__22076),
            .I(N__22061));
    Span4Mux_v I__5084 (
            .O(N__22071),
            .I(N__22055));
    Span4Mux_s2_v I__5083 (
            .O(N__22068),
            .I(N__22055));
    Span4Mux_h I__5082 (
            .O(N__22065),
            .I(N__22052));
    IoInMux I__5081 (
            .O(N__22064),
            .I(N__22049));
    Span4Mux_h I__5080 (
            .O(N__22061),
            .I(N__22046));
    IoInMux I__5079 (
            .O(N__22060),
            .I(N__22043));
    Span4Mux_h I__5078 (
            .O(N__22055),
            .I(N__22040));
    Span4Mux_h I__5077 (
            .O(N__22052),
            .I(N__22031));
    LocalMux I__5076 (
            .O(N__22049),
            .I(N__22031));
    Span4Mux_h I__5075 (
            .O(N__22046),
            .I(N__22031));
    LocalMux I__5074 (
            .O(N__22043),
            .I(N__22031));
    Odrv4 I__5073 (
            .O(N__22040),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__5072 (
            .O(N__22031),
            .I(CONSTANT_ONE_NET));
    InMux I__5071 (
            .O(N__22026),
            .I(N__22023));
    LocalMux I__5070 (
            .O(N__22023),
            .I(N__22020));
    Span4Mux_h I__5069 (
            .O(N__22020),
            .I(N__22017));
    Span4Mux_v I__5068 (
            .O(N__22017),
            .I(N__22014));
    Odrv4 I__5067 (
            .O(N__22014),
            .I(TVP_VIDEO_c_9));
    InMux I__5066 (
            .O(N__22011),
            .I(N__22008));
    LocalMux I__5065 (
            .O(N__22008),
            .I(\tvp_video_buffer.BUFFER_0_9 ));
    InMux I__5064 (
            .O(N__22005),
            .I(N__22002));
    LocalMux I__5063 (
            .O(N__22002),
            .I(\tvp_video_buffer.BUFFER_1_9 ));
    InMux I__5062 (
            .O(N__21999),
            .I(N__21996));
    LocalMux I__5061 (
            .O(N__21996),
            .I(N__21978));
    ClkMux I__5060 (
            .O(N__21995),
            .I(N__21789));
    ClkMux I__5059 (
            .O(N__21994),
            .I(N__21789));
    ClkMux I__5058 (
            .O(N__21993),
            .I(N__21789));
    ClkMux I__5057 (
            .O(N__21992),
            .I(N__21789));
    ClkMux I__5056 (
            .O(N__21991),
            .I(N__21789));
    ClkMux I__5055 (
            .O(N__21990),
            .I(N__21789));
    ClkMux I__5054 (
            .O(N__21989),
            .I(N__21789));
    ClkMux I__5053 (
            .O(N__21988),
            .I(N__21789));
    ClkMux I__5052 (
            .O(N__21987),
            .I(N__21789));
    ClkMux I__5051 (
            .O(N__21986),
            .I(N__21789));
    ClkMux I__5050 (
            .O(N__21985),
            .I(N__21789));
    ClkMux I__5049 (
            .O(N__21984),
            .I(N__21789));
    ClkMux I__5048 (
            .O(N__21983),
            .I(N__21789));
    ClkMux I__5047 (
            .O(N__21982),
            .I(N__21789));
    ClkMux I__5046 (
            .O(N__21981),
            .I(N__21789));
    Glb2LocalMux I__5045 (
            .O(N__21978),
            .I(N__21789));
    ClkMux I__5044 (
            .O(N__21977),
            .I(N__21789));
    ClkMux I__5043 (
            .O(N__21976),
            .I(N__21789));
    ClkMux I__5042 (
            .O(N__21975),
            .I(N__21789));
    ClkMux I__5041 (
            .O(N__21974),
            .I(N__21789));
    ClkMux I__5040 (
            .O(N__21973),
            .I(N__21789));
    ClkMux I__5039 (
            .O(N__21972),
            .I(N__21789));
    ClkMux I__5038 (
            .O(N__21971),
            .I(N__21789));
    ClkMux I__5037 (
            .O(N__21970),
            .I(N__21789));
    ClkMux I__5036 (
            .O(N__21969),
            .I(N__21789));
    ClkMux I__5035 (
            .O(N__21968),
            .I(N__21789));
    ClkMux I__5034 (
            .O(N__21967),
            .I(N__21789));
    ClkMux I__5033 (
            .O(N__21966),
            .I(N__21789));
    ClkMux I__5032 (
            .O(N__21965),
            .I(N__21789));
    ClkMux I__5031 (
            .O(N__21964),
            .I(N__21789));
    ClkMux I__5030 (
            .O(N__21963),
            .I(N__21789));
    ClkMux I__5029 (
            .O(N__21962),
            .I(N__21789));
    ClkMux I__5028 (
            .O(N__21961),
            .I(N__21789));
    ClkMux I__5027 (
            .O(N__21960),
            .I(N__21789));
    ClkMux I__5026 (
            .O(N__21959),
            .I(N__21789));
    ClkMux I__5025 (
            .O(N__21958),
            .I(N__21789));
    ClkMux I__5024 (
            .O(N__21957),
            .I(N__21789));
    ClkMux I__5023 (
            .O(N__21956),
            .I(N__21789));
    ClkMux I__5022 (
            .O(N__21955),
            .I(N__21789));
    ClkMux I__5021 (
            .O(N__21954),
            .I(N__21789));
    ClkMux I__5020 (
            .O(N__21953),
            .I(N__21789));
    ClkMux I__5019 (
            .O(N__21952),
            .I(N__21789));
    ClkMux I__5018 (
            .O(N__21951),
            .I(N__21789));
    ClkMux I__5017 (
            .O(N__21950),
            .I(N__21789));
    ClkMux I__5016 (
            .O(N__21949),
            .I(N__21789));
    ClkMux I__5015 (
            .O(N__21948),
            .I(N__21789));
    ClkMux I__5014 (
            .O(N__21947),
            .I(N__21789));
    ClkMux I__5013 (
            .O(N__21946),
            .I(N__21789));
    ClkMux I__5012 (
            .O(N__21945),
            .I(N__21789));
    ClkMux I__5011 (
            .O(N__21944),
            .I(N__21789));
    ClkMux I__5010 (
            .O(N__21943),
            .I(N__21789));
    ClkMux I__5009 (
            .O(N__21942),
            .I(N__21789));
    ClkMux I__5008 (
            .O(N__21941),
            .I(N__21789));
    ClkMux I__5007 (
            .O(N__21940),
            .I(N__21789));
    ClkMux I__5006 (
            .O(N__21939),
            .I(N__21789));
    ClkMux I__5005 (
            .O(N__21938),
            .I(N__21789));
    ClkMux I__5004 (
            .O(N__21937),
            .I(N__21789));
    ClkMux I__5003 (
            .O(N__21936),
            .I(N__21789));
    ClkMux I__5002 (
            .O(N__21935),
            .I(N__21789));
    ClkMux I__5001 (
            .O(N__21934),
            .I(N__21789));
    ClkMux I__5000 (
            .O(N__21933),
            .I(N__21789));
    ClkMux I__4999 (
            .O(N__21932),
            .I(N__21789));
    ClkMux I__4998 (
            .O(N__21931),
            .I(N__21789));
    ClkMux I__4997 (
            .O(N__21930),
            .I(N__21789));
    ClkMux I__4996 (
            .O(N__21929),
            .I(N__21789));
    ClkMux I__4995 (
            .O(N__21928),
            .I(N__21789));
    ClkMux I__4994 (
            .O(N__21927),
            .I(N__21789));
    ClkMux I__4993 (
            .O(N__21926),
            .I(N__21789));
    GlobalMux I__4992 (
            .O(N__21789),
            .I(N__21786));
    gio2CtrlBuf I__4991 (
            .O(N__21786),
            .I(DEBUG_c_3_c));
    InMux I__4990 (
            .O(N__21783),
            .I(N__21780));
    LocalMux I__4989 (
            .O(N__21780),
            .I(N__21777));
    Odrv4 I__4988 (
            .O(N__21777),
            .I(\transmit_module.Y_DELTA_PATTERN_88 ));
    InMux I__4987 (
            .O(N__21774),
            .I(N__21771));
    LocalMux I__4986 (
            .O(N__21771),
            .I(N__21768));
    Span4Mux_v I__4985 (
            .O(N__21768),
            .I(N__21765));
    Odrv4 I__4984 (
            .O(N__21765),
            .I(\transmit_module.Y_DELTA_PATTERN_84 ));
    InMux I__4983 (
            .O(N__21762),
            .I(N__21759));
    LocalMux I__4982 (
            .O(N__21759),
            .I(N__21756));
    Sp12to4 I__4981 (
            .O(N__21756),
            .I(N__21753));
    Odrv12 I__4980 (
            .O(N__21753),
            .I(\line_buffer.n3533 ));
    InMux I__4979 (
            .O(N__21750),
            .I(N__21747));
    LocalMux I__4978 (
            .O(N__21747),
            .I(N__21744));
    Odrv4 I__4977 (
            .O(N__21744),
            .I(\line_buffer.n3549 ));
    CascadeMux I__4976 (
            .O(N__21741),
            .I(\line_buffer.n3611_cascade_ ));
    InMux I__4975 (
            .O(N__21738),
            .I(N__21734));
    InMux I__4974 (
            .O(N__21737),
            .I(N__21731));
    LocalMux I__4973 (
            .O(N__21734),
            .I(N__21728));
    LocalMux I__4972 (
            .O(N__21731),
            .I(N__21721));
    Span4Mux_v I__4971 (
            .O(N__21728),
            .I(N__21718));
    InMux I__4970 (
            .O(N__21727),
            .I(N__21715));
    InMux I__4969 (
            .O(N__21726),
            .I(N__21711));
    InMux I__4968 (
            .O(N__21725),
            .I(N__21708));
    InMux I__4967 (
            .O(N__21724),
            .I(N__21705));
    Span4Mux_v I__4966 (
            .O(N__21721),
            .I(N__21701));
    Span4Mux_v I__4965 (
            .O(N__21718),
            .I(N__21696));
    LocalMux I__4964 (
            .O(N__21715),
            .I(N__21696));
    InMux I__4963 (
            .O(N__21714),
            .I(N__21693));
    LocalMux I__4962 (
            .O(N__21711),
            .I(N__21689));
    LocalMux I__4961 (
            .O(N__21708),
            .I(N__21686));
    LocalMux I__4960 (
            .O(N__21705),
            .I(N__21683));
    InMux I__4959 (
            .O(N__21704),
            .I(N__21680));
    Span4Mux_v I__4958 (
            .O(N__21701),
            .I(N__21673));
    Span4Mux_v I__4957 (
            .O(N__21696),
            .I(N__21673));
    LocalMux I__4956 (
            .O(N__21693),
            .I(N__21673));
    InMux I__4955 (
            .O(N__21692),
            .I(N__21670));
    Span12Mux_s5_v I__4954 (
            .O(N__21689),
            .I(N__21667));
    Span12Mux_s6_v I__4953 (
            .O(N__21686),
            .I(N__21664));
    Span12Mux_v I__4952 (
            .O(N__21683),
            .I(N__21659));
    LocalMux I__4951 (
            .O(N__21680),
            .I(N__21659));
    Span4Mux_v I__4950 (
            .O(N__21673),
            .I(N__21656));
    LocalMux I__4949 (
            .O(N__21670),
            .I(N__21653));
    Span12Mux_h I__4948 (
            .O(N__21667),
            .I(N__21650));
    Span12Mux_h I__4947 (
            .O(N__21664),
            .I(N__21645));
    Span12Mux_h I__4946 (
            .O(N__21659),
            .I(N__21645));
    Sp12to4 I__4945 (
            .O(N__21656),
            .I(N__21640));
    Span12Mux_v I__4944 (
            .O(N__21653),
            .I(N__21640));
    Odrv12 I__4943 (
            .O(N__21650),
            .I(RX_DATA_4));
    Odrv12 I__4942 (
            .O(N__21645),
            .I(RX_DATA_4));
    Odrv12 I__4941 (
            .O(N__21640),
            .I(RX_DATA_4));
    InMux I__4940 (
            .O(N__21633),
            .I(N__21630));
    LocalMux I__4939 (
            .O(N__21630),
            .I(\tvp_video_buffer.BUFFER_1_6 ));
    IoInMux I__4938 (
            .O(N__21627),
            .I(N__21624));
    LocalMux I__4937 (
            .O(N__21624),
            .I(N__21620));
    InMux I__4936 (
            .O(N__21623),
            .I(N__21617));
    IoSpan4Mux I__4935 (
            .O(N__21620),
            .I(N__21614));
    LocalMux I__4934 (
            .O(N__21617),
            .I(N__21611));
    Span4Mux_s0_h I__4933 (
            .O(N__21614),
            .I(N__21608));
    Span4Mux_h I__4932 (
            .O(N__21611),
            .I(N__21605));
    Sp12to4 I__4931 (
            .O(N__21608),
            .I(N__21602));
    Sp12to4 I__4930 (
            .O(N__21605),
            .I(N__21599));
    Span12Mux_s11_h I__4929 (
            .O(N__21602),
            .I(N__21596));
    Span12Mux_v I__4928 (
            .O(N__21599),
            .I(N__21593));
    Span12Mux_v I__4927 (
            .O(N__21596),
            .I(N__21588));
    Span12Mux_h I__4926 (
            .O(N__21593),
            .I(N__21588));
    Odrv12 I__4925 (
            .O(N__21588),
            .I(DEBUG_c_5_c));
    InMux I__4924 (
            .O(N__21585),
            .I(N__21582));
    LocalMux I__4923 (
            .O(N__21582),
            .I(\tvp_video_buffer.BUFFER_0_6 ));
    InMux I__4922 (
            .O(N__21579),
            .I(N__21576));
    LocalMux I__4921 (
            .O(N__21576),
            .I(N__21573));
    Span4Mux_h I__4920 (
            .O(N__21573),
            .I(N__21570));
    Span4Mux_h I__4919 (
            .O(N__21570),
            .I(N__21567));
    Odrv4 I__4918 (
            .O(N__21567),
            .I(\line_buffer.n468 ));
    InMux I__4917 (
            .O(N__21564),
            .I(N__21561));
    LocalMux I__4916 (
            .O(N__21561),
            .I(N__21558));
    Span12Mux_h I__4915 (
            .O(N__21558),
            .I(N__21555));
    Span12Mux_v I__4914 (
            .O(N__21555),
            .I(N__21552));
    Odrv12 I__4913 (
            .O(N__21552),
            .I(\line_buffer.n460 ));
    InMux I__4912 (
            .O(N__21549),
            .I(N__21546));
    LocalMux I__4911 (
            .O(N__21546),
            .I(N__21543));
    Odrv4 I__4910 (
            .O(N__21543),
            .I(\line_buffer.n3548 ));
    InMux I__4909 (
            .O(N__21540),
            .I(N__21537));
    LocalMux I__4908 (
            .O(N__21537),
            .I(N__21534));
    Span12Mux_v I__4907 (
            .O(N__21534),
            .I(N__21531));
    Odrv12 I__4906 (
            .O(N__21531),
            .I(\line_buffer.n567 ));
    InMux I__4905 (
            .O(N__21528),
            .I(N__21525));
    LocalMux I__4904 (
            .O(N__21525),
            .I(N__21522));
    Span4Mux_h I__4903 (
            .O(N__21522),
            .I(N__21519));
    Sp12to4 I__4902 (
            .O(N__21519),
            .I(N__21516));
    Span12Mux_s7_h I__4901 (
            .O(N__21516),
            .I(N__21513));
    Span12Mux_v I__4900 (
            .O(N__21513),
            .I(N__21510));
    Odrv12 I__4899 (
            .O(N__21510),
            .I(\line_buffer.n559 ));
    InMux I__4898 (
            .O(N__21507),
            .I(N__21494));
    InMux I__4897 (
            .O(N__21506),
            .I(N__21491));
    CascadeMux I__4896 (
            .O(N__21505),
            .I(N__21488));
    CascadeMux I__4895 (
            .O(N__21504),
            .I(N__21485));
    CascadeMux I__4894 (
            .O(N__21503),
            .I(N__21480));
    CascadeMux I__4893 (
            .O(N__21502),
            .I(N__21475));
    CascadeMux I__4892 (
            .O(N__21501),
            .I(N__21471));
    InMux I__4891 (
            .O(N__21500),
            .I(N__21468));
    CascadeMux I__4890 (
            .O(N__21499),
            .I(N__21465));
    InMux I__4889 (
            .O(N__21498),
            .I(N__21460));
    CascadeMux I__4888 (
            .O(N__21497),
            .I(N__21455));
    LocalMux I__4887 (
            .O(N__21494),
            .I(N__21452));
    LocalMux I__4886 (
            .O(N__21491),
            .I(N__21449));
    InMux I__4885 (
            .O(N__21488),
            .I(N__21446));
    InMux I__4884 (
            .O(N__21485),
            .I(N__21443));
    InMux I__4883 (
            .O(N__21484),
            .I(N__21440));
    InMux I__4882 (
            .O(N__21483),
            .I(N__21436));
    InMux I__4881 (
            .O(N__21480),
            .I(N__21433));
    InMux I__4880 (
            .O(N__21479),
            .I(N__21426));
    InMux I__4879 (
            .O(N__21478),
            .I(N__21426));
    InMux I__4878 (
            .O(N__21475),
            .I(N__21426));
    InMux I__4877 (
            .O(N__21474),
            .I(N__21421));
    InMux I__4876 (
            .O(N__21471),
            .I(N__21421));
    LocalMux I__4875 (
            .O(N__21468),
            .I(N__21418));
    InMux I__4874 (
            .O(N__21465),
            .I(N__21415));
    CascadeMux I__4873 (
            .O(N__21464),
            .I(N__21411));
    CascadeMux I__4872 (
            .O(N__21463),
            .I(N__21408));
    LocalMux I__4871 (
            .O(N__21460),
            .I(N__21405));
    InMux I__4870 (
            .O(N__21459),
            .I(N__21402));
    InMux I__4869 (
            .O(N__21458),
            .I(N__21397));
    InMux I__4868 (
            .O(N__21455),
            .I(N__21397));
    Span4Mux_v I__4867 (
            .O(N__21452),
            .I(N__21394));
    Span4Mux_h I__4866 (
            .O(N__21449),
            .I(N__21389));
    LocalMux I__4865 (
            .O(N__21446),
            .I(N__21389));
    LocalMux I__4864 (
            .O(N__21443),
            .I(N__21386));
    LocalMux I__4863 (
            .O(N__21440),
            .I(N__21383));
    InMux I__4862 (
            .O(N__21439),
            .I(N__21380));
    LocalMux I__4861 (
            .O(N__21436),
            .I(N__21367));
    LocalMux I__4860 (
            .O(N__21433),
            .I(N__21367));
    LocalMux I__4859 (
            .O(N__21426),
            .I(N__21367));
    LocalMux I__4858 (
            .O(N__21421),
            .I(N__21367));
    Span4Mux_h I__4857 (
            .O(N__21418),
            .I(N__21367));
    LocalMux I__4856 (
            .O(N__21415),
            .I(N__21367));
    InMux I__4855 (
            .O(N__21414),
            .I(N__21362));
    InMux I__4854 (
            .O(N__21411),
            .I(N__21362));
    InMux I__4853 (
            .O(N__21408),
            .I(N__21359));
    Span4Mux_v I__4852 (
            .O(N__21405),
            .I(N__21356));
    LocalMux I__4851 (
            .O(N__21402),
            .I(N__21351));
    LocalMux I__4850 (
            .O(N__21397),
            .I(N__21351));
    Span4Mux_h I__4849 (
            .O(N__21394),
            .I(N__21344));
    Span4Mux_h I__4848 (
            .O(N__21389),
            .I(N__21344));
    Span4Mux_h I__4847 (
            .O(N__21386),
            .I(N__21344));
    Span4Mux_v I__4846 (
            .O(N__21383),
            .I(N__21337));
    LocalMux I__4845 (
            .O(N__21380),
            .I(N__21337));
    Span4Mux_v I__4844 (
            .O(N__21367),
            .I(N__21337));
    LocalMux I__4843 (
            .O(N__21362),
            .I(TX_ADDR_12));
    LocalMux I__4842 (
            .O(N__21359),
            .I(TX_ADDR_12));
    Odrv4 I__4841 (
            .O(N__21356),
            .I(TX_ADDR_12));
    Odrv12 I__4840 (
            .O(N__21351),
            .I(TX_ADDR_12));
    Odrv4 I__4839 (
            .O(N__21344),
            .I(TX_ADDR_12));
    Odrv4 I__4838 (
            .O(N__21337),
            .I(TX_ADDR_12));
    InMux I__4837 (
            .O(N__21324),
            .I(N__21321));
    LocalMux I__4836 (
            .O(N__21321),
            .I(N__21318));
    Span12Mux_h I__4835 (
            .O(N__21318),
            .I(N__21315));
    Odrv12 I__4834 (
            .O(N__21315),
            .I(\line_buffer.n3540 ));
    InMux I__4833 (
            .O(N__21312),
            .I(N__21309));
    LocalMux I__4832 (
            .O(N__21309),
            .I(\line_buffer.n3573 ));
    CascadeMux I__4831 (
            .O(N__21306),
            .I(N__21301));
    CascadeMux I__4830 (
            .O(N__21305),
            .I(N__21296));
    InMux I__4829 (
            .O(N__21304),
            .I(N__21290));
    InMux I__4828 (
            .O(N__21301),
            .I(N__21287));
    CascadeMux I__4827 (
            .O(N__21300),
            .I(N__21284));
    CascadeMux I__4826 (
            .O(N__21299),
            .I(N__21280));
    InMux I__4825 (
            .O(N__21296),
            .I(N__21277));
    CascadeMux I__4824 (
            .O(N__21295),
            .I(N__21274));
    InMux I__4823 (
            .O(N__21294),
            .I(N__21271));
    InMux I__4822 (
            .O(N__21293),
            .I(N__21264));
    LocalMux I__4821 (
            .O(N__21290),
            .I(N__21261));
    LocalMux I__4820 (
            .O(N__21287),
            .I(N__21258));
    InMux I__4819 (
            .O(N__21284),
            .I(N__21255));
    InMux I__4818 (
            .O(N__21283),
            .I(N__21252));
    InMux I__4817 (
            .O(N__21280),
            .I(N__21249));
    LocalMux I__4816 (
            .O(N__21277),
            .I(N__21246));
    InMux I__4815 (
            .O(N__21274),
            .I(N__21243));
    LocalMux I__4814 (
            .O(N__21271),
            .I(N__21240));
    InMux I__4813 (
            .O(N__21270),
            .I(N__21237));
    InMux I__4812 (
            .O(N__21269),
            .I(N__21232));
    InMux I__4811 (
            .O(N__21268),
            .I(N__21232));
    InMux I__4810 (
            .O(N__21267),
            .I(N__21229));
    LocalMux I__4809 (
            .O(N__21264),
            .I(N__21225));
    Span4Mux_v I__4808 (
            .O(N__21261),
            .I(N__21220));
    Span4Mux_v I__4807 (
            .O(N__21258),
            .I(N__21220));
    LocalMux I__4806 (
            .O(N__21255),
            .I(N__21217));
    LocalMux I__4805 (
            .O(N__21252),
            .I(N__21212));
    LocalMux I__4804 (
            .O(N__21249),
            .I(N__21212));
    Span4Mux_v I__4803 (
            .O(N__21246),
            .I(N__21207));
    LocalMux I__4802 (
            .O(N__21243),
            .I(N__21207));
    Span4Mux_v I__4801 (
            .O(N__21240),
            .I(N__21202));
    LocalMux I__4800 (
            .O(N__21237),
            .I(N__21202));
    LocalMux I__4799 (
            .O(N__21232),
            .I(N__21197));
    LocalMux I__4798 (
            .O(N__21229),
            .I(N__21197));
    InMux I__4797 (
            .O(N__21228),
            .I(N__21194));
    Span4Mux_v I__4796 (
            .O(N__21225),
            .I(N__21189));
    Span4Mux_h I__4795 (
            .O(N__21220),
            .I(N__21189));
    Span4Mux_v I__4794 (
            .O(N__21217),
            .I(N__21186));
    Span4Mux_v I__4793 (
            .O(N__21212),
            .I(N__21181));
    Span4Mux_v I__4792 (
            .O(N__21207),
            .I(N__21181));
    Span4Mux_v I__4791 (
            .O(N__21202),
            .I(N__21174));
    Span4Mux_v I__4790 (
            .O(N__21197),
            .I(N__21174));
    LocalMux I__4789 (
            .O(N__21194),
            .I(N__21174));
    Odrv4 I__4788 (
            .O(N__21189),
            .I(TX_ADDR_13));
    Odrv4 I__4787 (
            .O(N__21186),
            .I(TX_ADDR_13));
    Odrv4 I__4786 (
            .O(N__21181),
            .I(TX_ADDR_13));
    Odrv4 I__4785 (
            .O(N__21174),
            .I(TX_ADDR_13));
    InMux I__4784 (
            .O(N__21165),
            .I(N__21162));
    LocalMux I__4783 (
            .O(N__21162),
            .I(\line_buffer.n3605 ));
    InMux I__4782 (
            .O(N__21159),
            .I(N__21156));
    LocalMux I__4781 (
            .O(N__21156),
            .I(\transmit_module.Y_DELTA_PATTERN_96 ));
    InMux I__4780 (
            .O(N__21153),
            .I(N__21150));
    LocalMux I__4779 (
            .O(N__21150),
            .I(\transmit_module.Y_DELTA_PATTERN_95 ));
    InMux I__4778 (
            .O(N__21147),
            .I(N__21144));
    LocalMux I__4777 (
            .O(N__21144),
            .I(\transmit_module.Y_DELTA_PATTERN_94 ));
    InMux I__4776 (
            .O(N__21141),
            .I(N__21138));
    LocalMux I__4775 (
            .O(N__21138),
            .I(\transmit_module.Y_DELTA_PATTERN_93 ));
    InMux I__4774 (
            .O(N__21135),
            .I(N__21132));
    LocalMux I__4773 (
            .O(N__21132),
            .I(N__21129));
    Odrv12 I__4772 (
            .O(N__21129),
            .I(\transmit_module.Y_DELTA_PATTERN_83 ));
    InMux I__4771 (
            .O(N__21126),
            .I(N__21123));
    LocalMux I__4770 (
            .O(N__21123),
            .I(N__21120));
    Span4Mux_v I__4769 (
            .O(N__21120),
            .I(N__21117));
    Sp12to4 I__4768 (
            .O(N__21117),
            .I(N__21114));
    Odrv12 I__4767 (
            .O(N__21114),
            .I(\line_buffer.n593 ));
    InMux I__4766 (
            .O(N__21111),
            .I(N__21108));
    LocalMux I__4765 (
            .O(N__21108),
            .I(N__21105));
    Span4Mux_v I__4764 (
            .O(N__21105),
            .I(N__21102));
    Sp12to4 I__4763 (
            .O(N__21102),
            .I(N__21099));
    Span12Mux_h I__4762 (
            .O(N__21099),
            .I(N__21096));
    Span12Mux_v I__4761 (
            .O(N__21096),
            .I(N__21093));
    Odrv12 I__4760 (
            .O(N__21093),
            .I(\line_buffer.n585 ));
    InMux I__4759 (
            .O(N__21090),
            .I(N__21087));
    LocalMux I__4758 (
            .O(N__21087),
            .I(\line_buffer.n3641 ));
    InMux I__4757 (
            .O(N__21084),
            .I(N__21081));
    LocalMux I__4756 (
            .O(N__21081),
            .I(N__21078));
    Span12Mux_v I__4755 (
            .O(N__21078),
            .I(N__21075));
    Odrv12 I__4754 (
            .O(N__21075),
            .I(\line_buffer.n533 ));
    InMux I__4753 (
            .O(N__21072),
            .I(N__21069));
    LocalMux I__4752 (
            .O(N__21069),
            .I(N__21066));
    Span4Mux_h I__4751 (
            .O(N__21066),
            .I(N__21063));
    Span4Mux_h I__4750 (
            .O(N__21063),
            .I(N__21060));
    Odrv4 I__4749 (
            .O(N__21060),
            .I(\line_buffer.n525 ));
    InMux I__4748 (
            .O(N__21057),
            .I(N__21054));
    LocalMux I__4747 (
            .O(N__21054),
            .I(N__21046));
    InMux I__4746 (
            .O(N__21053),
            .I(N__21043));
    InMux I__4745 (
            .O(N__21052),
            .I(N__21040));
    InMux I__4744 (
            .O(N__21051),
            .I(N__21037));
    InMux I__4743 (
            .O(N__21050),
            .I(N__21034));
    InMux I__4742 (
            .O(N__21049),
            .I(N__21030));
    Span4Mux_h I__4741 (
            .O(N__21046),
            .I(N__21026));
    LocalMux I__4740 (
            .O(N__21043),
            .I(N__21017));
    LocalMux I__4739 (
            .O(N__21040),
            .I(N__21017));
    LocalMux I__4738 (
            .O(N__21037),
            .I(N__21017));
    LocalMux I__4737 (
            .O(N__21034),
            .I(N__21017));
    InMux I__4736 (
            .O(N__21033),
            .I(N__21014));
    LocalMux I__4735 (
            .O(N__21030),
            .I(N__21011));
    InMux I__4734 (
            .O(N__21029),
            .I(N__21008));
    Span4Mux_h I__4733 (
            .O(N__21026),
            .I(N__21004));
    Span12Mux_v I__4732 (
            .O(N__21017),
            .I(N__20999));
    LocalMux I__4731 (
            .O(N__21014),
            .I(N__20999));
    Span4Mux_s1_v I__4730 (
            .O(N__21011),
            .I(N__20994));
    LocalMux I__4729 (
            .O(N__21008),
            .I(N__20994));
    InMux I__4728 (
            .O(N__21007),
            .I(N__20991));
    Sp12to4 I__4727 (
            .O(N__21004),
            .I(N__20988));
    Span12Mux_v I__4726 (
            .O(N__20999),
            .I(N__20985));
    Span4Mux_v I__4725 (
            .O(N__20994),
            .I(N__20982));
    LocalMux I__4724 (
            .O(N__20991),
            .I(N__20979));
    Span12Mux_v I__4723 (
            .O(N__20988),
            .I(N__20974));
    Span12Mux_h I__4722 (
            .O(N__20985),
            .I(N__20974));
    Span4Mux_h I__4721 (
            .O(N__20982),
            .I(N__20971));
    Span4Mux_h I__4720 (
            .O(N__20979),
            .I(N__20968));
    Odrv12 I__4719 (
            .O(N__20974),
            .I(RX_DATA_7));
    Odrv4 I__4718 (
            .O(N__20971),
            .I(RX_DATA_7));
    Odrv4 I__4717 (
            .O(N__20968),
            .I(RX_DATA_7));
    InMux I__4716 (
            .O(N__20961),
            .I(N__20958));
    LocalMux I__4715 (
            .O(N__20958),
            .I(N__20955));
    Span12Mux_v I__4714 (
            .O(N__20955),
            .I(N__20952));
    Odrv12 I__4713 (
            .O(N__20952),
            .I(\line_buffer.n565 ));
    InMux I__4712 (
            .O(N__20949),
            .I(N__20946));
    LocalMux I__4711 (
            .O(N__20946),
            .I(N__20943));
    Span4Mux_h I__4710 (
            .O(N__20943),
            .I(N__20940));
    Span4Mux_h I__4709 (
            .O(N__20940),
            .I(N__20937));
    Odrv4 I__4708 (
            .O(N__20937),
            .I(\line_buffer.n557 ));
    CascadeMux I__4707 (
            .O(N__20934),
            .I(\line_buffer.n3656_cascade_ ));
    InMux I__4706 (
            .O(N__20931),
            .I(N__20928));
    LocalMux I__4705 (
            .O(N__20928),
            .I(\line_buffer.n3596 ));
    InMux I__4704 (
            .O(N__20925),
            .I(N__20922));
    LocalMux I__4703 (
            .O(N__20922),
            .I(\line_buffer.n3638 ));
    InMux I__4702 (
            .O(N__20919),
            .I(N__20916));
    LocalMux I__4701 (
            .O(N__20916),
            .I(N__20913));
    Span4Mux_v I__4700 (
            .O(N__20913),
            .I(N__20910));
    Odrv4 I__4699 (
            .O(N__20910),
            .I(TX_DATA_0));
    InMux I__4698 (
            .O(N__20907),
            .I(N__20904));
    LocalMux I__4697 (
            .O(N__20904),
            .I(N__20901));
    Span4Mux_v I__4696 (
            .O(N__20901),
            .I(N__20898));
    Sp12to4 I__4695 (
            .O(N__20898),
            .I(N__20895));
    Span12Mux_h I__4694 (
            .O(N__20895),
            .I(N__20892));
    Span12Mux_v I__4693 (
            .O(N__20892),
            .I(N__20889));
    Odrv12 I__4692 (
            .O(N__20889),
            .I(\line_buffer.n530 ));
    CascadeMux I__4691 (
            .O(N__20886),
            .I(N__20883));
    InMux I__4690 (
            .O(N__20883),
            .I(N__20880));
    LocalMux I__4689 (
            .O(N__20880),
            .I(N__20877));
    Span4Mux_h I__4688 (
            .O(N__20877),
            .I(N__20874));
    Span4Mux_h I__4687 (
            .O(N__20874),
            .I(N__20871));
    Span4Mux_v I__4686 (
            .O(N__20871),
            .I(N__20868));
    Odrv4 I__4685 (
            .O(N__20868),
            .I(\line_buffer.n522 ));
    InMux I__4684 (
            .O(N__20865),
            .I(N__20862));
    LocalMux I__4683 (
            .O(N__20862),
            .I(\line_buffer.n3632 ));
    CascadeMux I__4682 (
            .O(N__20859),
            .I(\line_buffer.n3650_cascade_ ));
    InMux I__4681 (
            .O(N__20856),
            .I(N__20853));
    LocalMux I__4680 (
            .O(N__20853),
            .I(N__20850));
    Span12Mux_h I__4679 (
            .O(N__20850),
            .I(N__20847));
    Odrv12 I__4678 (
            .O(N__20847),
            .I(\line_buffer.n594 ));
    InMux I__4677 (
            .O(N__20844),
            .I(N__20841));
    LocalMux I__4676 (
            .O(N__20841),
            .I(N__20838));
    Span12Mux_h I__4675 (
            .O(N__20838),
            .I(N__20835));
    Span12Mux_v I__4674 (
            .O(N__20835),
            .I(N__20832));
    Odrv12 I__4673 (
            .O(N__20832),
            .I(\line_buffer.n586 ));
    InMux I__4672 (
            .O(N__20829),
            .I(N__20826));
    LocalMux I__4671 (
            .O(N__20826),
            .I(\line_buffer.n3647 ));
    InMux I__4670 (
            .O(N__20823),
            .I(N__20820));
    LocalMux I__4669 (
            .O(N__20820),
            .I(N__20817));
    Span4Mux_h I__4668 (
            .O(N__20817),
            .I(N__20814));
    Span4Mux_h I__4667 (
            .O(N__20814),
            .I(N__20811));
    Span4Mux_v I__4666 (
            .O(N__20811),
            .I(N__20808));
    Odrv4 I__4665 (
            .O(N__20808),
            .I(\line_buffer.n521 ));
    CascadeMux I__4664 (
            .O(N__20805),
            .I(N__20802));
    InMux I__4663 (
            .O(N__20802),
            .I(N__20799));
    LocalMux I__4662 (
            .O(N__20799),
            .I(N__20796));
    Span4Mux_v I__4661 (
            .O(N__20796),
            .I(N__20793));
    Sp12to4 I__4660 (
            .O(N__20793),
            .I(N__20790));
    Span12Mux_h I__4659 (
            .O(N__20790),
            .I(N__20787));
    Span12Mux_v I__4658 (
            .O(N__20787),
            .I(N__20784));
    Odrv12 I__4657 (
            .O(N__20784),
            .I(\line_buffer.n529 ));
    InMux I__4656 (
            .O(N__20781),
            .I(N__20778));
    LocalMux I__4655 (
            .O(N__20778),
            .I(\line_buffer.n3644 ));
    InMux I__4654 (
            .O(N__20775),
            .I(N__20772));
    LocalMux I__4653 (
            .O(N__20772),
            .I(N__20769));
    Odrv12 I__4652 (
            .O(N__20769),
            .I(TX_DATA_5));
    IoInMux I__4651 (
            .O(N__20766),
            .I(N__20763));
    LocalMux I__4650 (
            .O(N__20763),
            .I(N__20759));
    IoInMux I__4649 (
            .O(N__20762),
            .I(N__20756));
    Span4Mux_s0_h I__4648 (
            .O(N__20759),
            .I(N__20753));
    LocalMux I__4647 (
            .O(N__20756),
            .I(N__20750));
    Span4Mux_h I__4646 (
            .O(N__20753),
            .I(N__20747));
    Span4Mux_s3_v I__4645 (
            .O(N__20750),
            .I(N__20744));
    Span4Mux_h I__4644 (
            .O(N__20747),
            .I(N__20740));
    Span4Mux_h I__4643 (
            .O(N__20744),
            .I(N__20737));
    IoInMux I__4642 (
            .O(N__20743),
            .I(N__20734));
    Span4Mux_h I__4641 (
            .O(N__20740),
            .I(N__20731));
    Span4Mux_h I__4640 (
            .O(N__20737),
            .I(N__20728));
    LocalMux I__4639 (
            .O(N__20734),
            .I(N__20725));
    Span4Mux_h I__4638 (
            .O(N__20731),
            .I(N__20720));
    Span4Mux_v I__4637 (
            .O(N__20728),
            .I(N__20720));
    Span12Mux_s11_v I__4636 (
            .O(N__20725),
            .I(N__20717));
    Span4Mux_v I__4635 (
            .O(N__20720),
            .I(N__20714));
    Odrv12 I__4634 (
            .O(N__20717),
            .I(n1813));
    Odrv4 I__4633 (
            .O(N__20714),
            .I(n1813));
    InMux I__4632 (
            .O(N__20709),
            .I(N__20706));
    LocalMux I__4631 (
            .O(N__20706),
            .I(N__20703));
    Odrv12 I__4630 (
            .O(N__20703),
            .I(TX_DATA_1));
    IoInMux I__4629 (
            .O(N__20700),
            .I(N__20697));
    LocalMux I__4628 (
            .O(N__20697),
            .I(N__20693));
    IoInMux I__4627 (
            .O(N__20696),
            .I(N__20690));
    Span4Mux_s1_v I__4626 (
            .O(N__20693),
            .I(N__20687));
    LocalMux I__4625 (
            .O(N__20690),
            .I(N__20684));
    Span4Mux_v I__4624 (
            .O(N__20687),
            .I(N__20679));
    Span4Mux_s2_h I__4623 (
            .O(N__20684),
            .I(N__20679));
    Span4Mux_h I__4622 (
            .O(N__20679),
            .I(N__20675));
    IoInMux I__4621 (
            .O(N__20678),
            .I(N__20672));
    Sp12to4 I__4620 (
            .O(N__20675),
            .I(N__20669));
    LocalMux I__4619 (
            .O(N__20672),
            .I(N__20666));
    Span12Mux_s10_v I__4618 (
            .O(N__20669),
            .I(N__20661));
    Span12Mux_s10_v I__4617 (
            .O(N__20666),
            .I(N__20661));
    Odrv12 I__4616 (
            .O(N__20661),
            .I(n1817));
    InMux I__4615 (
            .O(N__20658),
            .I(N__20655));
    LocalMux I__4614 (
            .O(N__20655),
            .I(\transmit_module.Y_DELTA_PATTERN_97 ));
    InMux I__4613 (
            .O(N__20652),
            .I(N__20649));
    LocalMux I__4612 (
            .O(N__20649),
            .I(\transmit_module.Y_DELTA_PATTERN_92 ));
    InMux I__4611 (
            .O(N__20646),
            .I(N__20643));
    LocalMux I__4610 (
            .O(N__20643),
            .I(\transmit_module.Y_DELTA_PATTERN_91 ));
    InMux I__4609 (
            .O(N__20640),
            .I(N__20637));
    LocalMux I__4608 (
            .O(N__20637),
            .I(\transmit_module.Y_DELTA_PATTERN_90 ));
    InMux I__4607 (
            .O(N__20634),
            .I(N__20630));
    InMux I__4606 (
            .O(N__20633),
            .I(N__20622));
    LocalMux I__4605 (
            .O(N__20630),
            .I(N__20619));
    InMux I__4604 (
            .O(N__20629),
            .I(N__20614));
    InMux I__4603 (
            .O(N__20628),
            .I(N__20614));
    InMux I__4602 (
            .O(N__20627),
            .I(N__20609));
    InMux I__4601 (
            .O(N__20626),
            .I(N__20609));
    InMux I__4600 (
            .O(N__20625),
            .I(N__20606));
    LocalMux I__4599 (
            .O(N__20622),
            .I(N__20601));
    Span4Mux_h I__4598 (
            .O(N__20619),
            .I(N__20596));
    LocalMux I__4597 (
            .O(N__20614),
            .I(N__20596));
    LocalMux I__4596 (
            .O(N__20609),
            .I(N__20593));
    LocalMux I__4595 (
            .O(N__20606),
            .I(N__20587));
    InMux I__4594 (
            .O(N__20605),
            .I(N__20584));
    InMux I__4593 (
            .O(N__20604),
            .I(N__20581));
    Span4Mux_h I__4592 (
            .O(N__20601),
            .I(N__20576));
    Span4Mux_h I__4591 (
            .O(N__20596),
            .I(N__20573));
    Span4Mux_h I__4590 (
            .O(N__20593),
            .I(N__20570));
    InMux I__4589 (
            .O(N__20592),
            .I(N__20567));
    InMux I__4588 (
            .O(N__20591),
            .I(N__20564));
    InMux I__4587 (
            .O(N__20590),
            .I(N__20561));
    Span4Mux_v I__4586 (
            .O(N__20587),
            .I(N__20554));
    LocalMux I__4585 (
            .O(N__20584),
            .I(N__20554));
    LocalMux I__4584 (
            .O(N__20581),
            .I(N__20554));
    InMux I__4583 (
            .O(N__20580),
            .I(N__20549));
    InMux I__4582 (
            .O(N__20579),
            .I(N__20549));
    Odrv4 I__4581 (
            .O(N__20576),
            .I(\transmit_module.Y_DELTA_PATTERN_0 ));
    Odrv4 I__4580 (
            .O(N__20573),
            .I(\transmit_module.Y_DELTA_PATTERN_0 ));
    Odrv4 I__4579 (
            .O(N__20570),
            .I(\transmit_module.Y_DELTA_PATTERN_0 ));
    LocalMux I__4578 (
            .O(N__20567),
            .I(\transmit_module.Y_DELTA_PATTERN_0 ));
    LocalMux I__4577 (
            .O(N__20564),
            .I(\transmit_module.Y_DELTA_PATTERN_0 ));
    LocalMux I__4576 (
            .O(N__20561),
            .I(\transmit_module.Y_DELTA_PATTERN_0 ));
    Odrv4 I__4575 (
            .O(N__20554),
            .I(\transmit_module.Y_DELTA_PATTERN_0 ));
    LocalMux I__4574 (
            .O(N__20549),
            .I(\transmit_module.Y_DELTA_PATTERN_0 ));
    InMux I__4573 (
            .O(N__20532),
            .I(N__20529));
    LocalMux I__4572 (
            .O(N__20529),
            .I(\transmit_module.Y_DELTA_PATTERN_99 ));
    CEMux I__4571 (
            .O(N__20526),
            .I(N__20522));
    CEMux I__4570 (
            .O(N__20525),
            .I(N__20519));
    LocalMux I__4569 (
            .O(N__20522),
            .I(N__20511));
    LocalMux I__4568 (
            .O(N__20519),
            .I(N__20507));
    CEMux I__4567 (
            .O(N__20518),
            .I(N__20504));
    CEMux I__4566 (
            .O(N__20517),
            .I(N__20500));
    CEMux I__4565 (
            .O(N__20516),
            .I(N__20496));
    SRMux I__4564 (
            .O(N__20515),
            .I(N__20493));
    CEMux I__4563 (
            .O(N__20514),
            .I(N__20489));
    Span4Mux_v I__4562 (
            .O(N__20511),
            .I(N__20483));
    CEMux I__4561 (
            .O(N__20510),
            .I(N__20480));
    Span4Mux_v I__4560 (
            .O(N__20507),
            .I(N__20475));
    LocalMux I__4559 (
            .O(N__20504),
            .I(N__20475));
    CEMux I__4558 (
            .O(N__20503),
            .I(N__20472));
    LocalMux I__4557 (
            .O(N__20500),
            .I(N__20469));
    CEMux I__4556 (
            .O(N__20499),
            .I(N__20466));
    LocalMux I__4555 (
            .O(N__20496),
            .I(N__20463));
    LocalMux I__4554 (
            .O(N__20493),
            .I(N__20460));
    SRMux I__4553 (
            .O(N__20492),
            .I(N__20457));
    LocalMux I__4552 (
            .O(N__20489),
            .I(N__20454));
    CEMux I__4551 (
            .O(N__20488),
            .I(N__20451));
    CEMux I__4550 (
            .O(N__20487),
            .I(N__20448));
    SRMux I__4549 (
            .O(N__20486),
            .I(N__20445));
    Span4Mux_v I__4548 (
            .O(N__20483),
            .I(N__20440));
    LocalMux I__4547 (
            .O(N__20480),
            .I(N__20440));
    Span4Mux_h I__4546 (
            .O(N__20475),
            .I(N__20437));
    LocalMux I__4545 (
            .O(N__20472),
            .I(N__20434));
    Span4Mux_v I__4544 (
            .O(N__20469),
            .I(N__20429));
    LocalMux I__4543 (
            .O(N__20466),
            .I(N__20429));
    Span4Mux_v I__4542 (
            .O(N__20463),
            .I(N__20426));
    Span4Mux_v I__4541 (
            .O(N__20460),
            .I(N__20423));
    LocalMux I__4540 (
            .O(N__20457),
            .I(N__20420));
    Span4Mux_h I__4539 (
            .O(N__20454),
            .I(N__20414));
    LocalMux I__4538 (
            .O(N__20451),
            .I(N__20414));
    LocalMux I__4537 (
            .O(N__20448),
            .I(N__20411));
    LocalMux I__4536 (
            .O(N__20445),
            .I(N__20408));
    Span4Mux_v I__4535 (
            .O(N__20440),
            .I(N__20405));
    Span4Mux_h I__4534 (
            .O(N__20437),
            .I(N__20400));
    Span4Mux_v I__4533 (
            .O(N__20434),
            .I(N__20400));
    Span4Mux_h I__4532 (
            .O(N__20429),
            .I(N__20391));
    Span4Mux_h I__4531 (
            .O(N__20426),
            .I(N__20391));
    Span4Mux_h I__4530 (
            .O(N__20423),
            .I(N__20391));
    Span4Mux_v I__4529 (
            .O(N__20420),
            .I(N__20391));
    SRMux I__4528 (
            .O(N__20419),
            .I(N__20388));
    Span4Mux_h I__4527 (
            .O(N__20414),
            .I(N__20381));
    Span4Mux_v I__4526 (
            .O(N__20411),
            .I(N__20381));
    Span4Mux_h I__4525 (
            .O(N__20408),
            .I(N__20381));
    Odrv4 I__4524 (
            .O(N__20405),
            .I(\transmit_module.n3679 ));
    Odrv4 I__4523 (
            .O(N__20400),
            .I(\transmit_module.n3679 ));
    Odrv4 I__4522 (
            .O(N__20391),
            .I(\transmit_module.n3679 ));
    LocalMux I__4521 (
            .O(N__20388),
            .I(\transmit_module.n3679 ));
    Odrv4 I__4520 (
            .O(N__20381),
            .I(\transmit_module.n3679 ));
    InMux I__4519 (
            .O(N__20370),
            .I(N__20367));
    LocalMux I__4518 (
            .O(N__20367),
            .I(N__20364));
    Span4Mux_v I__4517 (
            .O(N__20364),
            .I(N__20361));
    Span4Mux_v I__4516 (
            .O(N__20361),
            .I(N__20358));
    Sp12to4 I__4515 (
            .O(N__20358),
            .I(N__20355));
    Odrv12 I__4514 (
            .O(N__20355),
            .I(\line_buffer.n566 ));
    InMux I__4513 (
            .O(N__20352),
            .I(N__20349));
    LocalMux I__4512 (
            .O(N__20349),
            .I(N__20346));
    Span4Mux_h I__4511 (
            .O(N__20346),
            .I(N__20343));
    Span4Mux_h I__4510 (
            .O(N__20343),
            .I(N__20340));
    Odrv4 I__4509 (
            .O(N__20340),
            .I(\line_buffer.n558 ));
    InMux I__4508 (
            .O(N__20337),
            .I(N__20334));
    LocalMux I__4507 (
            .O(N__20334),
            .I(N__20331));
    Span4Mux_h I__4506 (
            .O(N__20331),
            .I(N__20328));
    Span4Mux_v I__4505 (
            .O(N__20328),
            .I(N__20325));
    Span4Mux_h I__4504 (
            .O(N__20325),
            .I(N__20322));
    Odrv4 I__4503 (
            .O(N__20322),
            .I(\line_buffer.n465 ));
    CascadeMux I__4502 (
            .O(N__20319),
            .I(N__20316));
    InMux I__4501 (
            .O(N__20316),
            .I(N__20313));
    LocalMux I__4500 (
            .O(N__20313),
            .I(N__20310));
    Span12Mux_h I__4499 (
            .O(N__20310),
            .I(N__20307));
    Span12Mux_v I__4498 (
            .O(N__20307),
            .I(N__20304));
    Odrv12 I__4497 (
            .O(N__20304),
            .I(\line_buffer.n457 ));
    InMux I__4496 (
            .O(N__20301),
            .I(N__20298));
    LocalMux I__4495 (
            .O(N__20298),
            .I(\line_buffer.n3629 ));
    InMux I__4494 (
            .O(N__20295),
            .I(N__20292));
    LocalMux I__4493 (
            .O(N__20292),
            .I(N__20289));
    Span4Mux_v I__4492 (
            .O(N__20289),
            .I(N__20286));
    Span4Mux_v I__4491 (
            .O(N__20286),
            .I(N__20283));
    Sp12to4 I__4490 (
            .O(N__20283),
            .I(N__20280));
    Odrv12 I__4489 (
            .O(N__20280),
            .I(\line_buffer.n561 ));
    InMux I__4488 (
            .O(N__20277),
            .I(N__20274));
    LocalMux I__4487 (
            .O(N__20274),
            .I(N__20271));
    Span4Mux_h I__4486 (
            .O(N__20271),
            .I(N__20268));
    Span4Mux_h I__4485 (
            .O(N__20268),
            .I(N__20265));
    Odrv4 I__4484 (
            .O(N__20265),
            .I(\line_buffer.n553 ));
    InMux I__4483 (
            .O(N__20262),
            .I(N__20259));
    LocalMux I__4482 (
            .O(N__20259),
            .I(N__20256));
    Span4Mux_h I__4481 (
            .O(N__20256),
            .I(N__20253));
    Span4Mux_h I__4480 (
            .O(N__20253),
            .I(N__20250));
    Span4Mux_v I__4479 (
            .O(N__20250),
            .I(N__20247));
    Span4Mux_v I__4478 (
            .O(N__20247),
            .I(N__20244));
    Odrv4 I__4477 (
            .O(N__20244),
            .I(\line_buffer.n456 ));
    InMux I__4476 (
            .O(N__20241),
            .I(N__20238));
    LocalMux I__4475 (
            .O(N__20238),
            .I(N__20235));
    Span4Mux_v I__4474 (
            .O(N__20235),
            .I(N__20232));
    Span4Mux_h I__4473 (
            .O(N__20232),
            .I(N__20229));
    Span4Mux_h I__4472 (
            .O(N__20229),
            .I(N__20226));
    Odrv4 I__4471 (
            .O(N__20226),
            .I(\line_buffer.n464 ));
    CascadeMux I__4470 (
            .O(N__20223),
            .I(\line_buffer.n3635_cascade_ ));
    InMux I__4469 (
            .O(N__20220),
            .I(N__20217));
    LocalMux I__4468 (
            .O(N__20217),
            .I(N__20214));
    Span4Mux_h I__4467 (
            .O(N__20214),
            .I(N__20211));
    Span4Mux_h I__4466 (
            .O(N__20211),
            .I(N__20208));
    Odrv4 I__4465 (
            .O(N__20208),
            .I(\line_buffer.n469 ));
    InMux I__4464 (
            .O(N__20205),
            .I(N__20202));
    LocalMux I__4463 (
            .O(N__20202),
            .I(N__20199));
    Span12Mux_h I__4462 (
            .O(N__20199),
            .I(N__20196));
    Span12Mux_v I__4461 (
            .O(N__20196),
            .I(N__20193));
    Odrv12 I__4460 (
            .O(N__20193),
            .I(\line_buffer.n461 ));
    InMux I__4459 (
            .O(N__20190),
            .I(N__20187));
    LocalMux I__4458 (
            .O(N__20187),
            .I(N__20184));
    Odrv4 I__4457 (
            .O(N__20184),
            .I(\line_buffer.n3653 ));
    IoInMux I__4456 (
            .O(N__20181),
            .I(N__20178));
    LocalMux I__4455 (
            .O(N__20178),
            .I(N__20175));
    IoSpan4Mux I__4454 (
            .O(N__20175),
            .I(N__20172));
    Span4Mux_s2_h I__4453 (
            .O(N__20172),
            .I(N__20169));
    Span4Mux_h I__4452 (
            .O(N__20169),
            .I(N__20165));
    InMux I__4451 (
            .O(N__20168),
            .I(N__20162));
    Sp12to4 I__4450 (
            .O(N__20165),
            .I(N__20157));
    LocalMux I__4449 (
            .O(N__20162),
            .I(N__20157));
    Span12Mux_h I__4448 (
            .O(N__20157),
            .I(N__20154));
    Odrv12 I__4447 (
            .O(N__20154),
            .I(DEBUG_c_2_c));
    InMux I__4446 (
            .O(N__20151),
            .I(N__20148));
    LocalMux I__4445 (
            .O(N__20148),
            .I(\tvp_hs_buffer.BUFFER_0_0 ));
    InMux I__4444 (
            .O(N__20145),
            .I(N__20142));
    LocalMux I__4443 (
            .O(N__20142),
            .I(\tvp_hs_buffer.BUFFER_1_0 ));
    InMux I__4442 (
            .O(N__20139),
            .I(N__20126));
    InMux I__4441 (
            .O(N__20138),
            .I(N__20119));
    InMux I__4440 (
            .O(N__20137),
            .I(N__20119));
    InMux I__4439 (
            .O(N__20136),
            .I(N__20119));
    InMux I__4438 (
            .O(N__20135),
            .I(N__20112));
    InMux I__4437 (
            .O(N__20134),
            .I(N__20112));
    InMux I__4436 (
            .O(N__20133),
            .I(N__20112));
    InMux I__4435 (
            .O(N__20132),
            .I(N__20105));
    InMux I__4434 (
            .O(N__20131),
            .I(N__20105));
    InMux I__4433 (
            .O(N__20130),
            .I(N__20105));
    InMux I__4432 (
            .O(N__20129),
            .I(N__20101));
    LocalMux I__4431 (
            .O(N__20126),
            .I(N__20097));
    LocalMux I__4430 (
            .O(N__20119),
            .I(N__20089));
    LocalMux I__4429 (
            .O(N__20112),
            .I(N__20089));
    LocalMux I__4428 (
            .O(N__20105),
            .I(N__20089));
    InMux I__4427 (
            .O(N__20104),
            .I(N__20086));
    LocalMux I__4426 (
            .O(N__20101),
            .I(N__20083));
    InMux I__4425 (
            .O(N__20100),
            .I(N__20080));
    Span12Mux_s2_v I__4424 (
            .O(N__20097),
            .I(N__20076));
    InMux I__4423 (
            .O(N__20096),
            .I(N__20073));
    Span4Mux_v I__4422 (
            .O(N__20089),
            .I(N__20068));
    LocalMux I__4421 (
            .O(N__20086),
            .I(N__20068));
    Span4Mux_v I__4420 (
            .O(N__20083),
            .I(N__20063));
    LocalMux I__4419 (
            .O(N__20080),
            .I(N__20060));
    InMux I__4418 (
            .O(N__20079),
            .I(N__20057));
    Span12Mux_v I__4417 (
            .O(N__20076),
            .I(N__20051));
    LocalMux I__4416 (
            .O(N__20073),
            .I(N__20051));
    Span4Mux_v I__4415 (
            .O(N__20068),
            .I(N__20048));
    InMux I__4414 (
            .O(N__20067),
            .I(N__20043));
    InMux I__4413 (
            .O(N__20066),
            .I(N__20043));
    Span4Mux_v I__4412 (
            .O(N__20063),
            .I(N__20036));
    Span4Mux_v I__4411 (
            .O(N__20060),
            .I(N__20036));
    LocalMux I__4410 (
            .O(N__20057),
            .I(N__20036));
    InMux I__4409 (
            .O(N__20056),
            .I(N__20033));
    Odrv12 I__4408 (
            .O(N__20051),
            .I(TVP_VSYNC_buff));
    Odrv4 I__4407 (
            .O(N__20048),
            .I(TVP_VSYNC_buff));
    LocalMux I__4406 (
            .O(N__20043),
            .I(TVP_VSYNC_buff));
    Odrv4 I__4405 (
            .O(N__20036),
            .I(TVP_VSYNC_buff));
    LocalMux I__4404 (
            .O(N__20033),
            .I(TVP_VSYNC_buff));
    CEMux I__4403 (
            .O(N__20022),
            .I(N__20019));
    LocalMux I__4402 (
            .O(N__20019),
            .I(N__20015));
    CEMux I__4401 (
            .O(N__20018),
            .I(N__20012));
    Span4Mux_h I__4400 (
            .O(N__20015),
            .I(N__20009));
    LocalMux I__4399 (
            .O(N__20012),
            .I(N__20006));
    Odrv4 I__4398 (
            .O(N__20009),
            .I(\receive_module.rx_counter.n2078 ));
    Odrv12 I__4397 (
            .O(N__20006),
            .I(\receive_module.rx_counter.n2078 ));
    InMux I__4396 (
            .O(N__20001),
            .I(N__19996));
    InMux I__4395 (
            .O(N__20000),
            .I(N__19991));
    InMux I__4394 (
            .O(N__19999),
            .I(N__19991));
    LocalMux I__4393 (
            .O(N__19996),
            .I(N__19988));
    LocalMux I__4392 (
            .O(N__19991),
            .I(TVP_HSYNC_buff));
    Odrv4 I__4391 (
            .O(N__19988),
            .I(TVP_HSYNC_buff));
    InMux I__4390 (
            .O(N__19983),
            .I(N__19980));
    LocalMux I__4389 (
            .O(N__19980),
            .I(\receive_module.rx_counter.old_HS ));
    InMux I__4388 (
            .O(N__19977),
            .I(N__19974));
    LocalMux I__4387 (
            .O(N__19974),
            .I(\transmit_module.Y_DELTA_PATTERN_98 ));
    InMux I__4386 (
            .O(N__19971),
            .I(N__19968));
    LocalMux I__4385 (
            .O(N__19968),
            .I(\transmit_module.Y_DELTA_PATTERN_89 ));
    IoInMux I__4384 (
            .O(N__19965),
            .I(N__19962));
    LocalMux I__4383 (
            .O(N__19962),
            .I(N__19959));
    IoSpan4Mux I__4382 (
            .O(N__19959),
            .I(N__19956));
    Span4Mux_s3_h I__4381 (
            .O(N__19956),
            .I(N__19952));
    InMux I__4380 (
            .O(N__19955),
            .I(N__19949));
    Sp12to4 I__4379 (
            .O(N__19952),
            .I(N__19946));
    LocalMux I__4378 (
            .O(N__19949),
            .I(N__19943));
    Span12Mux_v I__4377 (
            .O(N__19946),
            .I(N__19940));
    Span12Mux_h I__4376 (
            .O(N__19943),
            .I(N__19937));
    Span12Mux_h I__4375 (
            .O(N__19940),
            .I(N__19934));
    Span12Mux_v I__4374 (
            .O(N__19937),
            .I(N__19931));
    Odrv12 I__4373 (
            .O(N__19934),
            .I(DEBUG_c_7_c));
    Odrv12 I__4372 (
            .O(N__19931),
            .I(DEBUG_c_7_c));
    InMux I__4371 (
            .O(N__19926),
            .I(N__19923));
    LocalMux I__4370 (
            .O(N__19923),
            .I(N__19918));
    InMux I__4369 (
            .O(N__19922),
            .I(N__19915));
    InMux I__4368 (
            .O(N__19921),
            .I(N__19911));
    Span4Mux_s2_v I__4367 (
            .O(N__19918),
            .I(N__19904));
    LocalMux I__4366 (
            .O(N__19915),
            .I(N__19904));
    InMux I__4365 (
            .O(N__19914),
            .I(N__19901));
    LocalMux I__4364 (
            .O(N__19911),
            .I(N__19898));
    InMux I__4363 (
            .O(N__19910),
            .I(N__19895));
    InMux I__4362 (
            .O(N__19909),
            .I(N__19892));
    Span4Mux_v I__4361 (
            .O(N__19904),
            .I(N__19888));
    LocalMux I__4360 (
            .O(N__19901),
            .I(N__19885));
    Span4Mux_v I__4359 (
            .O(N__19898),
            .I(N__19878));
    LocalMux I__4358 (
            .O(N__19895),
            .I(N__19878));
    LocalMux I__4357 (
            .O(N__19892),
            .I(N__19878));
    InMux I__4356 (
            .O(N__19891),
            .I(N__19875));
    Span4Mux_h I__4355 (
            .O(N__19888),
            .I(N__19870));
    Span4Mux_v I__4354 (
            .O(N__19885),
            .I(N__19867));
    Span4Mux_v I__4353 (
            .O(N__19878),
            .I(N__19862));
    LocalMux I__4352 (
            .O(N__19875),
            .I(N__19862));
    InMux I__4351 (
            .O(N__19874),
            .I(N__19859));
    InMux I__4350 (
            .O(N__19873),
            .I(N__19856));
    Sp12to4 I__4349 (
            .O(N__19870),
            .I(N__19853));
    Span4Mux_h I__4348 (
            .O(N__19867),
            .I(N__19850));
    Span4Mux_v I__4347 (
            .O(N__19862),
            .I(N__19845));
    LocalMux I__4346 (
            .O(N__19859),
            .I(N__19845));
    LocalMux I__4345 (
            .O(N__19856),
            .I(N__19842));
    Span12Mux_v I__4344 (
            .O(N__19853),
            .I(N__19837));
    Sp12to4 I__4343 (
            .O(N__19850),
            .I(N__19837));
    Span4Mux_v I__4342 (
            .O(N__19845),
            .I(N__19834));
    Span4Mux_h I__4341 (
            .O(N__19842),
            .I(N__19831));
    Span12Mux_v I__4340 (
            .O(N__19837),
            .I(N__19826));
    Sp12to4 I__4339 (
            .O(N__19834),
            .I(N__19826));
    Span4Mux_v I__4338 (
            .O(N__19831),
            .I(N__19823));
    Odrv12 I__4337 (
            .O(N__19826),
            .I(RX_DATA_6));
    Odrv4 I__4336 (
            .O(N__19823),
            .I(RX_DATA_6));
    InMux I__4335 (
            .O(N__19818),
            .I(N__19815));
    LocalMux I__4334 (
            .O(N__19815),
            .I(\tvp_video_buffer.BUFFER_0_8 ));
    InMux I__4333 (
            .O(N__19812),
            .I(N__19809));
    LocalMux I__4332 (
            .O(N__19809),
            .I(\tvp_video_buffer.BUFFER_1_8 ));
    InMux I__4331 (
            .O(N__19806),
            .I(N__19803));
    LocalMux I__4330 (
            .O(N__19803),
            .I(N__19800));
    Span4Mux_v I__4329 (
            .O(N__19800),
            .I(N__19797));
    Sp12to4 I__4328 (
            .O(N__19797),
            .I(N__19794));
    Odrv12 I__4327 (
            .O(N__19794),
            .I(\line_buffer.n598 ));
    InMux I__4326 (
            .O(N__19791),
            .I(N__19788));
    LocalMux I__4325 (
            .O(N__19788),
            .I(N__19785));
    Span12Mux_v I__4324 (
            .O(N__19785),
            .I(N__19782));
    Odrv12 I__4323 (
            .O(N__19782),
            .I(\line_buffer.n590 ));
    InMux I__4322 (
            .O(N__19779),
            .I(N__19776));
    LocalMux I__4321 (
            .O(N__19776),
            .I(N__19773));
    Sp12to4 I__4320 (
            .O(N__19773),
            .I(N__19770));
    Span12Mux_v I__4319 (
            .O(N__19770),
            .I(N__19767));
    Odrv12 I__4318 (
            .O(N__19767),
            .I(\line_buffer.n526 ));
    InMux I__4317 (
            .O(N__19764),
            .I(N__19761));
    LocalMux I__4316 (
            .O(N__19761),
            .I(N__19758));
    Span4Mux_v I__4315 (
            .O(N__19758),
            .I(N__19755));
    Sp12to4 I__4314 (
            .O(N__19755),
            .I(N__19752));
    Span12Mux_h I__4313 (
            .O(N__19752),
            .I(N__19749));
    Span12Mux_v I__4312 (
            .O(N__19749),
            .I(N__19746));
    Odrv12 I__4311 (
            .O(N__19746),
            .I(\line_buffer.n534 ));
    CascadeMux I__4310 (
            .O(N__19743),
            .I(\line_buffer.n3593_cascade_ ));
    InMux I__4309 (
            .O(N__19740),
            .I(N__19737));
    LocalMux I__4308 (
            .O(N__19737),
            .I(N__19734));
    Odrv12 I__4307 (
            .O(N__19734),
            .I(\line_buffer.n554 ));
    InMux I__4306 (
            .O(N__19731),
            .I(N__19728));
    LocalMux I__4305 (
            .O(N__19728),
            .I(N__19725));
    Span4Mux_v I__4304 (
            .O(N__19725),
            .I(N__19722));
    Span4Mux_h I__4303 (
            .O(N__19722),
            .I(N__19719));
    Span4Mux_h I__4302 (
            .O(N__19719),
            .I(N__19716));
    Odrv4 I__4301 (
            .O(N__19716),
            .I(\line_buffer.n562 ));
    InMux I__4300 (
            .O(N__19713),
            .I(N__19710));
    LocalMux I__4299 (
            .O(N__19710),
            .I(N__19707));
    Span4Mux_h I__4298 (
            .O(N__19707),
            .I(N__19704));
    Odrv4 I__4297 (
            .O(N__19704),
            .I(\receive_module.n132 ));
    IoInMux I__4296 (
            .O(N__19701),
            .I(N__19698));
    LocalMux I__4295 (
            .O(N__19698),
            .I(N__19694));
    CascadeMux I__4294 (
            .O(N__19697),
            .I(N__19691));
    Span4Mux_s3_h I__4293 (
            .O(N__19694),
            .I(N__19687));
    InMux I__4292 (
            .O(N__19691),
            .I(N__19681));
    CascadeMux I__4291 (
            .O(N__19690),
            .I(N__19677));
    Span4Mux_h I__4290 (
            .O(N__19687),
            .I(N__19673));
    CascadeMux I__4289 (
            .O(N__19686),
            .I(N__19664));
    CascadeMux I__4288 (
            .O(N__19685),
            .I(N__19661));
    CascadeMux I__4287 (
            .O(N__19684),
            .I(N__19656));
    LocalMux I__4286 (
            .O(N__19681),
            .I(N__19653));
    InMux I__4285 (
            .O(N__19680),
            .I(N__19650));
    InMux I__4284 (
            .O(N__19677),
            .I(N__19646));
    CascadeMux I__4283 (
            .O(N__19676),
            .I(N__19642));
    Span4Mux_h I__4282 (
            .O(N__19673),
            .I(N__19638));
    InMux I__4281 (
            .O(N__19672),
            .I(N__19631));
    InMux I__4280 (
            .O(N__19671),
            .I(N__19631));
    InMux I__4279 (
            .O(N__19670),
            .I(N__19631));
    InMux I__4278 (
            .O(N__19669),
            .I(N__19626));
    InMux I__4277 (
            .O(N__19668),
            .I(N__19626));
    InMux I__4276 (
            .O(N__19667),
            .I(N__19613));
    InMux I__4275 (
            .O(N__19664),
            .I(N__19613));
    InMux I__4274 (
            .O(N__19661),
            .I(N__19613));
    InMux I__4273 (
            .O(N__19660),
            .I(N__19613));
    InMux I__4272 (
            .O(N__19659),
            .I(N__19613));
    InMux I__4271 (
            .O(N__19656),
            .I(N__19613));
    Sp12to4 I__4270 (
            .O(N__19653),
            .I(N__19608));
    LocalMux I__4269 (
            .O(N__19650),
            .I(N__19608));
    InMux I__4268 (
            .O(N__19649),
            .I(N__19605));
    LocalMux I__4267 (
            .O(N__19646),
            .I(N__19602));
    InMux I__4266 (
            .O(N__19645),
            .I(N__19595));
    InMux I__4265 (
            .O(N__19642),
            .I(N__19595));
    InMux I__4264 (
            .O(N__19641),
            .I(N__19595));
    Span4Mux_h I__4263 (
            .O(N__19638),
            .I(N__19586));
    LocalMux I__4262 (
            .O(N__19631),
            .I(N__19586));
    LocalMux I__4261 (
            .O(N__19626),
            .I(N__19583));
    LocalMux I__4260 (
            .O(N__19613),
            .I(N__19576));
    Span12Mux_v I__4259 (
            .O(N__19608),
            .I(N__19576));
    LocalMux I__4258 (
            .O(N__19605),
            .I(N__19576));
    Span4Mux_v I__4257 (
            .O(N__19602),
            .I(N__19571));
    LocalMux I__4256 (
            .O(N__19595),
            .I(N__19571));
    InMux I__4255 (
            .O(N__19594),
            .I(N__19568));
    InMux I__4254 (
            .O(N__19593),
            .I(N__19565));
    InMux I__4253 (
            .O(N__19592),
            .I(N__19560));
    InMux I__4252 (
            .O(N__19591),
            .I(N__19560));
    Span4Mux_v I__4251 (
            .O(N__19586),
            .I(N__19555));
    Span4Mux_v I__4250 (
            .O(N__19583),
            .I(N__19555));
    Odrv12 I__4249 (
            .O(N__19576),
            .I(DEBUG_c_4));
    Odrv4 I__4248 (
            .O(N__19571),
            .I(DEBUG_c_4));
    LocalMux I__4247 (
            .O(N__19568),
            .I(DEBUG_c_4));
    LocalMux I__4246 (
            .O(N__19565),
            .I(DEBUG_c_4));
    LocalMux I__4245 (
            .O(N__19560),
            .I(DEBUG_c_4));
    Odrv4 I__4244 (
            .O(N__19555),
            .I(DEBUG_c_4));
    CascadeMux I__4243 (
            .O(N__19542),
            .I(N__19538));
    CascadeMux I__4242 (
            .O(N__19541),
            .I(N__19535));
    CascadeBuf I__4241 (
            .O(N__19538),
            .I(N__19532));
    CascadeBuf I__4240 (
            .O(N__19535),
            .I(N__19529));
    CascadeMux I__4239 (
            .O(N__19532),
            .I(N__19526));
    CascadeMux I__4238 (
            .O(N__19529),
            .I(N__19523));
    CascadeBuf I__4237 (
            .O(N__19526),
            .I(N__19520));
    CascadeBuf I__4236 (
            .O(N__19523),
            .I(N__19517));
    CascadeMux I__4235 (
            .O(N__19520),
            .I(N__19514));
    CascadeMux I__4234 (
            .O(N__19517),
            .I(N__19511));
    CascadeBuf I__4233 (
            .O(N__19514),
            .I(N__19508));
    CascadeBuf I__4232 (
            .O(N__19511),
            .I(N__19505));
    CascadeMux I__4231 (
            .O(N__19508),
            .I(N__19502));
    CascadeMux I__4230 (
            .O(N__19505),
            .I(N__19499));
    CascadeBuf I__4229 (
            .O(N__19502),
            .I(N__19496));
    CascadeBuf I__4228 (
            .O(N__19499),
            .I(N__19493));
    CascadeMux I__4227 (
            .O(N__19496),
            .I(N__19490));
    CascadeMux I__4226 (
            .O(N__19493),
            .I(N__19487));
    CascadeBuf I__4225 (
            .O(N__19490),
            .I(N__19484));
    CascadeBuf I__4224 (
            .O(N__19487),
            .I(N__19481));
    CascadeMux I__4223 (
            .O(N__19484),
            .I(N__19478));
    CascadeMux I__4222 (
            .O(N__19481),
            .I(N__19475));
    CascadeBuf I__4221 (
            .O(N__19478),
            .I(N__19472));
    CascadeBuf I__4220 (
            .O(N__19475),
            .I(N__19469));
    CascadeMux I__4219 (
            .O(N__19472),
            .I(N__19466));
    CascadeMux I__4218 (
            .O(N__19469),
            .I(N__19463));
    CascadeBuf I__4217 (
            .O(N__19466),
            .I(N__19460));
    CascadeBuf I__4216 (
            .O(N__19463),
            .I(N__19457));
    CascadeMux I__4215 (
            .O(N__19460),
            .I(N__19454));
    CascadeMux I__4214 (
            .O(N__19457),
            .I(N__19451));
    CascadeBuf I__4213 (
            .O(N__19454),
            .I(N__19448));
    CascadeBuf I__4212 (
            .O(N__19451),
            .I(N__19445));
    CascadeMux I__4211 (
            .O(N__19448),
            .I(N__19442));
    CascadeMux I__4210 (
            .O(N__19445),
            .I(N__19439));
    CascadeBuf I__4209 (
            .O(N__19442),
            .I(N__19436));
    CascadeBuf I__4208 (
            .O(N__19439),
            .I(N__19433));
    CascadeMux I__4207 (
            .O(N__19436),
            .I(N__19430));
    CascadeMux I__4206 (
            .O(N__19433),
            .I(N__19427));
    CascadeBuf I__4205 (
            .O(N__19430),
            .I(N__19424));
    CascadeBuf I__4204 (
            .O(N__19427),
            .I(N__19421));
    CascadeMux I__4203 (
            .O(N__19424),
            .I(N__19418));
    CascadeMux I__4202 (
            .O(N__19421),
            .I(N__19415));
    CascadeBuf I__4201 (
            .O(N__19418),
            .I(N__19412));
    CascadeBuf I__4200 (
            .O(N__19415),
            .I(N__19409));
    CascadeMux I__4199 (
            .O(N__19412),
            .I(N__19406));
    CascadeMux I__4198 (
            .O(N__19409),
            .I(N__19403));
    CascadeBuf I__4197 (
            .O(N__19406),
            .I(N__19400));
    CascadeBuf I__4196 (
            .O(N__19403),
            .I(N__19397));
    CascadeMux I__4195 (
            .O(N__19400),
            .I(N__19394));
    CascadeMux I__4194 (
            .O(N__19397),
            .I(N__19391));
    CascadeBuf I__4193 (
            .O(N__19394),
            .I(N__19388));
    CascadeBuf I__4192 (
            .O(N__19391),
            .I(N__19385));
    CascadeMux I__4191 (
            .O(N__19388),
            .I(N__19382));
    CascadeMux I__4190 (
            .O(N__19385),
            .I(N__19379));
    CascadeBuf I__4189 (
            .O(N__19382),
            .I(N__19376));
    CascadeBuf I__4188 (
            .O(N__19379),
            .I(N__19373));
    CascadeMux I__4187 (
            .O(N__19376),
            .I(N__19370));
    CascadeMux I__4186 (
            .O(N__19373),
            .I(N__19367));
    CascadeBuf I__4185 (
            .O(N__19370),
            .I(N__19364));
    CascadeBuf I__4184 (
            .O(N__19367),
            .I(N__19361));
    CascadeMux I__4183 (
            .O(N__19364),
            .I(N__19358));
    CascadeMux I__4182 (
            .O(N__19361),
            .I(N__19355));
    InMux I__4181 (
            .O(N__19358),
            .I(N__19352));
    InMux I__4180 (
            .O(N__19355),
            .I(N__19349));
    LocalMux I__4179 (
            .O(N__19352),
            .I(N__19345));
    LocalMux I__4178 (
            .O(N__19349),
            .I(N__19342));
    InMux I__4177 (
            .O(N__19348),
            .I(N__19339));
    Span4Mux_h I__4176 (
            .O(N__19345),
            .I(N__19336));
    Span4Mux_s2_v I__4175 (
            .O(N__19342),
            .I(N__19333));
    LocalMux I__4174 (
            .O(N__19339),
            .I(N__19330));
    Sp12to4 I__4173 (
            .O(N__19336),
            .I(N__19326));
    Sp12to4 I__4172 (
            .O(N__19333),
            .I(N__19323));
    Span4Mux_h I__4171 (
            .O(N__19330),
            .I(N__19320));
    InMux I__4170 (
            .O(N__19329),
            .I(N__19317));
    Span12Mux_v I__4169 (
            .O(N__19326),
            .I(N__19314));
    Span12Mux_h I__4168 (
            .O(N__19323),
            .I(N__19311));
    Odrv4 I__4167 (
            .O(N__19320),
            .I(RX_ADDR_5));
    LocalMux I__4166 (
            .O(N__19317),
            .I(RX_ADDR_5));
    Odrv12 I__4165 (
            .O(N__19314),
            .I(RX_ADDR_5));
    Odrv12 I__4164 (
            .O(N__19311),
            .I(RX_ADDR_5));
    SRMux I__4163 (
            .O(N__19302),
            .I(N__19295));
    SRMux I__4162 (
            .O(N__19301),
            .I(N__19292));
    SRMux I__4161 (
            .O(N__19300),
            .I(N__19288));
    SRMux I__4160 (
            .O(N__19299),
            .I(N__19285));
    SRMux I__4159 (
            .O(N__19298),
            .I(N__19282));
    LocalMux I__4158 (
            .O(N__19295),
            .I(N__19279));
    LocalMux I__4157 (
            .O(N__19292),
            .I(N__19276));
    SRMux I__4156 (
            .O(N__19291),
            .I(N__19273));
    LocalMux I__4155 (
            .O(N__19288),
            .I(N__19269));
    LocalMux I__4154 (
            .O(N__19285),
            .I(N__19266));
    LocalMux I__4153 (
            .O(N__19282),
            .I(N__19263));
    Sp12to4 I__4152 (
            .O(N__19279),
            .I(N__19260));
    Span4Mux_h I__4151 (
            .O(N__19276),
            .I(N__19255));
    LocalMux I__4150 (
            .O(N__19273),
            .I(N__19255));
    SRMux I__4149 (
            .O(N__19272),
            .I(N__19252));
    Span4Mux_v I__4148 (
            .O(N__19269),
            .I(N__19249));
    Span4Mux_h I__4147 (
            .O(N__19266),
            .I(N__19246));
    Span4Mux_h I__4146 (
            .O(N__19263),
            .I(N__19243));
    Span12Mux_s9_v I__4145 (
            .O(N__19260),
            .I(N__19236));
    Sp12to4 I__4144 (
            .O(N__19255),
            .I(N__19236));
    LocalMux I__4143 (
            .O(N__19252),
            .I(N__19236));
    Odrv4 I__4142 (
            .O(N__19249),
            .I(\receive_module.n3674 ));
    Odrv4 I__4141 (
            .O(N__19246),
            .I(\receive_module.n3674 ));
    Odrv4 I__4140 (
            .O(N__19243),
            .I(\receive_module.n3674 ));
    Odrv12 I__4139 (
            .O(N__19236),
            .I(\receive_module.n3674 ));
    InMux I__4138 (
            .O(N__19227),
            .I(N__19224));
    LocalMux I__4137 (
            .O(N__19224),
            .I(N__19221));
    Span4Mux_v I__4136 (
            .O(N__19221),
            .I(N__19218));
    Sp12to4 I__4135 (
            .O(N__19218),
            .I(N__19215));
    Odrv12 I__4134 (
            .O(N__19215),
            .I(\line_buffer.n596 ));
    InMux I__4133 (
            .O(N__19212),
            .I(N__19209));
    LocalMux I__4132 (
            .O(N__19209),
            .I(N__19206));
    Span12Mux_v I__4131 (
            .O(N__19206),
            .I(N__19203));
    Odrv12 I__4130 (
            .O(N__19203),
            .I(\line_buffer.n588 ));
    InMux I__4129 (
            .O(N__19200),
            .I(N__19197));
    LocalMux I__4128 (
            .O(N__19197),
            .I(\line_buffer.n3623 ));
    InMux I__4127 (
            .O(N__19194),
            .I(bfn_17_10_0_));
    InMux I__4126 (
            .O(N__19191),
            .I(N__19187));
    InMux I__4125 (
            .O(N__19190),
            .I(N__19184));
    LocalMux I__4124 (
            .O(N__19187),
            .I(N__19181));
    LocalMux I__4123 (
            .O(N__19184),
            .I(N__19174));
    Span4Mux_v I__4122 (
            .O(N__19181),
            .I(N__19174));
    InMux I__4121 (
            .O(N__19180),
            .I(N__19169));
    InMux I__4120 (
            .O(N__19179),
            .I(N__19169));
    Odrv4 I__4119 (
            .O(N__19174),
            .I(\receive_module.rx_counter.Y_8 ));
    LocalMux I__4118 (
            .O(N__19169),
            .I(\receive_module.rx_counter.Y_8 ));
    InMux I__4117 (
            .O(N__19164),
            .I(N__19161));
    LocalMux I__4116 (
            .O(N__19161),
            .I(N__19158));
    Odrv4 I__4115 (
            .O(N__19158),
            .I(\tvp_video_buffer.BUFFER_1_2 ));
    InMux I__4114 (
            .O(N__19155),
            .I(N__19152));
    LocalMux I__4113 (
            .O(N__19152),
            .I(N__19149));
    Span4Mux_s1_v I__4112 (
            .O(N__19149),
            .I(N__19145));
    InMux I__4111 (
            .O(N__19148),
            .I(N__19142));
    Span4Mux_v I__4110 (
            .O(N__19145),
            .I(N__19135));
    LocalMux I__4109 (
            .O(N__19142),
            .I(N__19135));
    InMux I__4108 (
            .O(N__19141),
            .I(N__19130));
    InMux I__4107 (
            .O(N__19140),
            .I(N__19126));
    Span4Mux_v I__4106 (
            .O(N__19135),
            .I(N__19123));
    InMux I__4105 (
            .O(N__19134),
            .I(N__19120));
    InMux I__4104 (
            .O(N__19133),
            .I(N__19116));
    LocalMux I__4103 (
            .O(N__19130),
            .I(N__19113));
    InMux I__4102 (
            .O(N__19129),
            .I(N__19110));
    LocalMux I__4101 (
            .O(N__19126),
            .I(N__19107));
    Span4Mux_v I__4100 (
            .O(N__19123),
            .I(N__19102));
    LocalMux I__4099 (
            .O(N__19120),
            .I(N__19102));
    InMux I__4098 (
            .O(N__19119),
            .I(N__19099));
    LocalMux I__4097 (
            .O(N__19116),
            .I(N__19096));
    Span4Mux_v I__4096 (
            .O(N__19113),
            .I(N__19093));
    LocalMux I__4095 (
            .O(N__19110),
            .I(N__19090));
    Span4Mux_v I__4094 (
            .O(N__19107),
            .I(N__19087));
    Span4Mux_v I__4093 (
            .O(N__19102),
            .I(N__19082));
    LocalMux I__4092 (
            .O(N__19099),
            .I(N__19082));
    Sp12to4 I__4091 (
            .O(N__19096),
            .I(N__19079));
    Span4Mux_v I__4090 (
            .O(N__19093),
            .I(N__19074));
    Span4Mux_v I__4089 (
            .O(N__19090),
            .I(N__19074));
    Span4Mux_v I__4088 (
            .O(N__19087),
            .I(N__19069));
    Span4Mux_v I__4087 (
            .O(N__19082),
            .I(N__19069));
    Span12Mux_v I__4086 (
            .O(N__19079),
            .I(N__19064));
    Sp12to4 I__4085 (
            .O(N__19074),
            .I(N__19064));
    Span4Mux_h I__4084 (
            .O(N__19069),
            .I(N__19061));
    Odrv12 I__4083 (
            .O(N__19064),
            .I(RX_DATA_0));
    Odrv4 I__4082 (
            .O(N__19061),
            .I(RX_DATA_0));
    InMux I__4081 (
            .O(N__19056),
            .I(N__19052));
    InMux I__4080 (
            .O(N__19055),
            .I(N__19049));
    LocalMux I__4079 (
            .O(N__19052),
            .I(\receive_module.rx_counter.FRAME_COUNTER_4 ));
    LocalMux I__4078 (
            .O(N__19049),
            .I(\receive_module.rx_counter.FRAME_COUNTER_4 ));
    InMux I__4077 (
            .O(N__19044),
            .I(N__19040));
    InMux I__4076 (
            .O(N__19043),
            .I(N__19037));
    LocalMux I__4075 (
            .O(N__19040),
            .I(\receive_module.rx_counter.FRAME_COUNTER_2 ));
    LocalMux I__4074 (
            .O(N__19037),
            .I(\receive_module.rx_counter.FRAME_COUNTER_2 ));
    InMux I__4073 (
            .O(N__19032),
            .I(N__19028));
    InMux I__4072 (
            .O(N__19031),
            .I(N__19025));
    LocalMux I__4071 (
            .O(N__19028),
            .I(\receive_module.rx_counter.FRAME_COUNTER_0 ));
    LocalMux I__4070 (
            .O(N__19025),
            .I(\receive_module.rx_counter.FRAME_COUNTER_0 ));
    InMux I__4069 (
            .O(N__19020),
            .I(N__19016));
    InMux I__4068 (
            .O(N__19019),
            .I(N__19013));
    LocalMux I__4067 (
            .O(N__19016),
            .I(\receive_module.rx_counter.FRAME_COUNTER_3 ));
    LocalMux I__4066 (
            .O(N__19013),
            .I(\receive_module.rx_counter.FRAME_COUNTER_3 ));
    CascadeMux I__4065 (
            .O(N__19008),
            .I(\receive_module.rx_counter.n7_adj_619_cascade_ ));
    InMux I__4064 (
            .O(N__19005),
            .I(N__19002));
    LocalMux I__4063 (
            .O(N__19002),
            .I(\receive_module.rx_counter.n3519 ));
    InMux I__4062 (
            .O(N__18999),
            .I(N__18995));
    InMux I__4061 (
            .O(N__18998),
            .I(N__18992));
    LocalMux I__4060 (
            .O(N__18995),
            .I(N__18989));
    LocalMux I__4059 (
            .O(N__18992),
            .I(\receive_module.rx_counter.old_VS ));
    Odrv4 I__4058 (
            .O(N__18989),
            .I(\receive_module.rx_counter.old_VS ));
    CascadeMux I__4057 (
            .O(N__18984),
            .I(\receive_module.rx_counter.n11_cascade_ ));
    SRMux I__4056 (
            .O(N__18981),
            .I(N__18978));
    LocalMux I__4055 (
            .O(N__18978),
            .I(N__18975));
    Odrv12 I__4054 (
            .O(N__18975),
            .I(\receive_module.rx_counter.n2547 ));
    InMux I__4053 (
            .O(N__18972),
            .I(N__18969));
    LocalMux I__4052 (
            .O(N__18969),
            .I(\receive_module.rx_counter.n11 ));
    InMux I__4051 (
            .O(N__18966),
            .I(N__18963));
    LocalMux I__4050 (
            .O(N__18963),
            .I(N__18960));
    Span12Mux_s6_v I__4049 (
            .O(N__18960),
            .I(N__18956));
    InMux I__4048 (
            .O(N__18959),
            .I(N__18953));
    Odrv12 I__4047 (
            .O(N__18956),
            .I(PULSE_1HZ));
    LocalMux I__4046 (
            .O(N__18953),
            .I(PULSE_1HZ));
    CEMux I__4045 (
            .O(N__18948),
            .I(N__18944));
    CEMux I__4044 (
            .O(N__18947),
            .I(N__18941));
    LocalMux I__4043 (
            .O(N__18944),
            .I(N__18938));
    LocalMux I__4042 (
            .O(N__18941),
            .I(N__18935));
    Odrv4 I__4041 (
            .O(N__18938),
            .I(\receive_module.rx_counter.n3672 ));
    Odrv4 I__4040 (
            .O(N__18935),
            .I(\receive_module.rx_counter.n3672 ));
    InMux I__4039 (
            .O(N__18930),
            .I(N__18926));
    InMux I__4038 (
            .O(N__18929),
            .I(N__18923));
    LocalMux I__4037 (
            .O(N__18926),
            .I(N__18913));
    LocalMux I__4036 (
            .O(N__18923),
            .I(N__18910));
    InMux I__4035 (
            .O(N__18922),
            .I(N__18903));
    InMux I__4034 (
            .O(N__18921),
            .I(N__18903));
    InMux I__4033 (
            .O(N__18920),
            .I(N__18903));
    InMux I__4032 (
            .O(N__18919),
            .I(N__18900));
    InMux I__4031 (
            .O(N__18918),
            .I(N__18895));
    InMux I__4030 (
            .O(N__18917),
            .I(N__18895));
    InMux I__4029 (
            .O(N__18916),
            .I(N__18892));
    Span4Mux_v I__4028 (
            .O(N__18913),
            .I(N__18889));
    Span4Mux_h I__4027 (
            .O(N__18910),
            .I(N__18884));
    LocalMux I__4026 (
            .O(N__18903),
            .I(N__18884));
    LocalMux I__4025 (
            .O(N__18900),
            .I(RX_ADDR_12));
    LocalMux I__4024 (
            .O(N__18895),
            .I(RX_ADDR_12));
    LocalMux I__4023 (
            .O(N__18892),
            .I(RX_ADDR_12));
    Odrv4 I__4022 (
            .O(N__18889),
            .I(RX_ADDR_12));
    Odrv4 I__4021 (
            .O(N__18884),
            .I(RX_ADDR_12));
    CascadeMux I__4020 (
            .O(N__18873),
            .I(N__18868));
    CascadeMux I__4019 (
            .O(N__18872),
            .I(N__18863));
    CascadeMux I__4018 (
            .O(N__18871),
            .I(N__18860));
    InMux I__4017 (
            .O(N__18868),
            .I(N__18857));
    CascadeMux I__4016 (
            .O(N__18867),
            .I(N__18854));
    CascadeMux I__4015 (
            .O(N__18866),
            .I(N__18851));
    InMux I__4014 (
            .O(N__18863),
            .I(N__18846));
    InMux I__4013 (
            .O(N__18860),
            .I(N__18843));
    LocalMux I__4012 (
            .O(N__18857),
            .I(N__18840));
    InMux I__4011 (
            .O(N__18854),
            .I(N__18835));
    InMux I__4010 (
            .O(N__18851),
            .I(N__18835));
    CascadeMux I__4009 (
            .O(N__18850),
            .I(N__18830));
    CascadeMux I__4008 (
            .O(N__18849),
            .I(N__18827));
    LocalMux I__4007 (
            .O(N__18846),
            .I(N__18824));
    LocalMux I__4006 (
            .O(N__18843),
            .I(N__18817));
    Span4Mux_h I__4005 (
            .O(N__18840),
            .I(N__18817));
    LocalMux I__4004 (
            .O(N__18835),
            .I(N__18817));
    InMux I__4003 (
            .O(N__18834),
            .I(N__18814));
    InMux I__4002 (
            .O(N__18833),
            .I(N__18809));
    InMux I__4001 (
            .O(N__18830),
            .I(N__18809));
    InMux I__4000 (
            .O(N__18827),
            .I(N__18806));
    Span4Mux_v I__3999 (
            .O(N__18824),
            .I(N__18803));
    Span4Mux_v I__3998 (
            .O(N__18817),
            .I(N__18800));
    LocalMux I__3997 (
            .O(N__18814),
            .I(RX_ADDR_13));
    LocalMux I__3996 (
            .O(N__18809),
            .I(RX_ADDR_13));
    LocalMux I__3995 (
            .O(N__18806),
            .I(RX_ADDR_13));
    Odrv4 I__3994 (
            .O(N__18803),
            .I(RX_ADDR_13));
    Odrv4 I__3993 (
            .O(N__18800),
            .I(RX_ADDR_13));
    InMux I__3992 (
            .O(N__18789),
            .I(N__18785));
    InMux I__3991 (
            .O(N__18788),
            .I(N__18782));
    LocalMux I__3990 (
            .O(N__18785),
            .I(N__18773));
    LocalMux I__3989 (
            .O(N__18782),
            .I(N__18770));
    InMux I__3988 (
            .O(N__18781),
            .I(N__18763));
    InMux I__3987 (
            .O(N__18780),
            .I(N__18763));
    InMux I__3986 (
            .O(N__18779),
            .I(N__18763));
    InMux I__3985 (
            .O(N__18778),
            .I(N__18759));
    InMux I__3984 (
            .O(N__18777),
            .I(N__18754));
    InMux I__3983 (
            .O(N__18776),
            .I(N__18754));
    Span4Mux_v I__3982 (
            .O(N__18773),
            .I(N__18751));
    Span4Mux_h I__3981 (
            .O(N__18770),
            .I(N__18748));
    LocalMux I__3980 (
            .O(N__18763),
            .I(N__18745));
    InMux I__3979 (
            .O(N__18762),
            .I(N__18742));
    LocalMux I__3978 (
            .O(N__18759),
            .I(RX_ADDR_11));
    LocalMux I__3977 (
            .O(N__18754),
            .I(RX_ADDR_11));
    Odrv4 I__3976 (
            .O(N__18751),
            .I(RX_ADDR_11));
    Odrv4 I__3975 (
            .O(N__18748),
            .I(RX_ADDR_11));
    Odrv4 I__3974 (
            .O(N__18745),
            .I(RX_ADDR_11));
    LocalMux I__3973 (
            .O(N__18742),
            .I(RX_ADDR_11));
    SRMux I__3972 (
            .O(N__18729),
            .I(N__18726));
    LocalMux I__3971 (
            .O(N__18726),
            .I(N__18722));
    SRMux I__3970 (
            .O(N__18725),
            .I(N__18719));
    Span4Mux_v I__3969 (
            .O(N__18722),
            .I(N__18712));
    LocalMux I__3968 (
            .O(N__18719),
            .I(N__18712));
    SRMux I__3967 (
            .O(N__18718),
            .I(N__18709));
    SRMux I__3966 (
            .O(N__18717),
            .I(N__18706));
    Span4Mux_v I__3965 (
            .O(N__18712),
            .I(N__18699));
    LocalMux I__3964 (
            .O(N__18709),
            .I(N__18699));
    LocalMux I__3963 (
            .O(N__18706),
            .I(N__18699));
    Span4Mux_v I__3962 (
            .O(N__18699),
            .I(N__18696));
    Span4Mux_h I__3961 (
            .O(N__18696),
            .I(N__18693));
    Odrv4 I__3960 (
            .O(N__18693),
            .I(\line_buffer.n538 ));
    InMux I__3959 (
            .O(N__18690),
            .I(N__18687));
    LocalMux I__3958 (
            .O(N__18687),
            .I(N__18683));
    InMux I__3957 (
            .O(N__18686),
            .I(N__18680));
    Odrv4 I__3956 (
            .O(N__18683),
            .I(\transmit_module.X_DELTA_PATTERN_0 ));
    LocalMux I__3955 (
            .O(N__18680),
            .I(\transmit_module.X_DELTA_PATTERN_0 ));
    InMux I__3954 (
            .O(N__18675),
            .I(N__18672));
    LocalMux I__3953 (
            .O(N__18672),
            .I(N__18669));
    Span4Mux_h I__3952 (
            .O(N__18669),
            .I(N__18666));
    Odrv4 I__3951 (
            .O(N__18666),
            .I(\transmit_module.X_DELTA_PATTERN_15 ));
    CEMux I__3950 (
            .O(N__18663),
            .I(N__18659));
    CEMux I__3949 (
            .O(N__18662),
            .I(N__18656));
    LocalMux I__3948 (
            .O(N__18659),
            .I(N__18652));
    LocalMux I__3947 (
            .O(N__18656),
            .I(N__18649));
    CEMux I__3946 (
            .O(N__18655),
            .I(N__18646));
    Span4Mux_v I__3945 (
            .O(N__18652),
            .I(N__18642));
    Span4Mux_h I__3944 (
            .O(N__18649),
            .I(N__18639));
    LocalMux I__3943 (
            .O(N__18646),
            .I(N__18636));
    CEMux I__3942 (
            .O(N__18645),
            .I(N__18633));
    Odrv4 I__3941 (
            .O(N__18642),
            .I(\transmit_module.n2084 ));
    Odrv4 I__3940 (
            .O(N__18639),
            .I(\transmit_module.n2084 ));
    Odrv12 I__3939 (
            .O(N__18636),
            .I(\transmit_module.n2084 ));
    LocalMux I__3938 (
            .O(N__18633),
            .I(\transmit_module.n2084 ));
    InMux I__3937 (
            .O(N__18624),
            .I(N__18618));
    InMux I__3936 (
            .O(N__18623),
            .I(N__18613));
    InMux I__3935 (
            .O(N__18622),
            .I(N__18613));
    InMux I__3934 (
            .O(N__18621),
            .I(N__18610));
    LocalMux I__3933 (
            .O(N__18618),
            .I(\receive_module.rx_counter.Y_0 ));
    LocalMux I__3932 (
            .O(N__18613),
            .I(\receive_module.rx_counter.Y_0 ));
    LocalMux I__3931 (
            .O(N__18610),
            .I(\receive_module.rx_counter.Y_0 ));
    InMux I__3930 (
            .O(N__18603),
            .I(bfn_17_9_0_));
    CascadeMux I__3929 (
            .O(N__18600),
            .I(N__18596));
    InMux I__3928 (
            .O(N__18599),
            .I(N__18591));
    InMux I__3927 (
            .O(N__18596),
            .I(N__18588));
    InMux I__3926 (
            .O(N__18595),
            .I(N__18583));
    InMux I__3925 (
            .O(N__18594),
            .I(N__18583));
    LocalMux I__3924 (
            .O(N__18591),
            .I(\receive_module.rx_counter.Y_1 ));
    LocalMux I__3923 (
            .O(N__18588),
            .I(\receive_module.rx_counter.Y_1 ));
    LocalMux I__3922 (
            .O(N__18583),
            .I(\receive_module.rx_counter.Y_1 ));
    InMux I__3921 (
            .O(N__18576),
            .I(\receive_module.rx_counter.n3172 ));
    InMux I__3920 (
            .O(N__18573),
            .I(N__18567));
    InMux I__3919 (
            .O(N__18572),
            .I(N__18562));
    InMux I__3918 (
            .O(N__18571),
            .I(N__18562));
    InMux I__3917 (
            .O(N__18570),
            .I(N__18559));
    LocalMux I__3916 (
            .O(N__18567),
            .I(\receive_module.rx_counter.Y_2 ));
    LocalMux I__3915 (
            .O(N__18562),
            .I(\receive_module.rx_counter.Y_2 ));
    LocalMux I__3914 (
            .O(N__18559),
            .I(\receive_module.rx_counter.Y_2 ));
    InMux I__3913 (
            .O(N__18552),
            .I(\receive_module.rx_counter.n3173 ));
    CascadeMux I__3912 (
            .O(N__18549),
            .I(N__18546));
    InMux I__3911 (
            .O(N__18546),
            .I(N__18540));
    InMux I__3910 (
            .O(N__18545),
            .I(N__18537));
    InMux I__3909 (
            .O(N__18544),
            .I(N__18532));
    InMux I__3908 (
            .O(N__18543),
            .I(N__18532));
    LocalMux I__3907 (
            .O(N__18540),
            .I(\receive_module.rx_counter.Y_3 ));
    LocalMux I__3906 (
            .O(N__18537),
            .I(\receive_module.rx_counter.Y_3 ));
    LocalMux I__3905 (
            .O(N__18532),
            .I(\receive_module.rx_counter.Y_3 ));
    InMux I__3904 (
            .O(N__18525),
            .I(\receive_module.rx_counter.n3174 ));
    InMux I__3903 (
            .O(N__18522),
            .I(N__18516));
    InMux I__3902 (
            .O(N__18521),
            .I(N__18509));
    InMux I__3901 (
            .O(N__18520),
            .I(N__18509));
    InMux I__3900 (
            .O(N__18519),
            .I(N__18509));
    LocalMux I__3899 (
            .O(N__18516),
            .I(\receive_module.rx_counter.Y_4 ));
    LocalMux I__3898 (
            .O(N__18509),
            .I(\receive_module.rx_counter.Y_4 ));
    InMux I__3897 (
            .O(N__18504),
            .I(\receive_module.rx_counter.n3175 ));
    InMux I__3896 (
            .O(N__18501),
            .I(N__18496));
    InMux I__3895 (
            .O(N__18500),
            .I(N__18491));
    InMux I__3894 (
            .O(N__18499),
            .I(N__18491));
    LocalMux I__3893 (
            .O(N__18496),
            .I(\receive_module.rx_counter.Y_5 ));
    LocalMux I__3892 (
            .O(N__18491),
            .I(\receive_module.rx_counter.Y_5 ));
    InMux I__3891 (
            .O(N__18486),
            .I(\receive_module.rx_counter.n3176 ));
    InMux I__3890 (
            .O(N__18483),
            .I(N__18478));
    InMux I__3889 (
            .O(N__18482),
            .I(N__18475));
    InMux I__3888 (
            .O(N__18481),
            .I(N__18472));
    LocalMux I__3887 (
            .O(N__18478),
            .I(\receive_module.rx_counter.Y_6 ));
    LocalMux I__3886 (
            .O(N__18475),
            .I(\receive_module.rx_counter.Y_6 ));
    LocalMux I__3885 (
            .O(N__18472),
            .I(\receive_module.rx_counter.Y_6 ));
    InMux I__3884 (
            .O(N__18465),
            .I(\receive_module.rx_counter.n3177 ));
    InMux I__3883 (
            .O(N__18462),
            .I(N__18456));
    InMux I__3882 (
            .O(N__18461),
            .I(N__18451));
    InMux I__3881 (
            .O(N__18460),
            .I(N__18451));
    InMux I__3880 (
            .O(N__18459),
            .I(N__18448));
    LocalMux I__3879 (
            .O(N__18456),
            .I(\receive_module.rx_counter.Y_7 ));
    LocalMux I__3878 (
            .O(N__18451),
            .I(\receive_module.rx_counter.Y_7 ));
    LocalMux I__3877 (
            .O(N__18448),
            .I(\receive_module.rx_counter.Y_7 ));
    InMux I__3876 (
            .O(N__18441),
            .I(\receive_module.rx_counter.n3178 ));
    InMux I__3875 (
            .O(N__18438),
            .I(N__18435));
    LocalMux I__3874 (
            .O(N__18435),
            .I(N__18432));
    Span4Mux_v I__3873 (
            .O(N__18432),
            .I(N__18429));
    Span4Mux_h I__3872 (
            .O(N__18429),
            .I(N__18426));
    Span4Mux_h I__3871 (
            .O(N__18426),
            .I(N__18423));
    Sp12to4 I__3870 (
            .O(N__18423),
            .I(N__18420));
    Span12Mux_v I__3869 (
            .O(N__18420),
            .I(N__18417));
    Odrv12 I__3868 (
            .O(N__18417),
            .I(\line_buffer.n532 ));
    CascadeMux I__3867 (
            .O(N__18414),
            .I(N__18411));
    InMux I__3866 (
            .O(N__18411),
            .I(N__18408));
    LocalMux I__3865 (
            .O(N__18408),
            .I(N__18405));
    Span4Mux_v I__3864 (
            .O(N__18405),
            .I(N__18402));
    Sp12to4 I__3863 (
            .O(N__18402),
            .I(N__18399));
    Span12Mux_v I__3862 (
            .O(N__18399),
            .I(N__18396));
    Odrv12 I__3861 (
            .O(N__18396),
            .I(\line_buffer.n524 ));
    InMux I__3860 (
            .O(N__18393),
            .I(N__18390));
    LocalMux I__3859 (
            .O(N__18390),
            .I(N__18387));
    Sp12to4 I__3858 (
            .O(N__18387),
            .I(N__18384));
    Odrv12 I__3857 (
            .O(N__18384),
            .I(\line_buffer.n467 ));
    CascadeMux I__3856 (
            .O(N__18381),
            .I(N__18378));
    InMux I__3855 (
            .O(N__18378),
            .I(N__18375));
    LocalMux I__3854 (
            .O(N__18375),
            .I(N__18372));
    Span4Mux_v I__3853 (
            .O(N__18372),
            .I(N__18369));
    Sp12to4 I__3852 (
            .O(N__18369),
            .I(N__18366));
    Span12Mux_h I__3851 (
            .O(N__18366),
            .I(N__18363));
    Odrv12 I__3850 (
            .O(N__18363),
            .I(\line_buffer.n459 ));
    InMux I__3849 (
            .O(N__18360),
            .I(N__18357));
    LocalMux I__3848 (
            .O(N__18357),
            .I(\line_buffer.n3587 ));
    CascadeMux I__3847 (
            .O(N__18354),
            .I(\line_buffer.n3590_cascade_ ));
    InMux I__3846 (
            .O(N__18351),
            .I(N__18348));
    LocalMux I__3845 (
            .O(N__18348),
            .I(\line_buffer.n3626 ));
    InMux I__3844 (
            .O(N__18345),
            .I(N__18342));
    LocalMux I__3843 (
            .O(N__18342),
            .I(TX_DATA_3));
    IoInMux I__3842 (
            .O(N__18339),
            .I(N__18334));
    IoInMux I__3841 (
            .O(N__18338),
            .I(N__18331));
    IoInMux I__3840 (
            .O(N__18337),
            .I(N__18328));
    LocalMux I__3839 (
            .O(N__18334),
            .I(N__18325));
    LocalMux I__3838 (
            .O(N__18331),
            .I(N__18322));
    LocalMux I__3837 (
            .O(N__18328),
            .I(N__18319));
    IoSpan4Mux I__3836 (
            .O(N__18325),
            .I(N__18316));
    IoSpan4Mux I__3835 (
            .O(N__18322),
            .I(N__18313));
    Span4Mux_s3_h I__3834 (
            .O(N__18319),
            .I(N__18310));
    Span4Mux_s3_v I__3833 (
            .O(N__18316),
            .I(N__18307));
    Span4Mux_s3_v I__3832 (
            .O(N__18313),
            .I(N__18304));
    Span4Mux_h I__3831 (
            .O(N__18310),
            .I(N__18301));
    Sp12to4 I__3830 (
            .O(N__18307),
            .I(N__18298));
    Sp12to4 I__3829 (
            .O(N__18304),
            .I(N__18295));
    Span4Mux_h I__3828 (
            .O(N__18301),
            .I(N__18292));
    Span12Mux_s10_v I__3827 (
            .O(N__18298),
            .I(N__18289));
    Span12Mux_h I__3826 (
            .O(N__18295),
            .I(N__18286));
    Span4Mux_h I__3825 (
            .O(N__18292),
            .I(N__18283));
    Odrv12 I__3824 (
            .O(N__18289),
            .I(n1815));
    Odrv12 I__3823 (
            .O(N__18286),
            .I(n1815));
    Odrv4 I__3822 (
            .O(N__18283),
            .I(n1815));
    SRMux I__3821 (
            .O(N__18276),
            .I(N__18272));
    SRMux I__3820 (
            .O(N__18275),
            .I(N__18267));
    LocalMux I__3819 (
            .O(N__18272),
            .I(N__18264));
    SRMux I__3818 (
            .O(N__18271),
            .I(N__18261));
    SRMux I__3817 (
            .O(N__18270),
            .I(N__18258));
    LocalMux I__3816 (
            .O(N__18267),
            .I(N__18255));
    Span4Mux_s2_v I__3815 (
            .O(N__18264),
            .I(N__18248));
    LocalMux I__3814 (
            .O(N__18261),
            .I(N__18248));
    LocalMux I__3813 (
            .O(N__18258),
            .I(N__18248));
    Span4Mux_v I__3812 (
            .O(N__18255),
            .I(N__18245));
    Span4Mux_v I__3811 (
            .O(N__18248),
            .I(N__18242));
    Span4Mux_v I__3810 (
            .O(N__18245),
            .I(N__18239));
    Span4Mux_h I__3809 (
            .O(N__18242),
            .I(N__18236));
    Span4Mux_h I__3808 (
            .O(N__18239),
            .I(N__18233));
    Span4Mux_h I__3807 (
            .O(N__18236),
            .I(N__18230));
    Odrv4 I__3806 (
            .O(N__18233),
            .I(\line_buffer.n602 ));
    Odrv4 I__3805 (
            .O(N__18230),
            .I(\line_buffer.n602 ));
    IoInMux I__3804 (
            .O(N__18225),
            .I(N__18222));
    LocalMux I__3803 (
            .O(N__18222),
            .I(N__18219));
    IoSpan4Mux I__3802 (
            .O(N__18219),
            .I(N__18216));
    Span4Mux_s2_h I__3801 (
            .O(N__18216),
            .I(N__18212));
    IoInMux I__3800 (
            .O(N__18215),
            .I(N__18209));
    Span4Mux_v I__3799 (
            .O(N__18212),
            .I(N__18206));
    LocalMux I__3798 (
            .O(N__18209),
            .I(N__18203));
    Sp12to4 I__3797 (
            .O(N__18206),
            .I(N__18200));
    IoSpan4Mux I__3796 (
            .O(N__18203),
            .I(N__18197));
    Span12Mux_h I__3795 (
            .O(N__18200),
            .I(N__18194));
    Span4Mux_s3_v I__3794 (
            .O(N__18197),
            .I(N__18191));
    Odrv12 I__3793 (
            .O(N__18194),
            .I(GB_BUFFER_DEBUG_c_3_c_THRU_CO));
    Odrv4 I__3792 (
            .O(N__18191),
            .I(GB_BUFFER_DEBUG_c_3_c_THRU_CO));
    IoInMux I__3791 (
            .O(N__18186),
            .I(N__18183));
    LocalMux I__3790 (
            .O(N__18183),
            .I(N__18180));
    IoSpan4Mux I__3789 (
            .O(N__18180),
            .I(N__18177));
    Span4Mux_s3_h I__3788 (
            .O(N__18177),
            .I(N__18173));
    InMux I__3787 (
            .O(N__18176),
            .I(N__18170));
    Span4Mux_h I__3786 (
            .O(N__18173),
            .I(N__18167));
    LocalMux I__3785 (
            .O(N__18170),
            .I(N__18164));
    Span4Mux_h I__3784 (
            .O(N__18167),
            .I(N__18160));
    Span4Mux_h I__3783 (
            .O(N__18164),
            .I(N__18157));
    InMux I__3782 (
            .O(N__18163),
            .I(N__18154));
    Odrv4 I__3781 (
            .O(N__18160),
            .I(DEBUG_c_0));
    Odrv4 I__3780 (
            .O(N__18157),
            .I(DEBUG_c_0));
    LocalMux I__3779 (
            .O(N__18154),
            .I(DEBUG_c_0));
    IoInMux I__3778 (
            .O(N__18147),
            .I(N__18144));
    LocalMux I__3777 (
            .O(N__18144),
            .I(N__18141));
    Span4Mux_s3_v I__3776 (
            .O(N__18141),
            .I(N__18138));
    Span4Mux_h I__3775 (
            .O(N__18138),
            .I(N__18135));
    Odrv4 I__3774 (
            .O(N__18135),
            .I(LED_c));
    InMux I__3773 (
            .O(N__18132),
            .I(N__18129));
    LocalMux I__3772 (
            .O(N__18129),
            .I(N__18126));
    Sp12to4 I__3771 (
            .O(N__18126),
            .I(N__18123));
    Span12Mux_v I__3770 (
            .O(N__18123),
            .I(N__18120));
    Span12Mux_h I__3769 (
            .O(N__18120),
            .I(N__18117));
    Odrv12 I__3768 (
            .O(N__18117),
            .I(TVP_VIDEO_c_2));
    InMux I__3767 (
            .O(N__18114),
            .I(N__18111));
    LocalMux I__3766 (
            .O(N__18111),
            .I(\tvp_video_buffer.BUFFER_0_2 ));
    SRMux I__3765 (
            .O(N__18108),
            .I(N__18105));
    LocalMux I__3764 (
            .O(N__18105),
            .I(N__18101));
    SRMux I__3763 (
            .O(N__18104),
            .I(N__18098));
    Span4Mux_v I__3762 (
            .O(N__18101),
            .I(N__18092));
    LocalMux I__3761 (
            .O(N__18098),
            .I(N__18092));
    SRMux I__3760 (
            .O(N__18097),
            .I(N__18088));
    Span4Mux_v I__3759 (
            .O(N__18092),
            .I(N__18085));
    SRMux I__3758 (
            .O(N__18091),
            .I(N__18082));
    LocalMux I__3757 (
            .O(N__18088),
            .I(N__18075));
    Sp12to4 I__3756 (
            .O(N__18085),
            .I(N__18075));
    LocalMux I__3755 (
            .O(N__18082),
            .I(N__18075));
    Span12Mux_v I__3754 (
            .O(N__18075),
            .I(N__18072));
    Odrv12 I__3753 (
            .O(N__18072),
            .I(\line_buffer.n474 ));
    InMux I__3752 (
            .O(N__18069),
            .I(N__18066));
    LocalMux I__3751 (
            .O(N__18066),
            .I(N__18063));
    Odrv4 I__3750 (
            .O(N__18063),
            .I(\receive_module.n128 ));
    CascadeMux I__3749 (
            .O(N__18060),
            .I(N__18056));
    CascadeMux I__3748 (
            .O(N__18059),
            .I(N__18053));
    CascadeBuf I__3747 (
            .O(N__18056),
            .I(N__18050));
    CascadeBuf I__3746 (
            .O(N__18053),
            .I(N__18047));
    CascadeMux I__3745 (
            .O(N__18050),
            .I(N__18044));
    CascadeMux I__3744 (
            .O(N__18047),
            .I(N__18041));
    CascadeBuf I__3743 (
            .O(N__18044),
            .I(N__18038));
    CascadeBuf I__3742 (
            .O(N__18041),
            .I(N__18035));
    CascadeMux I__3741 (
            .O(N__18038),
            .I(N__18032));
    CascadeMux I__3740 (
            .O(N__18035),
            .I(N__18029));
    CascadeBuf I__3739 (
            .O(N__18032),
            .I(N__18026));
    CascadeBuf I__3738 (
            .O(N__18029),
            .I(N__18023));
    CascadeMux I__3737 (
            .O(N__18026),
            .I(N__18020));
    CascadeMux I__3736 (
            .O(N__18023),
            .I(N__18017));
    CascadeBuf I__3735 (
            .O(N__18020),
            .I(N__18014));
    CascadeBuf I__3734 (
            .O(N__18017),
            .I(N__18011));
    CascadeMux I__3733 (
            .O(N__18014),
            .I(N__18008));
    CascadeMux I__3732 (
            .O(N__18011),
            .I(N__18005));
    CascadeBuf I__3731 (
            .O(N__18008),
            .I(N__18002));
    CascadeBuf I__3730 (
            .O(N__18005),
            .I(N__17999));
    CascadeMux I__3729 (
            .O(N__18002),
            .I(N__17996));
    CascadeMux I__3728 (
            .O(N__17999),
            .I(N__17993));
    CascadeBuf I__3727 (
            .O(N__17996),
            .I(N__17990));
    CascadeBuf I__3726 (
            .O(N__17993),
            .I(N__17987));
    CascadeMux I__3725 (
            .O(N__17990),
            .I(N__17984));
    CascadeMux I__3724 (
            .O(N__17987),
            .I(N__17981));
    CascadeBuf I__3723 (
            .O(N__17984),
            .I(N__17978));
    CascadeBuf I__3722 (
            .O(N__17981),
            .I(N__17975));
    CascadeMux I__3721 (
            .O(N__17978),
            .I(N__17972));
    CascadeMux I__3720 (
            .O(N__17975),
            .I(N__17969));
    CascadeBuf I__3719 (
            .O(N__17972),
            .I(N__17966));
    CascadeBuf I__3718 (
            .O(N__17969),
            .I(N__17963));
    CascadeMux I__3717 (
            .O(N__17966),
            .I(N__17960));
    CascadeMux I__3716 (
            .O(N__17963),
            .I(N__17957));
    CascadeBuf I__3715 (
            .O(N__17960),
            .I(N__17954));
    CascadeBuf I__3714 (
            .O(N__17957),
            .I(N__17951));
    CascadeMux I__3713 (
            .O(N__17954),
            .I(N__17948));
    CascadeMux I__3712 (
            .O(N__17951),
            .I(N__17945));
    CascadeBuf I__3711 (
            .O(N__17948),
            .I(N__17942));
    CascadeBuf I__3710 (
            .O(N__17945),
            .I(N__17939));
    CascadeMux I__3709 (
            .O(N__17942),
            .I(N__17936));
    CascadeMux I__3708 (
            .O(N__17939),
            .I(N__17933));
    CascadeBuf I__3707 (
            .O(N__17936),
            .I(N__17930));
    CascadeBuf I__3706 (
            .O(N__17933),
            .I(N__17927));
    CascadeMux I__3705 (
            .O(N__17930),
            .I(N__17924));
    CascadeMux I__3704 (
            .O(N__17927),
            .I(N__17921));
    CascadeBuf I__3703 (
            .O(N__17924),
            .I(N__17918));
    CascadeBuf I__3702 (
            .O(N__17921),
            .I(N__17915));
    CascadeMux I__3701 (
            .O(N__17918),
            .I(N__17912));
    CascadeMux I__3700 (
            .O(N__17915),
            .I(N__17909));
    CascadeBuf I__3699 (
            .O(N__17912),
            .I(N__17906));
    CascadeBuf I__3698 (
            .O(N__17909),
            .I(N__17903));
    CascadeMux I__3697 (
            .O(N__17906),
            .I(N__17900));
    CascadeMux I__3696 (
            .O(N__17903),
            .I(N__17897));
    CascadeBuf I__3695 (
            .O(N__17900),
            .I(N__17894));
    CascadeBuf I__3694 (
            .O(N__17897),
            .I(N__17891));
    CascadeMux I__3693 (
            .O(N__17894),
            .I(N__17888));
    CascadeMux I__3692 (
            .O(N__17891),
            .I(N__17885));
    CascadeBuf I__3691 (
            .O(N__17888),
            .I(N__17882));
    CascadeBuf I__3690 (
            .O(N__17885),
            .I(N__17879));
    CascadeMux I__3689 (
            .O(N__17882),
            .I(N__17876));
    CascadeMux I__3688 (
            .O(N__17879),
            .I(N__17873));
    InMux I__3687 (
            .O(N__17876),
            .I(N__17870));
    InMux I__3686 (
            .O(N__17873),
            .I(N__17867));
    LocalMux I__3685 (
            .O(N__17870),
            .I(N__17864));
    LocalMux I__3684 (
            .O(N__17867),
            .I(N__17861));
    Span4Mux_s1_v I__3683 (
            .O(N__17864),
            .I(N__17858));
    Span4Mux_s1_v I__3682 (
            .O(N__17861),
            .I(N__17855));
    Span4Mux_v I__3681 (
            .O(N__17858),
            .I(N__17850));
    Span4Mux_v I__3680 (
            .O(N__17855),
            .I(N__17847));
    CascadeMux I__3679 (
            .O(N__17854),
            .I(N__17844));
    InMux I__3678 (
            .O(N__17853),
            .I(N__17841));
    Sp12to4 I__3677 (
            .O(N__17850),
            .I(N__17838));
    Sp12to4 I__3676 (
            .O(N__17847),
            .I(N__17835));
    InMux I__3675 (
            .O(N__17844),
            .I(N__17832));
    LocalMux I__3674 (
            .O(N__17841),
            .I(N__17829));
    Span12Mux_h I__3673 (
            .O(N__17838),
            .I(N__17824));
    Span12Mux_h I__3672 (
            .O(N__17835),
            .I(N__17824));
    LocalMux I__3671 (
            .O(N__17832),
            .I(RX_ADDR_9));
    Odrv4 I__3670 (
            .O(N__17829),
            .I(RX_ADDR_9));
    Odrv12 I__3669 (
            .O(N__17824),
            .I(RX_ADDR_9));
    InMux I__3668 (
            .O(N__17817),
            .I(N__17814));
    LocalMux I__3667 (
            .O(N__17814),
            .I(N__17811));
    Odrv4 I__3666 (
            .O(N__17811),
            .I(\receive_module.n134 ));
    CascadeMux I__3665 (
            .O(N__17808),
            .I(N__17805));
    CascadeBuf I__3664 (
            .O(N__17805),
            .I(N__17801));
    CascadeMux I__3663 (
            .O(N__17804),
            .I(N__17798));
    CascadeMux I__3662 (
            .O(N__17801),
            .I(N__17795));
    CascadeBuf I__3661 (
            .O(N__17798),
            .I(N__17792));
    CascadeBuf I__3660 (
            .O(N__17795),
            .I(N__17789));
    CascadeMux I__3659 (
            .O(N__17792),
            .I(N__17786));
    CascadeMux I__3658 (
            .O(N__17789),
            .I(N__17783));
    CascadeBuf I__3657 (
            .O(N__17786),
            .I(N__17780));
    CascadeBuf I__3656 (
            .O(N__17783),
            .I(N__17777));
    CascadeMux I__3655 (
            .O(N__17780),
            .I(N__17774));
    CascadeMux I__3654 (
            .O(N__17777),
            .I(N__17771));
    CascadeBuf I__3653 (
            .O(N__17774),
            .I(N__17768));
    CascadeBuf I__3652 (
            .O(N__17771),
            .I(N__17765));
    CascadeMux I__3651 (
            .O(N__17768),
            .I(N__17762));
    CascadeMux I__3650 (
            .O(N__17765),
            .I(N__17759));
    CascadeBuf I__3649 (
            .O(N__17762),
            .I(N__17756));
    CascadeBuf I__3648 (
            .O(N__17759),
            .I(N__17753));
    CascadeMux I__3647 (
            .O(N__17756),
            .I(N__17750));
    CascadeMux I__3646 (
            .O(N__17753),
            .I(N__17747));
    CascadeBuf I__3645 (
            .O(N__17750),
            .I(N__17744));
    CascadeBuf I__3644 (
            .O(N__17747),
            .I(N__17741));
    CascadeMux I__3643 (
            .O(N__17744),
            .I(N__17738));
    CascadeMux I__3642 (
            .O(N__17741),
            .I(N__17735));
    CascadeBuf I__3641 (
            .O(N__17738),
            .I(N__17732));
    CascadeBuf I__3640 (
            .O(N__17735),
            .I(N__17729));
    CascadeMux I__3639 (
            .O(N__17732),
            .I(N__17726));
    CascadeMux I__3638 (
            .O(N__17729),
            .I(N__17723));
    CascadeBuf I__3637 (
            .O(N__17726),
            .I(N__17720));
    CascadeBuf I__3636 (
            .O(N__17723),
            .I(N__17717));
    CascadeMux I__3635 (
            .O(N__17720),
            .I(N__17714));
    CascadeMux I__3634 (
            .O(N__17717),
            .I(N__17711));
    CascadeBuf I__3633 (
            .O(N__17714),
            .I(N__17708));
    CascadeBuf I__3632 (
            .O(N__17711),
            .I(N__17705));
    CascadeMux I__3631 (
            .O(N__17708),
            .I(N__17702));
    CascadeMux I__3630 (
            .O(N__17705),
            .I(N__17699));
    CascadeBuf I__3629 (
            .O(N__17702),
            .I(N__17696));
    CascadeBuf I__3628 (
            .O(N__17699),
            .I(N__17693));
    CascadeMux I__3627 (
            .O(N__17696),
            .I(N__17690));
    CascadeMux I__3626 (
            .O(N__17693),
            .I(N__17687));
    CascadeBuf I__3625 (
            .O(N__17690),
            .I(N__17684));
    CascadeBuf I__3624 (
            .O(N__17687),
            .I(N__17681));
    CascadeMux I__3623 (
            .O(N__17684),
            .I(N__17678));
    CascadeMux I__3622 (
            .O(N__17681),
            .I(N__17675));
    CascadeBuf I__3621 (
            .O(N__17678),
            .I(N__17672));
    CascadeBuf I__3620 (
            .O(N__17675),
            .I(N__17669));
    CascadeMux I__3619 (
            .O(N__17672),
            .I(N__17666));
    CascadeMux I__3618 (
            .O(N__17669),
            .I(N__17663));
    CascadeBuf I__3617 (
            .O(N__17666),
            .I(N__17660));
    CascadeBuf I__3616 (
            .O(N__17663),
            .I(N__17657));
    CascadeMux I__3615 (
            .O(N__17660),
            .I(N__17654));
    CascadeMux I__3614 (
            .O(N__17657),
            .I(N__17651));
    CascadeBuf I__3613 (
            .O(N__17654),
            .I(N__17648));
    CascadeBuf I__3612 (
            .O(N__17651),
            .I(N__17645));
    CascadeMux I__3611 (
            .O(N__17648),
            .I(N__17642));
    CascadeMux I__3610 (
            .O(N__17645),
            .I(N__17639));
    CascadeBuf I__3609 (
            .O(N__17642),
            .I(N__17636));
    CascadeBuf I__3608 (
            .O(N__17639),
            .I(N__17633));
    CascadeMux I__3607 (
            .O(N__17636),
            .I(N__17630));
    CascadeMux I__3606 (
            .O(N__17633),
            .I(N__17627));
    CascadeBuf I__3605 (
            .O(N__17630),
            .I(N__17624));
    InMux I__3604 (
            .O(N__17627),
            .I(N__17621));
    CascadeMux I__3603 (
            .O(N__17624),
            .I(N__17618));
    LocalMux I__3602 (
            .O(N__17621),
            .I(N__17614));
    InMux I__3601 (
            .O(N__17618),
            .I(N__17611));
    InMux I__3600 (
            .O(N__17617),
            .I(N__17608));
    Span4Mux_s2_v I__3599 (
            .O(N__17614),
            .I(N__17605));
    LocalMux I__3598 (
            .O(N__17611),
            .I(N__17602));
    LocalMux I__3597 (
            .O(N__17608),
            .I(N__17599));
    Sp12to4 I__3596 (
            .O(N__17605),
            .I(N__17595));
    Sp12to4 I__3595 (
            .O(N__17602),
            .I(N__17592));
    Span4Mux_h I__3594 (
            .O(N__17599),
            .I(N__17589));
    InMux I__3593 (
            .O(N__17598),
            .I(N__17586));
    Span12Mux_h I__3592 (
            .O(N__17595),
            .I(N__17583));
    Span12Mux_v I__3591 (
            .O(N__17592),
            .I(N__17580));
    Odrv4 I__3590 (
            .O(N__17589),
            .I(RX_ADDR_3));
    LocalMux I__3589 (
            .O(N__17586),
            .I(RX_ADDR_3));
    Odrv12 I__3588 (
            .O(N__17583),
            .I(RX_ADDR_3));
    Odrv12 I__3587 (
            .O(N__17580),
            .I(RX_ADDR_3));
    InMux I__3586 (
            .O(N__17571),
            .I(N__17568));
    LocalMux I__3585 (
            .O(N__17568),
            .I(N__17565));
    Odrv4 I__3584 (
            .O(N__17565),
            .I(\receive_module.n133 ));
    CascadeMux I__3583 (
            .O(N__17562),
            .I(N__17558));
    CascadeMux I__3582 (
            .O(N__17561),
            .I(N__17555));
    CascadeBuf I__3581 (
            .O(N__17558),
            .I(N__17552));
    CascadeBuf I__3580 (
            .O(N__17555),
            .I(N__17549));
    CascadeMux I__3579 (
            .O(N__17552),
            .I(N__17546));
    CascadeMux I__3578 (
            .O(N__17549),
            .I(N__17543));
    CascadeBuf I__3577 (
            .O(N__17546),
            .I(N__17540));
    CascadeBuf I__3576 (
            .O(N__17543),
            .I(N__17537));
    CascadeMux I__3575 (
            .O(N__17540),
            .I(N__17534));
    CascadeMux I__3574 (
            .O(N__17537),
            .I(N__17531));
    CascadeBuf I__3573 (
            .O(N__17534),
            .I(N__17528));
    CascadeBuf I__3572 (
            .O(N__17531),
            .I(N__17525));
    CascadeMux I__3571 (
            .O(N__17528),
            .I(N__17522));
    CascadeMux I__3570 (
            .O(N__17525),
            .I(N__17519));
    CascadeBuf I__3569 (
            .O(N__17522),
            .I(N__17516));
    CascadeBuf I__3568 (
            .O(N__17519),
            .I(N__17513));
    CascadeMux I__3567 (
            .O(N__17516),
            .I(N__17510));
    CascadeMux I__3566 (
            .O(N__17513),
            .I(N__17507));
    CascadeBuf I__3565 (
            .O(N__17510),
            .I(N__17504));
    CascadeBuf I__3564 (
            .O(N__17507),
            .I(N__17501));
    CascadeMux I__3563 (
            .O(N__17504),
            .I(N__17498));
    CascadeMux I__3562 (
            .O(N__17501),
            .I(N__17495));
    CascadeBuf I__3561 (
            .O(N__17498),
            .I(N__17492));
    CascadeBuf I__3560 (
            .O(N__17495),
            .I(N__17489));
    CascadeMux I__3559 (
            .O(N__17492),
            .I(N__17486));
    CascadeMux I__3558 (
            .O(N__17489),
            .I(N__17483));
    CascadeBuf I__3557 (
            .O(N__17486),
            .I(N__17480));
    CascadeBuf I__3556 (
            .O(N__17483),
            .I(N__17477));
    CascadeMux I__3555 (
            .O(N__17480),
            .I(N__17474));
    CascadeMux I__3554 (
            .O(N__17477),
            .I(N__17471));
    CascadeBuf I__3553 (
            .O(N__17474),
            .I(N__17468));
    CascadeBuf I__3552 (
            .O(N__17471),
            .I(N__17465));
    CascadeMux I__3551 (
            .O(N__17468),
            .I(N__17462));
    CascadeMux I__3550 (
            .O(N__17465),
            .I(N__17459));
    CascadeBuf I__3549 (
            .O(N__17462),
            .I(N__17456));
    CascadeBuf I__3548 (
            .O(N__17459),
            .I(N__17453));
    CascadeMux I__3547 (
            .O(N__17456),
            .I(N__17450));
    CascadeMux I__3546 (
            .O(N__17453),
            .I(N__17447));
    CascadeBuf I__3545 (
            .O(N__17450),
            .I(N__17444));
    CascadeBuf I__3544 (
            .O(N__17447),
            .I(N__17441));
    CascadeMux I__3543 (
            .O(N__17444),
            .I(N__17438));
    CascadeMux I__3542 (
            .O(N__17441),
            .I(N__17435));
    CascadeBuf I__3541 (
            .O(N__17438),
            .I(N__17432));
    CascadeBuf I__3540 (
            .O(N__17435),
            .I(N__17429));
    CascadeMux I__3539 (
            .O(N__17432),
            .I(N__17426));
    CascadeMux I__3538 (
            .O(N__17429),
            .I(N__17423));
    CascadeBuf I__3537 (
            .O(N__17426),
            .I(N__17420));
    CascadeBuf I__3536 (
            .O(N__17423),
            .I(N__17417));
    CascadeMux I__3535 (
            .O(N__17420),
            .I(N__17414));
    CascadeMux I__3534 (
            .O(N__17417),
            .I(N__17411));
    CascadeBuf I__3533 (
            .O(N__17414),
            .I(N__17408));
    CascadeBuf I__3532 (
            .O(N__17411),
            .I(N__17405));
    CascadeMux I__3531 (
            .O(N__17408),
            .I(N__17402));
    CascadeMux I__3530 (
            .O(N__17405),
            .I(N__17399));
    CascadeBuf I__3529 (
            .O(N__17402),
            .I(N__17396));
    CascadeBuf I__3528 (
            .O(N__17399),
            .I(N__17393));
    CascadeMux I__3527 (
            .O(N__17396),
            .I(N__17390));
    CascadeMux I__3526 (
            .O(N__17393),
            .I(N__17387));
    CascadeBuf I__3525 (
            .O(N__17390),
            .I(N__17384));
    CascadeBuf I__3524 (
            .O(N__17387),
            .I(N__17381));
    CascadeMux I__3523 (
            .O(N__17384),
            .I(N__17378));
    CascadeMux I__3522 (
            .O(N__17381),
            .I(N__17375));
    InMux I__3521 (
            .O(N__17378),
            .I(N__17372));
    InMux I__3520 (
            .O(N__17375),
            .I(N__17369));
    LocalMux I__3519 (
            .O(N__17372),
            .I(N__17366));
    LocalMux I__3518 (
            .O(N__17369),
            .I(N__17363));
    Span4Mux_s1_v I__3517 (
            .O(N__17366),
            .I(N__17358));
    Span4Mux_s1_v I__3516 (
            .O(N__17363),
            .I(N__17355));
    CascadeMux I__3515 (
            .O(N__17362),
            .I(N__17352));
    CascadeMux I__3514 (
            .O(N__17361),
            .I(N__17349));
    Sp12to4 I__3513 (
            .O(N__17358),
            .I(N__17346));
    Sp12to4 I__3512 (
            .O(N__17355),
            .I(N__17343));
    InMux I__3511 (
            .O(N__17352),
            .I(N__17340));
    InMux I__3510 (
            .O(N__17349),
            .I(N__17337));
    Span12Mux_h I__3509 (
            .O(N__17346),
            .I(N__17332));
    Span12Mux_h I__3508 (
            .O(N__17343),
            .I(N__17332));
    LocalMux I__3507 (
            .O(N__17340),
            .I(N__17329));
    LocalMux I__3506 (
            .O(N__17337),
            .I(N__17324));
    Span12Mux_v I__3505 (
            .O(N__17332),
            .I(N__17324));
    Odrv4 I__3504 (
            .O(N__17329),
            .I(RX_ADDR_4));
    Odrv12 I__3503 (
            .O(N__17324),
            .I(RX_ADDR_4));
    InMux I__3502 (
            .O(N__17319),
            .I(N__17316));
    LocalMux I__3501 (
            .O(N__17316),
            .I(N__17313));
    Odrv4 I__3500 (
            .O(N__17313),
            .I(\receive_module.n129 ));
    CascadeMux I__3499 (
            .O(N__17310),
            .I(N__17306));
    CascadeMux I__3498 (
            .O(N__17309),
            .I(N__17303));
    CascadeBuf I__3497 (
            .O(N__17306),
            .I(N__17300));
    CascadeBuf I__3496 (
            .O(N__17303),
            .I(N__17297));
    CascadeMux I__3495 (
            .O(N__17300),
            .I(N__17294));
    CascadeMux I__3494 (
            .O(N__17297),
            .I(N__17291));
    CascadeBuf I__3493 (
            .O(N__17294),
            .I(N__17288));
    CascadeBuf I__3492 (
            .O(N__17291),
            .I(N__17285));
    CascadeMux I__3491 (
            .O(N__17288),
            .I(N__17282));
    CascadeMux I__3490 (
            .O(N__17285),
            .I(N__17279));
    CascadeBuf I__3489 (
            .O(N__17282),
            .I(N__17276));
    CascadeBuf I__3488 (
            .O(N__17279),
            .I(N__17273));
    CascadeMux I__3487 (
            .O(N__17276),
            .I(N__17270));
    CascadeMux I__3486 (
            .O(N__17273),
            .I(N__17267));
    CascadeBuf I__3485 (
            .O(N__17270),
            .I(N__17264));
    CascadeBuf I__3484 (
            .O(N__17267),
            .I(N__17261));
    CascadeMux I__3483 (
            .O(N__17264),
            .I(N__17258));
    CascadeMux I__3482 (
            .O(N__17261),
            .I(N__17255));
    CascadeBuf I__3481 (
            .O(N__17258),
            .I(N__17252));
    CascadeBuf I__3480 (
            .O(N__17255),
            .I(N__17249));
    CascadeMux I__3479 (
            .O(N__17252),
            .I(N__17246));
    CascadeMux I__3478 (
            .O(N__17249),
            .I(N__17243));
    CascadeBuf I__3477 (
            .O(N__17246),
            .I(N__17240));
    CascadeBuf I__3476 (
            .O(N__17243),
            .I(N__17237));
    CascadeMux I__3475 (
            .O(N__17240),
            .I(N__17234));
    CascadeMux I__3474 (
            .O(N__17237),
            .I(N__17231));
    CascadeBuf I__3473 (
            .O(N__17234),
            .I(N__17228));
    CascadeBuf I__3472 (
            .O(N__17231),
            .I(N__17225));
    CascadeMux I__3471 (
            .O(N__17228),
            .I(N__17222));
    CascadeMux I__3470 (
            .O(N__17225),
            .I(N__17219));
    CascadeBuf I__3469 (
            .O(N__17222),
            .I(N__17216));
    CascadeBuf I__3468 (
            .O(N__17219),
            .I(N__17213));
    CascadeMux I__3467 (
            .O(N__17216),
            .I(N__17210));
    CascadeMux I__3466 (
            .O(N__17213),
            .I(N__17207));
    CascadeBuf I__3465 (
            .O(N__17210),
            .I(N__17204));
    CascadeBuf I__3464 (
            .O(N__17207),
            .I(N__17201));
    CascadeMux I__3463 (
            .O(N__17204),
            .I(N__17198));
    CascadeMux I__3462 (
            .O(N__17201),
            .I(N__17195));
    CascadeBuf I__3461 (
            .O(N__17198),
            .I(N__17192));
    CascadeBuf I__3460 (
            .O(N__17195),
            .I(N__17189));
    CascadeMux I__3459 (
            .O(N__17192),
            .I(N__17186));
    CascadeMux I__3458 (
            .O(N__17189),
            .I(N__17183));
    CascadeBuf I__3457 (
            .O(N__17186),
            .I(N__17180));
    CascadeBuf I__3456 (
            .O(N__17183),
            .I(N__17177));
    CascadeMux I__3455 (
            .O(N__17180),
            .I(N__17174));
    CascadeMux I__3454 (
            .O(N__17177),
            .I(N__17171));
    CascadeBuf I__3453 (
            .O(N__17174),
            .I(N__17168));
    CascadeBuf I__3452 (
            .O(N__17171),
            .I(N__17165));
    CascadeMux I__3451 (
            .O(N__17168),
            .I(N__17162));
    CascadeMux I__3450 (
            .O(N__17165),
            .I(N__17159));
    CascadeBuf I__3449 (
            .O(N__17162),
            .I(N__17156));
    CascadeBuf I__3448 (
            .O(N__17159),
            .I(N__17153));
    CascadeMux I__3447 (
            .O(N__17156),
            .I(N__17150));
    CascadeMux I__3446 (
            .O(N__17153),
            .I(N__17147));
    CascadeBuf I__3445 (
            .O(N__17150),
            .I(N__17144));
    CascadeBuf I__3444 (
            .O(N__17147),
            .I(N__17141));
    CascadeMux I__3443 (
            .O(N__17144),
            .I(N__17138));
    CascadeMux I__3442 (
            .O(N__17141),
            .I(N__17135));
    CascadeBuf I__3441 (
            .O(N__17138),
            .I(N__17132));
    CascadeBuf I__3440 (
            .O(N__17135),
            .I(N__17129));
    CascadeMux I__3439 (
            .O(N__17132),
            .I(N__17126));
    CascadeMux I__3438 (
            .O(N__17129),
            .I(N__17123));
    InMux I__3437 (
            .O(N__17126),
            .I(N__17120));
    InMux I__3436 (
            .O(N__17123),
            .I(N__17117));
    LocalMux I__3435 (
            .O(N__17120),
            .I(N__17113));
    LocalMux I__3434 (
            .O(N__17117),
            .I(N__17110));
    InMux I__3433 (
            .O(N__17116),
            .I(N__17107));
    Span4Mux_h I__3432 (
            .O(N__17113),
            .I(N__17104));
    Span4Mux_h I__3431 (
            .O(N__17110),
            .I(N__17101));
    LocalMux I__3430 (
            .O(N__17107),
            .I(N__17097));
    Sp12to4 I__3429 (
            .O(N__17104),
            .I(N__17094));
    Sp12to4 I__3428 (
            .O(N__17101),
            .I(N__17091));
    InMux I__3427 (
            .O(N__17100),
            .I(N__17088));
    Span12Mux_v I__3426 (
            .O(N__17097),
            .I(N__17083));
    Span12Mux_v I__3425 (
            .O(N__17094),
            .I(N__17083));
    Span12Mux_v I__3424 (
            .O(N__17091),
            .I(N__17080));
    LocalMux I__3423 (
            .O(N__17088),
            .I(RX_ADDR_8));
    Odrv12 I__3422 (
            .O(N__17083),
            .I(RX_ADDR_8));
    Odrv12 I__3421 (
            .O(N__17080),
            .I(RX_ADDR_8));
    InMux I__3420 (
            .O(N__17073),
            .I(N__17070));
    LocalMux I__3419 (
            .O(N__17070),
            .I(N__17067));
    Span4Mux_h I__3418 (
            .O(N__17067),
            .I(N__17064));
    Odrv4 I__3417 (
            .O(N__17064),
            .I(\receive_module.n131 ));
    CascadeMux I__3416 (
            .O(N__17061),
            .I(N__17057));
    CascadeMux I__3415 (
            .O(N__17060),
            .I(N__17054));
    CascadeBuf I__3414 (
            .O(N__17057),
            .I(N__17051));
    CascadeBuf I__3413 (
            .O(N__17054),
            .I(N__17048));
    CascadeMux I__3412 (
            .O(N__17051),
            .I(N__17045));
    CascadeMux I__3411 (
            .O(N__17048),
            .I(N__17042));
    CascadeBuf I__3410 (
            .O(N__17045),
            .I(N__17039));
    CascadeBuf I__3409 (
            .O(N__17042),
            .I(N__17036));
    CascadeMux I__3408 (
            .O(N__17039),
            .I(N__17033));
    CascadeMux I__3407 (
            .O(N__17036),
            .I(N__17030));
    CascadeBuf I__3406 (
            .O(N__17033),
            .I(N__17027));
    CascadeBuf I__3405 (
            .O(N__17030),
            .I(N__17024));
    CascadeMux I__3404 (
            .O(N__17027),
            .I(N__17021));
    CascadeMux I__3403 (
            .O(N__17024),
            .I(N__17018));
    CascadeBuf I__3402 (
            .O(N__17021),
            .I(N__17015));
    CascadeBuf I__3401 (
            .O(N__17018),
            .I(N__17012));
    CascadeMux I__3400 (
            .O(N__17015),
            .I(N__17009));
    CascadeMux I__3399 (
            .O(N__17012),
            .I(N__17006));
    CascadeBuf I__3398 (
            .O(N__17009),
            .I(N__17003));
    CascadeBuf I__3397 (
            .O(N__17006),
            .I(N__17000));
    CascadeMux I__3396 (
            .O(N__17003),
            .I(N__16997));
    CascadeMux I__3395 (
            .O(N__17000),
            .I(N__16994));
    CascadeBuf I__3394 (
            .O(N__16997),
            .I(N__16991));
    CascadeBuf I__3393 (
            .O(N__16994),
            .I(N__16988));
    CascadeMux I__3392 (
            .O(N__16991),
            .I(N__16985));
    CascadeMux I__3391 (
            .O(N__16988),
            .I(N__16982));
    CascadeBuf I__3390 (
            .O(N__16985),
            .I(N__16979));
    CascadeBuf I__3389 (
            .O(N__16982),
            .I(N__16976));
    CascadeMux I__3388 (
            .O(N__16979),
            .I(N__16973));
    CascadeMux I__3387 (
            .O(N__16976),
            .I(N__16970));
    CascadeBuf I__3386 (
            .O(N__16973),
            .I(N__16967));
    CascadeBuf I__3385 (
            .O(N__16970),
            .I(N__16964));
    CascadeMux I__3384 (
            .O(N__16967),
            .I(N__16961));
    CascadeMux I__3383 (
            .O(N__16964),
            .I(N__16958));
    CascadeBuf I__3382 (
            .O(N__16961),
            .I(N__16955));
    CascadeBuf I__3381 (
            .O(N__16958),
            .I(N__16952));
    CascadeMux I__3380 (
            .O(N__16955),
            .I(N__16949));
    CascadeMux I__3379 (
            .O(N__16952),
            .I(N__16946));
    CascadeBuf I__3378 (
            .O(N__16949),
            .I(N__16943));
    CascadeBuf I__3377 (
            .O(N__16946),
            .I(N__16940));
    CascadeMux I__3376 (
            .O(N__16943),
            .I(N__16937));
    CascadeMux I__3375 (
            .O(N__16940),
            .I(N__16934));
    CascadeBuf I__3374 (
            .O(N__16937),
            .I(N__16931));
    CascadeBuf I__3373 (
            .O(N__16934),
            .I(N__16928));
    CascadeMux I__3372 (
            .O(N__16931),
            .I(N__16925));
    CascadeMux I__3371 (
            .O(N__16928),
            .I(N__16922));
    CascadeBuf I__3370 (
            .O(N__16925),
            .I(N__16919));
    CascadeBuf I__3369 (
            .O(N__16922),
            .I(N__16916));
    CascadeMux I__3368 (
            .O(N__16919),
            .I(N__16913));
    CascadeMux I__3367 (
            .O(N__16916),
            .I(N__16910));
    CascadeBuf I__3366 (
            .O(N__16913),
            .I(N__16907));
    CascadeBuf I__3365 (
            .O(N__16910),
            .I(N__16904));
    CascadeMux I__3364 (
            .O(N__16907),
            .I(N__16901));
    CascadeMux I__3363 (
            .O(N__16904),
            .I(N__16898));
    CascadeBuf I__3362 (
            .O(N__16901),
            .I(N__16895));
    CascadeBuf I__3361 (
            .O(N__16898),
            .I(N__16892));
    CascadeMux I__3360 (
            .O(N__16895),
            .I(N__16889));
    CascadeMux I__3359 (
            .O(N__16892),
            .I(N__16886));
    CascadeBuf I__3358 (
            .O(N__16889),
            .I(N__16883));
    CascadeBuf I__3357 (
            .O(N__16886),
            .I(N__16880));
    CascadeMux I__3356 (
            .O(N__16883),
            .I(N__16877));
    CascadeMux I__3355 (
            .O(N__16880),
            .I(N__16874));
    InMux I__3354 (
            .O(N__16877),
            .I(N__16871));
    InMux I__3353 (
            .O(N__16874),
            .I(N__16868));
    LocalMux I__3352 (
            .O(N__16871),
            .I(N__16865));
    LocalMux I__3351 (
            .O(N__16868),
            .I(N__16861));
    Span4Mux_s1_v I__3350 (
            .O(N__16865),
            .I(N__16858));
    InMux I__3349 (
            .O(N__16864),
            .I(N__16854));
    Span4Mux_s1_v I__3348 (
            .O(N__16861),
            .I(N__16851));
    Sp12to4 I__3347 (
            .O(N__16858),
            .I(N__16848));
    CascadeMux I__3346 (
            .O(N__16857),
            .I(N__16845));
    LocalMux I__3345 (
            .O(N__16854),
            .I(N__16842));
    Sp12to4 I__3344 (
            .O(N__16851),
            .I(N__16839));
    Span12Mux_h I__3343 (
            .O(N__16848),
            .I(N__16836));
    InMux I__3342 (
            .O(N__16845),
            .I(N__16833));
    Span4Mux_h I__3341 (
            .O(N__16842),
            .I(N__16830));
    Span12Mux_v I__3340 (
            .O(N__16839),
            .I(N__16825));
    Span12Mux_v I__3339 (
            .O(N__16836),
            .I(N__16825));
    LocalMux I__3338 (
            .O(N__16833),
            .I(RX_ADDR_6));
    Odrv4 I__3337 (
            .O(N__16830),
            .I(RX_ADDR_6));
    Odrv12 I__3336 (
            .O(N__16825),
            .I(RX_ADDR_6));
    InMux I__3335 (
            .O(N__16818),
            .I(N__16815));
    LocalMux I__3334 (
            .O(N__16815),
            .I(N__16812));
    Odrv4 I__3333 (
            .O(N__16812),
            .I(\receive_module.n130 ));
    CascadeMux I__3332 (
            .O(N__16809),
            .I(N__16805));
    CascadeMux I__3331 (
            .O(N__16808),
            .I(N__16802));
    CascadeBuf I__3330 (
            .O(N__16805),
            .I(N__16799));
    CascadeBuf I__3329 (
            .O(N__16802),
            .I(N__16796));
    CascadeMux I__3328 (
            .O(N__16799),
            .I(N__16793));
    CascadeMux I__3327 (
            .O(N__16796),
            .I(N__16790));
    CascadeBuf I__3326 (
            .O(N__16793),
            .I(N__16787));
    CascadeBuf I__3325 (
            .O(N__16790),
            .I(N__16784));
    CascadeMux I__3324 (
            .O(N__16787),
            .I(N__16781));
    CascadeMux I__3323 (
            .O(N__16784),
            .I(N__16778));
    CascadeBuf I__3322 (
            .O(N__16781),
            .I(N__16775));
    CascadeBuf I__3321 (
            .O(N__16778),
            .I(N__16772));
    CascadeMux I__3320 (
            .O(N__16775),
            .I(N__16769));
    CascadeMux I__3319 (
            .O(N__16772),
            .I(N__16766));
    CascadeBuf I__3318 (
            .O(N__16769),
            .I(N__16763));
    CascadeBuf I__3317 (
            .O(N__16766),
            .I(N__16760));
    CascadeMux I__3316 (
            .O(N__16763),
            .I(N__16757));
    CascadeMux I__3315 (
            .O(N__16760),
            .I(N__16754));
    CascadeBuf I__3314 (
            .O(N__16757),
            .I(N__16751));
    CascadeBuf I__3313 (
            .O(N__16754),
            .I(N__16748));
    CascadeMux I__3312 (
            .O(N__16751),
            .I(N__16745));
    CascadeMux I__3311 (
            .O(N__16748),
            .I(N__16742));
    CascadeBuf I__3310 (
            .O(N__16745),
            .I(N__16739));
    CascadeBuf I__3309 (
            .O(N__16742),
            .I(N__16736));
    CascadeMux I__3308 (
            .O(N__16739),
            .I(N__16733));
    CascadeMux I__3307 (
            .O(N__16736),
            .I(N__16730));
    CascadeBuf I__3306 (
            .O(N__16733),
            .I(N__16727));
    CascadeBuf I__3305 (
            .O(N__16730),
            .I(N__16724));
    CascadeMux I__3304 (
            .O(N__16727),
            .I(N__16721));
    CascadeMux I__3303 (
            .O(N__16724),
            .I(N__16718));
    CascadeBuf I__3302 (
            .O(N__16721),
            .I(N__16715));
    CascadeBuf I__3301 (
            .O(N__16718),
            .I(N__16712));
    CascadeMux I__3300 (
            .O(N__16715),
            .I(N__16709));
    CascadeMux I__3299 (
            .O(N__16712),
            .I(N__16706));
    CascadeBuf I__3298 (
            .O(N__16709),
            .I(N__16703));
    CascadeBuf I__3297 (
            .O(N__16706),
            .I(N__16700));
    CascadeMux I__3296 (
            .O(N__16703),
            .I(N__16697));
    CascadeMux I__3295 (
            .O(N__16700),
            .I(N__16694));
    CascadeBuf I__3294 (
            .O(N__16697),
            .I(N__16691));
    CascadeBuf I__3293 (
            .O(N__16694),
            .I(N__16688));
    CascadeMux I__3292 (
            .O(N__16691),
            .I(N__16685));
    CascadeMux I__3291 (
            .O(N__16688),
            .I(N__16682));
    CascadeBuf I__3290 (
            .O(N__16685),
            .I(N__16679));
    CascadeBuf I__3289 (
            .O(N__16682),
            .I(N__16676));
    CascadeMux I__3288 (
            .O(N__16679),
            .I(N__16673));
    CascadeMux I__3287 (
            .O(N__16676),
            .I(N__16670));
    CascadeBuf I__3286 (
            .O(N__16673),
            .I(N__16667));
    CascadeBuf I__3285 (
            .O(N__16670),
            .I(N__16664));
    CascadeMux I__3284 (
            .O(N__16667),
            .I(N__16661));
    CascadeMux I__3283 (
            .O(N__16664),
            .I(N__16658));
    CascadeBuf I__3282 (
            .O(N__16661),
            .I(N__16655));
    CascadeBuf I__3281 (
            .O(N__16658),
            .I(N__16652));
    CascadeMux I__3280 (
            .O(N__16655),
            .I(N__16649));
    CascadeMux I__3279 (
            .O(N__16652),
            .I(N__16646));
    CascadeBuf I__3278 (
            .O(N__16649),
            .I(N__16643));
    CascadeBuf I__3277 (
            .O(N__16646),
            .I(N__16640));
    CascadeMux I__3276 (
            .O(N__16643),
            .I(N__16637));
    CascadeMux I__3275 (
            .O(N__16640),
            .I(N__16634));
    CascadeBuf I__3274 (
            .O(N__16637),
            .I(N__16631));
    CascadeBuf I__3273 (
            .O(N__16634),
            .I(N__16628));
    CascadeMux I__3272 (
            .O(N__16631),
            .I(N__16625));
    CascadeMux I__3271 (
            .O(N__16628),
            .I(N__16622));
    InMux I__3270 (
            .O(N__16625),
            .I(N__16619));
    InMux I__3269 (
            .O(N__16622),
            .I(N__16615));
    LocalMux I__3268 (
            .O(N__16619),
            .I(N__16612));
    InMux I__3267 (
            .O(N__16618),
            .I(N__16609));
    LocalMux I__3266 (
            .O(N__16615),
            .I(N__16606));
    Span4Mux_h I__3265 (
            .O(N__16612),
            .I(N__16603));
    LocalMux I__3264 (
            .O(N__16609),
            .I(N__16600));
    Span12Mux_s1_v I__3263 (
            .O(N__16606),
            .I(N__16596));
    Sp12to4 I__3262 (
            .O(N__16603),
            .I(N__16593));
    Span4Mux_h I__3261 (
            .O(N__16600),
            .I(N__16590));
    InMux I__3260 (
            .O(N__16599),
            .I(N__16587));
    Span12Mux_v I__3259 (
            .O(N__16596),
            .I(N__16584));
    Span12Mux_v I__3258 (
            .O(N__16593),
            .I(N__16581));
    Odrv4 I__3257 (
            .O(N__16590),
            .I(RX_ADDR_7));
    LocalMux I__3256 (
            .O(N__16587),
            .I(RX_ADDR_7));
    Odrv12 I__3255 (
            .O(N__16584),
            .I(RX_ADDR_7));
    Odrv12 I__3254 (
            .O(N__16581),
            .I(RX_ADDR_7));
    InMux I__3253 (
            .O(N__16572),
            .I(N__16569));
    LocalMux I__3252 (
            .O(N__16569),
            .I(N__16566));
    Span4Mux_v I__3251 (
            .O(N__16566),
            .I(N__16563));
    Span4Mux_h I__3250 (
            .O(N__16563),
            .I(N__16560));
    Span4Mux_h I__3249 (
            .O(N__16560),
            .I(N__16557));
    Span4Mux_v I__3248 (
            .O(N__16557),
            .I(N__16554));
    Odrv4 I__3247 (
            .O(N__16554),
            .I(\line_buffer.n564 ));
    InMux I__3246 (
            .O(N__16551),
            .I(N__16548));
    LocalMux I__3245 (
            .O(N__16548),
            .I(N__16545));
    Span4Mux_v I__3244 (
            .O(N__16545),
            .I(N__16542));
    Span4Mux_h I__3243 (
            .O(N__16542),
            .I(N__16539));
    Span4Mux_h I__3242 (
            .O(N__16539),
            .I(N__16536));
    Odrv4 I__3241 (
            .O(N__16536),
            .I(\line_buffer.n556 ));
    SRMux I__3240 (
            .O(N__16533),
            .I(N__16529));
    SRMux I__3239 (
            .O(N__16532),
            .I(N__16524));
    LocalMux I__3238 (
            .O(N__16529),
            .I(N__16521));
    SRMux I__3237 (
            .O(N__16528),
            .I(N__16518));
    SRMux I__3236 (
            .O(N__16527),
            .I(N__16515));
    LocalMux I__3235 (
            .O(N__16524),
            .I(N__16512));
    Span4Mux_h I__3234 (
            .O(N__16521),
            .I(N__16509));
    LocalMux I__3233 (
            .O(N__16518),
            .I(N__16506));
    LocalMux I__3232 (
            .O(N__16515),
            .I(N__16503));
    Span4Mux_h I__3231 (
            .O(N__16512),
            .I(N__16500));
    Span4Mux_h I__3230 (
            .O(N__16509),
            .I(N__16497));
    Span4Mux_h I__3229 (
            .O(N__16506),
            .I(N__16492));
    Span4Mux_v I__3228 (
            .O(N__16503),
            .I(N__16492));
    Sp12to4 I__3227 (
            .O(N__16500),
            .I(N__16489));
    Sp12to4 I__3226 (
            .O(N__16497),
            .I(N__16486));
    Sp12to4 I__3225 (
            .O(N__16492),
            .I(N__16481));
    Span12Mux_s5_v I__3224 (
            .O(N__16489),
            .I(N__16481));
    Span12Mux_v I__3223 (
            .O(N__16486),
            .I(N__16476));
    Span12Mux_v I__3222 (
            .O(N__16481),
            .I(N__16476));
    Odrv12 I__3221 (
            .O(N__16476),
            .I(\line_buffer.n473 ));
    SRMux I__3220 (
            .O(N__16473),
            .I(N__16470));
    LocalMux I__3219 (
            .O(N__16470),
            .I(N__16467));
    Span4Mux_v I__3218 (
            .O(N__16467),
            .I(N__16461));
    SRMux I__3217 (
            .O(N__16466),
            .I(N__16458));
    SRMux I__3216 (
            .O(N__16465),
            .I(N__16455));
    SRMux I__3215 (
            .O(N__16464),
            .I(N__16452));
    Span4Mux_v I__3214 (
            .O(N__16461),
            .I(N__16447));
    LocalMux I__3213 (
            .O(N__16458),
            .I(N__16447));
    LocalMux I__3212 (
            .O(N__16455),
            .I(N__16442));
    LocalMux I__3211 (
            .O(N__16452),
            .I(N__16442));
    Span4Mux_v I__3210 (
            .O(N__16447),
            .I(N__16437));
    Span4Mux_v I__3209 (
            .O(N__16442),
            .I(N__16437));
    Span4Mux_h I__3208 (
            .O(N__16437),
            .I(N__16434));
    Span4Mux_h I__3207 (
            .O(N__16434),
            .I(N__16431));
    Odrv4 I__3206 (
            .O(N__16431),
            .I(\line_buffer.n570 ));
    SRMux I__3205 (
            .O(N__16428),
            .I(N__16424));
    SRMux I__3204 (
            .O(N__16427),
            .I(N__16420));
    LocalMux I__3203 (
            .O(N__16424),
            .I(N__16417));
    SRMux I__3202 (
            .O(N__16423),
            .I(N__16414));
    LocalMux I__3201 (
            .O(N__16420),
            .I(N__16410));
    Span4Mux_h I__3200 (
            .O(N__16417),
            .I(N__16405));
    LocalMux I__3199 (
            .O(N__16414),
            .I(N__16405));
    SRMux I__3198 (
            .O(N__16413),
            .I(N__16402));
    Span4Mux_v I__3197 (
            .O(N__16410),
            .I(N__16399));
    Span4Mux_v I__3196 (
            .O(N__16405),
            .I(N__16394));
    LocalMux I__3195 (
            .O(N__16402),
            .I(N__16394));
    Sp12to4 I__3194 (
            .O(N__16399),
            .I(N__16391));
    Span4Mux_h I__3193 (
            .O(N__16394),
            .I(N__16388));
    Span12Mux_h I__3192 (
            .O(N__16391),
            .I(N__16385));
    Span4Mux_h I__3191 (
            .O(N__16388),
            .I(N__16382));
    Odrv12 I__3190 (
            .O(N__16385),
            .I(\line_buffer.n571 ));
    Odrv4 I__3189 (
            .O(N__16382),
            .I(\line_buffer.n571 ));
    InMux I__3188 (
            .O(N__16377),
            .I(N__16374));
    LocalMux I__3187 (
            .O(N__16374),
            .I(N__16371));
    Span4Mux_h I__3186 (
            .O(N__16371),
            .I(N__16368));
    Odrv4 I__3185 (
            .O(N__16368),
            .I(\transmit_module.ADDR_Y_COMPONENT_11 ));
    InMux I__3184 (
            .O(N__16365),
            .I(N__16362));
    LocalMux I__3183 (
            .O(N__16362),
            .I(N__16359));
    Odrv4 I__3182 (
            .O(N__16359),
            .I(\transmit_module.n121 ));
    InMux I__3181 (
            .O(N__16356),
            .I(N__16353));
    LocalMux I__3180 (
            .O(N__16353),
            .I(N__16350));
    Span4Mux_h I__3179 (
            .O(N__16350),
            .I(N__16347));
    Odrv4 I__3178 (
            .O(N__16347),
            .I(\transmit_module.ADDR_Y_COMPONENT_13 ));
    InMux I__3177 (
            .O(N__16344),
            .I(N__16341));
    LocalMux I__3176 (
            .O(N__16341),
            .I(N__16338));
    Odrv4 I__3175 (
            .O(N__16338),
            .I(\transmit_module.n119 ));
    InMux I__3174 (
            .O(N__16335),
            .I(N__16332));
    LocalMux I__3173 (
            .O(N__16332),
            .I(N__16329));
    Span4Mux_v I__3172 (
            .O(N__16329),
            .I(N__16326));
    Odrv4 I__3171 (
            .O(N__16326),
            .I(\transmit_module.ADDR_Y_COMPONENT_12 ));
    InMux I__3170 (
            .O(N__16323),
            .I(N__16309));
    InMux I__3169 (
            .O(N__16322),
            .I(N__16309));
    InMux I__3168 (
            .O(N__16321),
            .I(N__16301));
    InMux I__3167 (
            .O(N__16320),
            .I(N__16291));
    InMux I__3166 (
            .O(N__16319),
            .I(N__16291));
    InMux I__3165 (
            .O(N__16318),
            .I(N__16291));
    InMux I__3164 (
            .O(N__16317),
            .I(N__16282));
    InMux I__3163 (
            .O(N__16316),
            .I(N__16282));
    InMux I__3162 (
            .O(N__16315),
            .I(N__16282));
    InMux I__3161 (
            .O(N__16314),
            .I(N__16282));
    LocalMux I__3160 (
            .O(N__16309),
            .I(N__16279));
    InMux I__3159 (
            .O(N__16308),
            .I(N__16276));
    InMux I__3158 (
            .O(N__16307),
            .I(N__16267));
    InMux I__3157 (
            .O(N__16306),
            .I(N__16267));
    InMux I__3156 (
            .O(N__16305),
            .I(N__16267));
    InMux I__3155 (
            .O(N__16304),
            .I(N__16267));
    LocalMux I__3154 (
            .O(N__16301),
            .I(N__16261));
    InMux I__3153 (
            .O(N__16300),
            .I(N__16254));
    InMux I__3152 (
            .O(N__16299),
            .I(N__16254));
    InMux I__3151 (
            .O(N__16298),
            .I(N__16254));
    LocalMux I__3150 (
            .O(N__16291),
            .I(N__16251));
    LocalMux I__3149 (
            .O(N__16282),
            .I(N__16242));
    Span4Mux_v I__3148 (
            .O(N__16279),
            .I(N__16242));
    LocalMux I__3147 (
            .O(N__16276),
            .I(N__16242));
    LocalMux I__3146 (
            .O(N__16267),
            .I(N__16242));
    CascadeMux I__3145 (
            .O(N__16266),
            .I(N__16234));
    InMux I__3144 (
            .O(N__16265),
            .I(N__16230));
    InMux I__3143 (
            .O(N__16264),
            .I(N__16227));
    Sp12to4 I__3142 (
            .O(N__16261),
            .I(N__16222));
    LocalMux I__3141 (
            .O(N__16254),
            .I(N__16222));
    Span4Mux_v I__3140 (
            .O(N__16251),
            .I(N__16217));
    Span4Mux_v I__3139 (
            .O(N__16242),
            .I(N__16217));
    InMux I__3138 (
            .O(N__16241),
            .I(N__16210));
    InMux I__3137 (
            .O(N__16240),
            .I(N__16210));
    InMux I__3136 (
            .O(N__16239),
            .I(N__16210));
    InMux I__3135 (
            .O(N__16238),
            .I(N__16201));
    InMux I__3134 (
            .O(N__16237),
            .I(N__16201));
    InMux I__3133 (
            .O(N__16234),
            .I(N__16201));
    InMux I__3132 (
            .O(N__16233),
            .I(N__16201));
    LocalMux I__3131 (
            .O(N__16230),
            .I(\transmit_module.n3675 ));
    LocalMux I__3130 (
            .O(N__16227),
            .I(\transmit_module.n3675 ));
    Odrv12 I__3129 (
            .O(N__16222),
            .I(\transmit_module.n3675 ));
    Odrv4 I__3128 (
            .O(N__16217),
            .I(\transmit_module.n3675 ));
    LocalMux I__3127 (
            .O(N__16210),
            .I(\transmit_module.n3675 ));
    LocalMux I__3126 (
            .O(N__16201),
            .I(\transmit_module.n3675 ));
    InMux I__3125 (
            .O(N__16188),
            .I(N__16185));
    LocalMux I__3124 (
            .O(N__16185),
            .I(N__16182));
    Odrv4 I__3123 (
            .O(N__16182),
            .I(\transmit_module.n120 ));
    CEMux I__3122 (
            .O(N__16179),
            .I(N__16176));
    LocalMux I__3121 (
            .O(N__16176),
            .I(N__16173));
    Span4Mux_v I__3120 (
            .O(N__16173),
            .I(N__16170));
    Span4Mux_h I__3119 (
            .O(N__16170),
            .I(N__16167));
    Odrv4 I__3118 (
            .O(N__16167),
            .I(\transmit_module.n2070 ));
    CEMux I__3117 (
            .O(N__16164),
            .I(N__16161));
    LocalMux I__3116 (
            .O(N__16161),
            .I(N__16158));
    Span4Mux_v I__3115 (
            .O(N__16158),
            .I(N__16155));
    Odrv4 I__3114 (
            .O(N__16155),
            .I(\receive_module.n3671 ));
    SRMux I__3113 (
            .O(N__16152),
            .I(N__16149));
    LocalMux I__3112 (
            .O(N__16149),
            .I(N__16145));
    SRMux I__3111 (
            .O(N__16148),
            .I(N__16142));
    Span4Mux_v I__3110 (
            .O(N__16145),
            .I(N__16135));
    LocalMux I__3109 (
            .O(N__16142),
            .I(N__16135));
    SRMux I__3108 (
            .O(N__16141),
            .I(N__16132));
    SRMux I__3107 (
            .O(N__16140),
            .I(N__16129));
    Span4Mux_v I__3106 (
            .O(N__16135),
            .I(N__16124));
    LocalMux I__3105 (
            .O(N__16132),
            .I(N__16124));
    LocalMux I__3104 (
            .O(N__16129),
            .I(N__16121));
    Span4Mux_h I__3103 (
            .O(N__16124),
            .I(N__16118));
    Span4Mux_h I__3102 (
            .O(N__16121),
            .I(N__16115));
    Span4Mux_h I__3101 (
            .O(N__16118),
            .I(N__16112));
    Span4Mux_h I__3100 (
            .O(N__16115),
            .I(N__16107));
    Span4Mux_h I__3099 (
            .O(N__16112),
            .I(N__16107));
    Odrv4 I__3098 (
            .O(N__16107),
            .I(\line_buffer.n603 ));
    SRMux I__3097 (
            .O(N__16104),
            .I(N__16100));
    SRMux I__3096 (
            .O(N__16103),
            .I(N__16097));
    LocalMux I__3095 (
            .O(N__16100),
            .I(N__16091));
    LocalMux I__3094 (
            .O(N__16097),
            .I(N__16091));
    SRMux I__3093 (
            .O(N__16096),
            .I(N__16088));
    Span4Mux_v I__3092 (
            .O(N__16091),
            .I(N__16082));
    LocalMux I__3091 (
            .O(N__16088),
            .I(N__16082));
    SRMux I__3090 (
            .O(N__16087),
            .I(N__16079));
    Span4Mux_v I__3089 (
            .O(N__16082),
            .I(N__16076));
    LocalMux I__3088 (
            .O(N__16079),
            .I(N__16073));
    Span4Mux_v I__3087 (
            .O(N__16076),
            .I(N__16070));
    Span4Mux_v I__3086 (
            .O(N__16073),
            .I(N__16067));
    Span4Mux_h I__3085 (
            .O(N__16070),
            .I(N__16064));
    Span4Mux_h I__3084 (
            .O(N__16067),
            .I(N__16061));
    Span4Mux_h I__3083 (
            .O(N__16064),
            .I(N__16058));
    Span4Mux_h I__3082 (
            .O(N__16061),
            .I(N__16055));
    Odrv4 I__3081 (
            .O(N__16058),
            .I(\line_buffer.n539 ));
    Odrv4 I__3080 (
            .O(N__16055),
            .I(\line_buffer.n539 ));
    InMux I__3079 (
            .O(N__16050),
            .I(\receive_module.rx_counter.n3205 ));
    InMux I__3078 (
            .O(N__16047),
            .I(\receive_module.rx_counter.n3206 ));
    InMux I__3077 (
            .O(N__16044),
            .I(N__16041));
    LocalMux I__3076 (
            .O(N__16041),
            .I(\receive_module.rx_counter.n6 ));
    InMux I__3075 (
            .O(N__16038),
            .I(N__16035));
    LocalMux I__3074 (
            .O(N__16035),
            .I(\receive_module.rx_counter.n7 ));
    InMux I__3073 (
            .O(N__16032),
            .I(N__16028));
    InMux I__3072 (
            .O(N__16031),
            .I(N__16025));
    LocalMux I__3071 (
            .O(N__16028),
            .I(\receive_module.rx_counter.FRAME_COUNTER_5 ));
    LocalMux I__3070 (
            .O(N__16025),
            .I(\receive_module.rx_counter.FRAME_COUNTER_5 ));
    InMux I__3069 (
            .O(N__16020),
            .I(N__16016));
    InMux I__3068 (
            .O(N__16019),
            .I(N__16013));
    LocalMux I__3067 (
            .O(N__16016),
            .I(\receive_module.rx_counter.FRAME_COUNTER_1 ));
    LocalMux I__3066 (
            .O(N__16013),
            .I(\receive_module.rx_counter.FRAME_COUNTER_1 ));
    InMux I__3065 (
            .O(N__16008),
            .I(N__16005));
    LocalMux I__3064 (
            .O(N__16005),
            .I(N__16000));
    InMux I__3063 (
            .O(N__16004),
            .I(N__15997));
    InMux I__3062 (
            .O(N__16003),
            .I(N__15994));
    Span4Mux_v I__3061 (
            .O(N__16000),
            .I(N__15991));
    LocalMux I__3060 (
            .O(N__15997),
            .I(N__15988));
    LocalMux I__3059 (
            .O(N__15994),
            .I(\receive_module.rx_counter.X_3 ));
    Odrv4 I__3058 (
            .O(N__15991),
            .I(\receive_module.rx_counter.X_3 ));
    Odrv4 I__3057 (
            .O(N__15988),
            .I(\receive_module.rx_counter.X_3 ));
    InMux I__3056 (
            .O(N__15981),
            .I(N__15978));
    LocalMux I__3055 (
            .O(N__15978),
            .I(N__15973));
    InMux I__3054 (
            .O(N__15977),
            .I(N__15970));
    InMux I__3053 (
            .O(N__15976),
            .I(N__15967));
    Span4Mux_v I__3052 (
            .O(N__15973),
            .I(N__15964));
    LocalMux I__3051 (
            .O(N__15970),
            .I(N__15961));
    LocalMux I__3050 (
            .O(N__15967),
            .I(\receive_module.rx_counter.X_5 ));
    Odrv4 I__3049 (
            .O(N__15964),
            .I(\receive_module.rx_counter.X_5 ));
    Odrv4 I__3048 (
            .O(N__15961),
            .I(\receive_module.rx_counter.X_5 ));
    CascadeMux I__3047 (
            .O(N__15954),
            .I(N__15951));
    InMux I__3046 (
            .O(N__15951),
            .I(N__15947));
    InMux I__3045 (
            .O(N__15950),
            .I(N__15943));
    LocalMux I__3044 (
            .O(N__15947),
            .I(N__15940));
    InMux I__3043 (
            .O(N__15946),
            .I(N__15937));
    LocalMux I__3042 (
            .O(N__15943),
            .I(N__15934));
    Span4Mux_v I__3041 (
            .O(N__15940),
            .I(N__15931));
    LocalMux I__3040 (
            .O(N__15937),
            .I(\receive_module.rx_counter.X_4 ));
    Odrv4 I__3039 (
            .O(N__15934),
            .I(\receive_module.rx_counter.X_4 ));
    Odrv4 I__3038 (
            .O(N__15931),
            .I(\receive_module.rx_counter.X_4 ));
    InMux I__3037 (
            .O(N__15924),
            .I(N__15920));
    InMux I__3036 (
            .O(N__15923),
            .I(N__15917));
    LocalMux I__3035 (
            .O(N__15920),
            .I(N__15912));
    LocalMux I__3034 (
            .O(N__15917),
            .I(N__15912));
    Odrv4 I__3033 (
            .O(N__15912),
            .I(\receive_module.rx_counter.n3222 ));
    CascadeMux I__3032 (
            .O(N__15909),
            .I(N__15905));
    InMux I__3031 (
            .O(N__15908),
            .I(N__15902));
    InMux I__3030 (
            .O(N__15905),
            .I(N__15898));
    LocalMux I__3029 (
            .O(N__15902),
            .I(N__15895));
    InMux I__3028 (
            .O(N__15901),
            .I(N__15892));
    LocalMux I__3027 (
            .O(N__15898),
            .I(N__15889));
    Span4Mux_v I__3026 (
            .O(N__15895),
            .I(N__15886));
    LocalMux I__3025 (
            .O(N__15892),
            .I(\receive_module.rx_counter.X_7 ));
    Odrv4 I__3024 (
            .O(N__15889),
            .I(\receive_module.rx_counter.X_7 ));
    Odrv4 I__3023 (
            .O(N__15886),
            .I(\receive_module.rx_counter.X_7 ));
    CascadeMux I__3022 (
            .O(N__15879),
            .I(\receive_module.rx_counter.n3455_cascade_ ));
    InMux I__3021 (
            .O(N__15876),
            .I(N__15873));
    LocalMux I__3020 (
            .O(N__15873),
            .I(N__15868));
    InMux I__3019 (
            .O(N__15872),
            .I(N__15865));
    InMux I__3018 (
            .O(N__15871),
            .I(N__15862));
    Span4Mux_v I__3017 (
            .O(N__15868),
            .I(N__15859));
    LocalMux I__3016 (
            .O(N__15865),
            .I(N__15856));
    LocalMux I__3015 (
            .O(N__15862),
            .I(\receive_module.rx_counter.X_6 ));
    Odrv4 I__3014 (
            .O(N__15859),
            .I(\receive_module.rx_counter.X_6 ));
    Odrv4 I__3013 (
            .O(N__15856),
            .I(\receive_module.rx_counter.X_6 ));
    InMux I__3012 (
            .O(N__15849),
            .I(N__15843));
    InMux I__3011 (
            .O(N__15848),
            .I(N__15843));
    LocalMux I__3010 (
            .O(N__15843),
            .I(N__15839));
    InMux I__3009 (
            .O(N__15842),
            .I(N__15836));
    Span4Mux_v I__3008 (
            .O(N__15839),
            .I(N__15833));
    LocalMux I__3007 (
            .O(N__15836),
            .I(\receive_module.rx_counter.X_8 ));
    Odrv4 I__3006 (
            .O(N__15833),
            .I(\receive_module.rx_counter.X_8 ));
    InMux I__3005 (
            .O(N__15828),
            .I(N__15825));
    LocalMux I__3004 (
            .O(N__15825),
            .I(N__15821));
    InMux I__3003 (
            .O(N__15824),
            .I(N__15818));
    Span4Mux_v I__3002 (
            .O(N__15821),
            .I(N__15815));
    LocalMux I__3001 (
            .O(N__15818),
            .I(\receive_module.rx_counter.X_9 ));
    Odrv4 I__3000 (
            .O(N__15815),
            .I(\receive_module.rx_counter.X_9 ));
    CascadeMux I__2999 (
            .O(N__15810),
            .I(\receive_module.rx_counter.n39_cascade_ ));
    InMux I__2998 (
            .O(N__15807),
            .I(N__15804));
    LocalMux I__2997 (
            .O(N__15804),
            .I(\receive_module.rx_counter.n3426 ));
    InMux I__2996 (
            .O(N__15801),
            .I(N__15798));
    LocalMux I__2995 (
            .O(N__15798),
            .I(N__15795));
    Odrv12 I__2994 (
            .O(N__15795),
            .I(\receive_module.rx_counter.n3478 ));
    CascadeMux I__2993 (
            .O(N__15792),
            .I(\receive_module.rx_counter.n54_cascade_ ));
    InMux I__2992 (
            .O(N__15789),
            .I(N__15786));
    LocalMux I__2991 (
            .O(N__15786),
            .I(N__15783));
    Odrv12 I__2990 (
            .O(N__15783),
            .I(\receive_module.rx_counter.n4_adj_612 ));
    InMux I__2989 (
            .O(N__15780),
            .I(N__15777));
    LocalMux I__2988 (
            .O(N__15777),
            .I(N__15774));
    Odrv4 I__2987 (
            .O(N__15774),
            .I(\receive_module.rx_counter.n4 ));
    CascadeMux I__2986 (
            .O(N__15771),
            .I(\receive_module.rx_counter.n5_cascade_ ));
    InMux I__2985 (
            .O(N__15768),
            .I(N__15765));
    LocalMux I__2984 (
            .O(N__15765),
            .I(\receive_module.rx_counter.n3450 ));
    InMux I__2983 (
            .O(N__15762),
            .I(N__15758));
    InMux I__2982 (
            .O(N__15761),
            .I(N__15755));
    LocalMux I__2981 (
            .O(N__15758),
            .I(\receive_module.rx_counter.n3677 ));
    LocalMux I__2980 (
            .O(N__15755),
            .I(\receive_module.rx_counter.n3677 ));
    SRMux I__2979 (
            .O(N__15750),
            .I(N__15747));
    LocalMux I__2978 (
            .O(N__15747),
            .I(N__15743));
    SRMux I__2977 (
            .O(N__15746),
            .I(N__15740));
    Span4Mux_h I__2976 (
            .O(N__15743),
            .I(N__15737));
    LocalMux I__2975 (
            .O(N__15740),
            .I(N__15734));
    Odrv4 I__2974 (
            .O(N__15737),
            .I(\receive_module.rx_counter.n3 ));
    Odrv12 I__2973 (
            .O(N__15734),
            .I(\receive_module.rx_counter.n3 ));
    InMux I__2972 (
            .O(N__15729),
            .I(N__15725));
    InMux I__2971 (
            .O(N__15728),
            .I(N__15722));
    LocalMux I__2970 (
            .O(N__15725),
            .I(\receive_module.rx_counter.X_1 ));
    LocalMux I__2969 (
            .O(N__15722),
            .I(\receive_module.rx_counter.X_1 ));
    InMux I__2968 (
            .O(N__15717),
            .I(N__15713));
    InMux I__2967 (
            .O(N__15716),
            .I(N__15710));
    LocalMux I__2966 (
            .O(N__15713),
            .I(\receive_module.rx_counter.X_2 ));
    LocalMux I__2965 (
            .O(N__15710),
            .I(\receive_module.rx_counter.X_2 ));
    InMux I__2964 (
            .O(N__15705),
            .I(N__15701));
    InMux I__2963 (
            .O(N__15704),
            .I(N__15698));
    LocalMux I__2962 (
            .O(N__15701),
            .I(\receive_module.rx_counter.X_0 ));
    LocalMux I__2961 (
            .O(N__15698),
            .I(\receive_module.rx_counter.X_0 ));
    InMux I__2960 (
            .O(N__15693),
            .I(bfn_16_12_0_));
    InMux I__2959 (
            .O(N__15690),
            .I(\receive_module.rx_counter.n3202 ));
    InMux I__2958 (
            .O(N__15687),
            .I(\receive_module.rx_counter.n3203 ));
    InMux I__2957 (
            .O(N__15684),
            .I(\receive_module.rx_counter.n3204 ));
    InMux I__2956 (
            .O(N__15681),
            .I(N__15678));
    LocalMux I__2955 (
            .O(N__15678),
            .I(N__15675));
    Odrv4 I__2954 (
            .O(N__15675),
            .I(\tvp_video_buffer.BUFFER_0_5 ));
    CascadeMux I__2953 (
            .O(N__15672),
            .I(\receive_module.rx_counter.n3452_cascade_ ));
    InMux I__2952 (
            .O(N__15669),
            .I(N__15666));
    LocalMux I__2951 (
            .O(N__15666),
            .I(N__15663));
    Span4Mux_v I__2950 (
            .O(N__15663),
            .I(N__15660));
    Odrv4 I__2949 (
            .O(N__15660),
            .I(\tvp_video_buffer.BUFFER_1_5 ));
    InMux I__2948 (
            .O(N__15657),
            .I(N__15654));
    LocalMux I__2947 (
            .O(N__15654),
            .I(N__15650));
    InMux I__2946 (
            .O(N__15653),
            .I(N__15647));
    Span4Mux_s3_v I__2945 (
            .O(N__15650),
            .I(N__15644));
    LocalMux I__2944 (
            .O(N__15647),
            .I(N__15641));
    Span4Mux_v I__2943 (
            .O(N__15644),
            .I(N__15637));
    Span4Mux_v I__2942 (
            .O(N__15641),
            .I(N__15632));
    InMux I__2941 (
            .O(N__15640),
            .I(N__15628));
    Span4Mux_v I__2940 (
            .O(N__15637),
            .I(N__15625));
    InMux I__2939 (
            .O(N__15636),
            .I(N__15622));
    InMux I__2938 (
            .O(N__15635),
            .I(N__15619));
    Span4Mux_v I__2937 (
            .O(N__15632),
            .I(N__15616));
    InMux I__2936 (
            .O(N__15631),
            .I(N__15613));
    LocalMux I__2935 (
            .O(N__15628),
            .I(N__15610));
    Span4Mux_v I__2934 (
            .O(N__15625),
            .I(N__15605));
    LocalMux I__2933 (
            .O(N__15622),
            .I(N__15605));
    LocalMux I__2932 (
            .O(N__15619),
            .I(N__15602));
    Sp12to4 I__2931 (
            .O(N__15616),
            .I(N__15597));
    LocalMux I__2930 (
            .O(N__15613),
            .I(N__15597));
    Span4Mux_v I__2929 (
            .O(N__15610),
            .I(N__15594));
    Span4Mux_v I__2928 (
            .O(N__15605),
            .I(N__15590));
    Span4Mux_v I__2927 (
            .O(N__15602),
            .I(N__15587));
    Span12Mux_h I__2926 (
            .O(N__15597),
            .I(N__15583));
    Span4Mux_v I__2925 (
            .O(N__15594),
            .I(N__15580));
    InMux I__2924 (
            .O(N__15593),
            .I(N__15577));
    Span4Mux_v I__2923 (
            .O(N__15590),
            .I(N__15572));
    Span4Mux_v I__2922 (
            .O(N__15587),
            .I(N__15572));
    InMux I__2921 (
            .O(N__15586),
            .I(N__15569));
    Span12Mux_v I__2920 (
            .O(N__15583),
            .I(N__15562));
    Sp12to4 I__2919 (
            .O(N__15580),
            .I(N__15562));
    LocalMux I__2918 (
            .O(N__15577),
            .I(N__15562));
    Sp12to4 I__2917 (
            .O(N__15572),
            .I(N__15557));
    LocalMux I__2916 (
            .O(N__15569),
            .I(N__15557));
    Odrv12 I__2915 (
            .O(N__15562),
            .I(RX_DATA_3));
    Odrv12 I__2914 (
            .O(N__15557),
            .I(RX_DATA_3));
    InMux I__2913 (
            .O(N__15552),
            .I(N__15549));
    LocalMux I__2912 (
            .O(N__15549),
            .I(N__15546));
    Odrv4 I__2911 (
            .O(N__15546),
            .I(\receive_module.rx_counter.n10 ));
    CascadeMux I__2910 (
            .O(N__15543),
            .I(\receive_module.rx_counter.n14_cascade_ ));
    InMux I__2909 (
            .O(N__15540),
            .I(N__15537));
    LocalMux I__2908 (
            .O(N__15537),
            .I(N__15534));
    Span4Mux_h I__2907 (
            .O(N__15534),
            .I(N__15531));
    Odrv4 I__2906 (
            .O(N__15531),
            .I(RX_TX_SYNC));
    InMux I__2905 (
            .O(N__15528),
            .I(\receive_module.n3158 ));
    InMux I__2904 (
            .O(N__15525),
            .I(N__15521));
    InMux I__2903 (
            .O(N__15524),
            .I(N__15518));
    LocalMux I__2902 (
            .O(N__15521),
            .I(N__15515));
    LocalMux I__2901 (
            .O(N__15518),
            .I(N__15508));
    Span4Mux_v I__2900 (
            .O(N__15515),
            .I(N__15508));
    InMux I__2899 (
            .O(N__15514),
            .I(N__15505));
    InMux I__2898 (
            .O(N__15513),
            .I(N__15502));
    Odrv4 I__2897 (
            .O(N__15508),
            .I(\transmit_module.TX_ADDR_4 ));
    LocalMux I__2896 (
            .O(N__15505),
            .I(\transmit_module.TX_ADDR_4 ));
    LocalMux I__2895 (
            .O(N__15502),
            .I(\transmit_module.TX_ADDR_4 ));
    InMux I__2894 (
            .O(N__15495),
            .I(N__15492));
    LocalMux I__2893 (
            .O(N__15492),
            .I(\transmit_module.ADDR_Y_COMPONENT_4 ));
    InMux I__2892 (
            .O(N__15489),
            .I(N__15484));
    InMux I__2891 (
            .O(N__15488),
            .I(N__15481));
    InMux I__2890 (
            .O(N__15487),
            .I(N__15478));
    LocalMux I__2889 (
            .O(N__15484),
            .I(N__15474));
    LocalMux I__2888 (
            .O(N__15481),
            .I(N__15469));
    LocalMux I__2887 (
            .O(N__15478),
            .I(N__15469));
    CascadeMux I__2886 (
            .O(N__15477),
            .I(N__15466));
    Span4Mux_h I__2885 (
            .O(N__15474),
            .I(N__15463));
    Span4Mux_v I__2884 (
            .O(N__15469),
            .I(N__15460));
    InMux I__2883 (
            .O(N__15466),
            .I(N__15457));
    Odrv4 I__2882 (
            .O(N__15463),
            .I(\transmit_module.TX_ADDR_7 ));
    Odrv4 I__2881 (
            .O(N__15460),
            .I(\transmit_module.TX_ADDR_7 ));
    LocalMux I__2880 (
            .O(N__15457),
            .I(\transmit_module.TX_ADDR_7 ));
    InMux I__2879 (
            .O(N__15450),
            .I(N__15447));
    LocalMux I__2878 (
            .O(N__15447),
            .I(\transmit_module.ADDR_Y_COMPONENT_7 ));
    InMux I__2877 (
            .O(N__15444),
            .I(N__15440));
    InMux I__2876 (
            .O(N__15443),
            .I(N__15436));
    LocalMux I__2875 (
            .O(N__15440),
            .I(N__15433));
    CascadeMux I__2874 (
            .O(N__15439),
            .I(N__15429));
    LocalMux I__2873 (
            .O(N__15436),
            .I(N__15426));
    Span4Mux_v I__2872 (
            .O(N__15433),
            .I(N__15423));
    InMux I__2871 (
            .O(N__15432),
            .I(N__15420));
    InMux I__2870 (
            .O(N__15429),
            .I(N__15417));
    Odrv12 I__2869 (
            .O(N__15426),
            .I(\transmit_module.TX_ADDR_6 ));
    Odrv4 I__2868 (
            .O(N__15423),
            .I(\transmit_module.TX_ADDR_6 ));
    LocalMux I__2867 (
            .O(N__15420),
            .I(\transmit_module.TX_ADDR_6 ));
    LocalMux I__2866 (
            .O(N__15417),
            .I(\transmit_module.TX_ADDR_6 ));
    InMux I__2865 (
            .O(N__15408),
            .I(N__15405));
    LocalMux I__2864 (
            .O(N__15405),
            .I(\transmit_module.ADDR_Y_COMPONENT_6 ));
    CEMux I__2863 (
            .O(N__15402),
            .I(N__15398));
    CEMux I__2862 (
            .O(N__15401),
            .I(N__15394));
    LocalMux I__2861 (
            .O(N__15398),
            .I(N__15391));
    CEMux I__2860 (
            .O(N__15397),
            .I(N__15385));
    LocalMux I__2859 (
            .O(N__15394),
            .I(N__15382));
    Span4Mux_v I__2858 (
            .O(N__15391),
            .I(N__15379));
    CEMux I__2857 (
            .O(N__15390),
            .I(N__15376));
    CEMux I__2856 (
            .O(N__15389),
            .I(N__15373));
    CEMux I__2855 (
            .O(N__15388),
            .I(N__15370));
    LocalMux I__2854 (
            .O(N__15385),
            .I(N__15367));
    Span4Mux_v I__2853 (
            .O(N__15382),
            .I(N__15364));
    Span4Mux_h I__2852 (
            .O(N__15379),
            .I(N__15361));
    LocalMux I__2851 (
            .O(N__15376),
            .I(N__15358));
    LocalMux I__2850 (
            .O(N__15373),
            .I(N__15355));
    LocalMux I__2849 (
            .O(N__15370),
            .I(N__15350));
    Span4Mux_h I__2848 (
            .O(N__15367),
            .I(N__15350));
    Span4Mux_h I__2847 (
            .O(N__15364),
            .I(N__15345));
    Span4Mux_h I__2846 (
            .O(N__15361),
            .I(N__15345));
    Span4Mux_v I__2845 (
            .O(N__15358),
            .I(N__15342));
    Span4Mux_v I__2844 (
            .O(N__15355),
            .I(N__15339));
    Span4Mux_h I__2843 (
            .O(N__15350),
            .I(N__15336));
    Odrv4 I__2842 (
            .O(N__15345),
            .I(\transmit_module.n2310 ));
    Odrv4 I__2841 (
            .O(N__15342),
            .I(\transmit_module.n2310 ));
    Odrv4 I__2840 (
            .O(N__15339),
            .I(\transmit_module.n2310 ));
    Odrv4 I__2839 (
            .O(N__15336),
            .I(\transmit_module.n2310 ));
    InMux I__2838 (
            .O(N__15327),
            .I(N__15324));
    LocalMux I__2837 (
            .O(N__15324),
            .I(N__15321));
    Odrv12 I__2836 (
            .O(N__15321),
            .I(\receive_module.n136 ));
    CascadeMux I__2835 (
            .O(N__15318),
            .I(N__15314));
    CascadeMux I__2834 (
            .O(N__15317),
            .I(N__15311));
    CascadeBuf I__2833 (
            .O(N__15314),
            .I(N__15308));
    CascadeBuf I__2832 (
            .O(N__15311),
            .I(N__15305));
    CascadeMux I__2831 (
            .O(N__15308),
            .I(N__15302));
    CascadeMux I__2830 (
            .O(N__15305),
            .I(N__15299));
    CascadeBuf I__2829 (
            .O(N__15302),
            .I(N__15296));
    CascadeBuf I__2828 (
            .O(N__15299),
            .I(N__15293));
    CascadeMux I__2827 (
            .O(N__15296),
            .I(N__15290));
    CascadeMux I__2826 (
            .O(N__15293),
            .I(N__15287));
    CascadeBuf I__2825 (
            .O(N__15290),
            .I(N__15284));
    CascadeBuf I__2824 (
            .O(N__15287),
            .I(N__15281));
    CascadeMux I__2823 (
            .O(N__15284),
            .I(N__15278));
    CascadeMux I__2822 (
            .O(N__15281),
            .I(N__15275));
    CascadeBuf I__2821 (
            .O(N__15278),
            .I(N__15272));
    CascadeBuf I__2820 (
            .O(N__15275),
            .I(N__15269));
    CascadeMux I__2819 (
            .O(N__15272),
            .I(N__15266));
    CascadeMux I__2818 (
            .O(N__15269),
            .I(N__15263));
    CascadeBuf I__2817 (
            .O(N__15266),
            .I(N__15260));
    CascadeBuf I__2816 (
            .O(N__15263),
            .I(N__15257));
    CascadeMux I__2815 (
            .O(N__15260),
            .I(N__15254));
    CascadeMux I__2814 (
            .O(N__15257),
            .I(N__15251));
    CascadeBuf I__2813 (
            .O(N__15254),
            .I(N__15248));
    CascadeBuf I__2812 (
            .O(N__15251),
            .I(N__15245));
    CascadeMux I__2811 (
            .O(N__15248),
            .I(N__15242));
    CascadeMux I__2810 (
            .O(N__15245),
            .I(N__15239));
    CascadeBuf I__2809 (
            .O(N__15242),
            .I(N__15236));
    CascadeBuf I__2808 (
            .O(N__15239),
            .I(N__15233));
    CascadeMux I__2807 (
            .O(N__15236),
            .I(N__15230));
    CascadeMux I__2806 (
            .O(N__15233),
            .I(N__15227));
    CascadeBuf I__2805 (
            .O(N__15230),
            .I(N__15224));
    CascadeBuf I__2804 (
            .O(N__15227),
            .I(N__15221));
    CascadeMux I__2803 (
            .O(N__15224),
            .I(N__15218));
    CascadeMux I__2802 (
            .O(N__15221),
            .I(N__15215));
    CascadeBuf I__2801 (
            .O(N__15218),
            .I(N__15212));
    CascadeBuf I__2800 (
            .O(N__15215),
            .I(N__15209));
    CascadeMux I__2799 (
            .O(N__15212),
            .I(N__15206));
    CascadeMux I__2798 (
            .O(N__15209),
            .I(N__15203));
    CascadeBuf I__2797 (
            .O(N__15206),
            .I(N__15200));
    CascadeBuf I__2796 (
            .O(N__15203),
            .I(N__15197));
    CascadeMux I__2795 (
            .O(N__15200),
            .I(N__15194));
    CascadeMux I__2794 (
            .O(N__15197),
            .I(N__15191));
    CascadeBuf I__2793 (
            .O(N__15194),
            .I(N__15188));
    CascadeBuf I__2792 (
            .O(N__15191),
            .I(N__15185));
    CascadeMux I__2791 (
            .O(N__15188),
            .I(N__15182));
    CascadeMux I__2790 (
            .O(N__15185),
            .I(N__15179));
    CascadeBuf I__2789 (
            .O(N__15182),
            .I(N__15176));
    CascadeBuf I__2788 (
            .O(N__15179),
            .I(N__15173));
    CascadeMux I__2787 (
            .O(N__15176),
            .I(N__15170));
    CascadeMux I__2786 (
            .O(N__15173),
            .I(N__15167));
    CascadeBuf I__2785 (
            .O(N__15170),
            .I(N__15164));
    CascadeBuf I__2784 (
            .O(N__15167),
            .I(N__15161));
    CascadeMux I__2783 (
            .O(N__15164),
            .I(N__15158));
    CascadeMux I__2782 (
            .O(N__15161),
            .I(N__15155));
    CascadeBuf I__2781 (
            .O(N__15158),
            .I(N__15152));
    CascadeBuf I__2780 (
            .O(N__15155),
            .I(N__15149));
    CascadeMux I__2779 (
            .O(N__15152),
            .I(N__15146));
    CascadeMux I__2778 (
            .O(N__15149),
            .I(N__15143));
    CascadeBuf I__2777 (
            .O(N__15146),
            .I(N__15140));
    CascadeBuf I__2776 (
            .O(N__15143),
            .I(N__15137));
    CascadeMux I__2775 (
            .O(N__15140),
            .I(N__15134));
    CascadeMux I__2774 (
            .O(N__15137),
            .I(N__15131));
    InMux I__2773 (
            .O(N__15134),
            .I(N__15128));
    InMux I__2772 (
            .O(N__15131),
            .I(N__15125));
    LocalMux I__2771 (
            .O(N__15128),
            .I(N__15120));
    LocalMux I__2770 (
            .O(N__15125),
            .I(N__15117));
    CascadeMux I__2769 (
            .O(N__15124),
            .I(N__15114));
    InMux I__2768 (
            .O(N__15123),
            .I(N__15111));
    Span12Mux_h I__2767 (
            .O(N__15120),
            .I(N__15106));
    Span12Mux_h I__2766 (
            .O(N__15117),
            .I(N__15106));
    InMux I__2765 (
            .O(N__15114),
            .I(N__15103));
    LocalMux I__2764 (
            .O(N__15111),
            .I(N__15100));
    Span12Mux_v I__2763 (
            .O(N__15106),
            .I(N__15097));
    LocalMux I__2762 (
            .O(N__15103),
            .I(RX_ADDR_1));
    Odrv4 I__2761 (
            .O(N__15100),
            .I(RX_ADDR_1));
    Odrv12 I__2760 (
            .O(N__15097),
            .I(RX_ADDR_1));
    InMux I__2759 (
            .O(N__15090),
            .I(N__15087));
    LocalMux I__2758 (
            .O(N__15087),
            .I(N__15084));
    Odrv12 I__2757 (
            .O(N__15084),
            .I(\receive_module.n127 ));
    CascadeMux I__2756 (
            .O(N__15081),
            .I(N__15077));
    CascadeMux I__2755 (
            .O(N__15080),
            .I(N__15074));
    CascadeBuf I__2754 (
            .O(N__15077),
            .I(N__15071));
    CascadeBuf I__2753 (
            .O(N__15074),
            .I(N__15068));
    CascadeMux I__2752 (
            .O(N__15071),
            .I(N__15065));
    CascadeMux I__2751 (
            .O(N__15068),
            .I(N__15062));
    CascadeBuf I__2750 (
            .O(N__15065),
            .I(N__15059));
    CascadeBuf I__2749 (
            .O(N__15062),
            .I(N__15056));
    CascadeMux I__2748 (
            .O(N__15059),
            .I(N__15053));
    CascadeMux I__2747 (
            .O(N__15056),
            .I(N__15050));
    CascadeBuf I__2746 (
            .O(N__15053),
            .I(N__15047));
    CascadeBuf I__2745 (
            .O(N__15050),
            .I(N__15044));
    CascadeMux I__2744 (
            .O(N__15047),
            .I(N__15041));
    CascadeMux I__2743 (
            .O(N__15044),
            .I(N__15038));
    CascadeBuf I__2742 (
            .O(N__15041),
            .I(N__15035));
    CascadeBuf I__2741 (
            .O(N__15038),
            .I(N__15032));
    CascadeMux I__2740 (
            .O(N__15035),
            .I(N__15029));
    CascadeMux I__2739 (
            .O(N__15032),
            .I(N__15026));
    CascadeBuf I__2738 (
            .O(N__15029),
            .I(N__15023));
    CascadeBuf I__2737 (
            .O(N__15026),
            .I(N__15020));
    CascadeMux I__2736 (
            .O(N__15023),
            .I(N__15017));
    CascadeMux I__2735 (
            .O(N__15020),
            .I(N__15014));
    CascadeBuf I__2734 (
            .O(N__15017),
            .I(N__15011));
    CascadeBuf I__2733 (
            .O(N__15014),
            .I(N__15008));
    CascadeMux I__2732 (
            .O(N__15011),
            .I(N__15005));
    CascadeMux I__2731 (
            .O(N__15008),
            .I(N__15002));
    CascadeBuf I__2730 (
            .O(N__15005),
            .I(N__14999));
    CascadeBuf I__2729 (
            .O(N__15002),
            .I(N__14996));
    CascadeMux I__2728 (
            .O(N__14999),
            .I(N__14993));
    CascadeMux I__2727 (
            .O(N__14996),
            .I(N__14990));
    CascadeBuf I__2726 (
            .O(N__14993),
            .I(N__14987));
    CascadeBuf I__2725 (
            .O(N__14990),
            .I(N__14984));
    CascadeMux I__2724 (
            .O(N__14987),
            .I(N__14981));
    CascadeMux I__2723 (
            .O(N__14984),
            .I(N__14978));
    CascadeBuf I__2722 (
            .O(N__14981),
            .I(N__14975));
    CascadeBuf I__2721 (
            .O(N__14978),
            .I(N__14972));
    CascadeMux I__2720 (
            .O(N__14975),
            .I(N__14969));
    CascadeMux I__2719 (
            .O(N__14972),
            .I(N__14966));
    CascadeBuf I__2718 (
            .O(N__14969),
            .I(N__14963));
    CascadeBuf I__2717 (
            .O(N__14966),
            .I(N__14960));
    CascadeMux I__2716 (
            .O(N__14963),
            .I(N__14957));
    CascadeMux I__2715 (
            .O(N__14960),
            .I(N__14954));
    CascadeBuf I__2714 (
            .O(N__14957),
            .I(N__14951));
    CascadeBuf I__2713 (
            .O(N__14954),
            .I(N__14948));
    CascadeMux I__2712 (
            .O(N__14951),
            .I(N__14945));
    CascadeMux I__2711 (
            .O(N__14948),
            .I(N__14942));
    CascadeBuf I__2710 (
            .O(N__14945),
            .I(N__14939));
    CascadeBuf I__2709 (
            .O(N__14942),
            .I(N__14936));
    CascadeMux I__2708 (
            .O(N__14939),
            .I(N__14933));
    CascadeMux I__2707 (
            .O(N__14936),
            .I(N__14930));
    CascadeBuf I__2706 (
            .O(N__14933),
            .I(N__14927));
    CascadeBuf I__2705 (
            .O(N__14930),
            .I(N__14924));
    CascadeMux I__2704 (
            .O(N__14927),
            .I(N__14921));
    CascadeMux I__2703 (
            .O(N__14924),
            .I(N__14918));
    CascadeBuf I__2702 (
            .O(N__14921),
            .I(N__14915));
    CascadeBuf I__2701 (
            .O(N__14918),
            .I(N__14912));
    CascadeMux I__2700 (
            .O(N__14915),
            .I(N__14909));
    CascadeMux I__2699 (
            .O(N__14912),
            .I(N__14906));
    CascadeBuf I__2698 (
            .O(N__14909),
            .I(N__14903));
    CascadeBuf I__2697 (
            .O(N__14906),
            .I(N__14900));
    CascadeMux I__2696 (
            .O(N__14903),
            .I(N__14897));
    CascadeMux I__2695 (
            .O(N__14900),
            .I(N__14894));
    InMux I__2694 (
            .O(N__14897),
            .I(N__14891));
    InMux I__2693 (
            .O(N__14894),
            .I(N__14888));
    LocalMux I__2692 (
            .O(N__14891),
            .I(N__14885));
    LocalMux I__2691 (
            .O(N__14888),
            .I(N__14882));
    Span4Mux_s3_v I__2690 (
            .O(N__14885),
            .I(N__14877));
    Span4Mux_s3_v I__2689 (
            .O(N__14882),
            .I(N__14874));
    CascadeMux I__2688 (
            .O(N__14881),
            .I(N__14871));
    InMux I__2687 (
            .O(N__14880),
            .I(N__14868));
    Sp12to4 I__2686 (
            .O(N__14877),
            .I(N__14865));
    Sp12to4 I__2685 (
            .O(N__14874),
            .I(N__14862));
    InMux I__2684 (
            .O(N__14871),
            .I(N__14859));
    LocalMux I__2683 (
            .O(N__14868),
            .I(N__14856));
    Span12Mux_h I__2682 (
            .O(N__14865),
            .I(N__14851));
    Span12Mux_h I__2681 (
            .O(N__14862),
            .I(N__14851));
    LocalMux I__2680 (
            .O(N__14859),
            .I(RX_ADDR_10));
    Odrv4 I__2679 (
            .O(N__14856),
            .I(RX_ADDR_10));
    Odrv12 I__2678 (
            .O(N__14851),
            .I(RX_ADDR_10));
    InMux I__2677 (
            .O(N__14844),
            .I(N__14841));
    LocalMux I__2676 (
            .O(N__14841),
            .I(N__14838));
    Odrv12 I__2675 (
            .O(N__14838),
            .I(\receive_module.n137 ));
    CascadeMux I__2674 (
            .O(N__14835),
            .I(N__14831));
    CascadeMux I__2673 (
            .O(N__14834),
            .I(N__14828));
    CascadeBuf I__2672 (
            .O(N__14831),
            .I(N__14825));
    CascadeBuf I__2671 (
            .O(N__14828),
            .I(N__14822));
    CascadeMux I__2670 (
            .O(N__14825),
            .I(N__14819));
    CascadeMux I__2669 (
            .O(N__14822),
            .I(N__14816));
    CascadeBuf I__2668 (
            .O(N__14819),
            .I(N__14813));
    CascadeBuf I__2667 (
            .O(N__14816),
            .I(N__14810));
    CascadeMux I__2666 (
            .O(N__14813),
            .I(N__14807));
    CascadeMux I__2665 (
            .O(N__14810),
            .I(N__14804));
    CascadeBuf I__2664 (
            .O(N__14807),
            .I(N__14801));
    CascadeBuf I__2663 (
            .O(N__14804),
            .I(N__14798));
    CascadeMux I__2662 (
            .O(N__14801),
            .I(N__14795));
    CascadeMux I__2661 (
            .O(N__14798),
            .I(N__14792));
    CascadeBuf I__2660 (
            .O(N__14795),
            .I(N__14789));
    CascadeBuf I__2659 (
            .O(N__14792),
            .I(N__14786));
    CascadeMux I__2658 (
            .O(N__14789),
            .I(N__14783));
    CascadeMux I__2657 (
            .O(N__14786),
            .I(N__14780));
    CascadeBuf I__2656 (
            .O(N__14783),
            .I(N__14777));
    CascadeBuf I__2655 (
            .O(N__14780),
            .I(N__14774));
    CascadeMux I__2654 (
            .O(N__14777),
            .I(N__14771));
    CascadeMux I__2653 (
            .O(N__14774),
            .I(N__14768));
    CascadeBuf I__2652 (
            .O(N__14771),
            .I(N__14765));
    CascadeBuf I__2651 (
            .O(N__14768),
            .I(N__14762));
    CascadeMux I__2650 (
            .O(N__14765),
            .I(N__14759));
    CascadeMux I__2649 (
            .O(N__14762),
            .I(N__14756));
    CascadeBuf I__2648 (
            .O(N__14759),
            .I(N__14753));
    CascadeBuf I__2647 (
            .O(N__14756),
            .I(N__14750));
    CascadeMux I__2646 (
            .O(N__14753),
            .I(N__14747));
    CascadeMux I__2645 (
            .O(N__14750),
            .I(N__14744));
    CascadeBuf I__2644 (
            .O(N__14747),
            .I(N__14741));
    CascadeBuf I__2643 (
            .O(N__14744),
            .I(N__14738));
    CascadeMux I__2642 (
            .O(N__14741),
            .I(N__14735));
    CascadeMux I__2641 (
            .O(N__14738),
            .I(N__14732));
    CascadeBuf I__2640 (
            .O(N__14735),
            .I(N__14729));
    CascadeBuf I__2639 (
            .O(N__14732),
            .I(N__14726));
    CascadeMux I__2638 (
            .O(N__14729),
            .I(N__14723));
    CascadeMux I__2637 (
            .O(N__14726),
            .I(N__14720));
    CascadeBuf I__2636 (
            .O(N__14723),
            .I(N__14717));
    CascadeBuf I__2635 (
            .O(N__14720),
            .I(N__14714));
    CascadeMux I__2634 (
            .O(N__14717),
            .I(N__14711));
    CascadeMux I__2633 (
            .O(N__14714),
            .I(N__14708));
    CascadeBuf I__2632 (
            .O(N__14711),
            .I(N__14705));
    CascadeBuf I__2631 (
            .O(N__14708),
            .I(N__14702));
    CascadeMux I__2630 (
            .O(N__14705),
            .I(N__14699));
    CascadeMux I__2629 (
            .O(N__14702),
            .I(N__14696));
    CascadeBuf I__2628 (
            .O(N__14699),
            .I(N__14693));
    CascadeBuf I__2627 (
            .O(N__14696),
            .I(N__14690));
    CascadeMux I__2626 (
            .O(N__14693),
            .I(N__14687));
    CascadeMux I__2625 (
            .O(N__14690),
            .I(N__14684));
    CascadeBuf I__2624 (
            .O(N__14687),
            .I(N__14681));
    CascadeBuf I__2623 (
            .O(N__14684),
            .I(N__14678));
    CascadeMux I__2622 (
            .O(N__14681),
            .I(N__14675));
    CascadeMux I__2621 (
            .O(N__14678),
            .I(N__14672));
    CascadeBuf I__2620 (
            .O(N__14675),
            .I(N__14669));
    CascadeBuf I__2619 (
            .O(N__14672),
            .I(N__14666));
    CascadeMux I__2618 (
            .O(N__14669),
            .I(N__14663));
    CascadeMux I__2617 (
            .O(N__14666),
            .I(N__14660));
    CascadeBuf I__2616 (
            .O(N__14663),
            .I(N__14657));
    CascadeBuf I__2615 (
            .O(N__14660),
            .I(N__14654));
    CascadeMux I__2614 (
            .O(N__14657),
            .I(N__14651));
    CascadeMux I__2613 (
            .O(N__14654),
            .I(N__14648));
    InMux I__2612 (
            .O(N__14651),
            .I(N__14645));
    InMux I__2611 (
            .O(N__14648),
            .I(N__14642));
    LocalMux I__2610 (
            .O(N__14645),
            .I(N__14639));
    LocalMux I__2609 (
            .O(N__14642),
            .I(N__14634));
    Span4Mux_s2_v I__2608 (
            .O(N__14639),
            .I(N__14631));
    CascadeMux I__2607 (
            .O(N__14638),
            .I(N__14628));
    InMux I__2606 (
            .O(N__14637),
            .I(N__14625));
    Span12Mux_s1_v I__2605 (
            .O(N__14634),
            .I(N__14622));
    Sp12to4 I__2604 (
            .O(N__14631),
            .I(N__14619));
    InMux I__2603 (
            .O(N__14628),
            .I(N__14616));
    LocalMux I__2602 (
            .O(N__14625),
            .I(N__14613));
    Span12Mux_v I__2601 (
            .O(N__14622),
            .I(N__14610));
    Span12Mux_h I__2600 (
            .O(N__14619),
            .I(N__14607));
    LocalMux I__2599 (
            .O(N__14616),
            .I(RX_ADDR_0));
    Odrv4 I__2598 (
            .O(N__14613),
            .I(RX_ADDR_0));
    Odrv12 I__2597 (
            .O(N__14610),
            .I(RX_ADDR_0));
    Odrv12 I__2596 (
            .O(N__14607),
            .I(RX_ADDR_0));
    IoInMux I__2595 (
            .O(N__14598),
            .I(N__14594));
    IoInMux I__2594 (
            .O(N__14597),
            .I(N__14590));
    LocalMux I__2593 (
            .O(N__14594),
            .I(N__14587));
    IoInMux I__2592 (
            .O(N__14593),
            .I(N__14584));
    LocalMux I__2591 (
            .O(N__14590),
            .I(N__14581));
    Span4Mux_s1_h I__2590 (
            .O(N__14587),
            .I(N__14578));
    LocalMux I__2589 (
            .O(N__14584),
            .I(N__14575));
    Sp12to4 I__2588 (
            .O(N__14581),
            .I(N__14570));
    Sp12to4 I__2587 (
            .O(N__14578),
            .I(N__14570));
    IoSpan4Mux I__2586 (
            .O(N__14575),
            .I(N__14567));
    Span12Mux_v I__2585 (
            .O(N__14570),
            .I(N__14564));
    Sp12to4 I__2584 (
            .O(N__14567),
            .I(N__14561));
    Span12Mux_h I__2583 (
            .O(N__14564),
            .I(N__14556));
    Span12Mux_v I__2582 (
            .O(N__14561),
            .I(N__14556));
    Odrv12 I__2581 (
            .O(N__14556),
            .I(n1818));
    InMux I__2580 (
            .O(N__14553),
            .I(N__14550));
    LocalMux I__2579 (
            .O(N__14550),
            .I(N__14547));
    Span12Mux_s6_v I__2578 (
            .O(N__14547),
            .I(N__14544));
    Odrv12 I__2577 (
            .O(N__14544),
            .I(\receive_module.n135 ));
    CascadeMux I__2576 (
            .O(N__14541),
            .I(N__14538));
    CascadeBuf I__2575 (
            .O(N__14538),
            .I(N__14534));
    CascadeMux I__2574 (
            .O(N__14537),
            .I(N__14531));
    CascadeMux I__2573 (
            .O(N__14534),
            .I(N__14528));
    CascadeBuf I__2572 (
            .O(N__14531),
            .I(N__14525));
    CascadeBuf I__2571 (
            .O(N__14528),
            .I(N__14522));
    CascadeMux I__2570 (
            .O(N__14525),
            .I(N__14519));
    CascadeMux I__2569 (
            .O(N__14522),
            .I(N__14516));
    CascadeBuf I__2568 (
            .O(N__14519),
            .I(N__14513));
    CascadeBuf I__2567 (
            .O(N__14516),
            .I(N__14510));
    CascadeMux I__2566 (
            .O(N__14513),
            .I(N__14507));
    CascadeMux I__2565 (
            .O(N__14510),
            .I(N__14504));
    CascadeBuf I__2564 (
            .O(N__14507),
            .I(N__14501));
    CascadeBuf I__2563 (
            .O(N__14504),
            .I(N__14498));
    CascadeMux I__2562 (
            .O(N__14501),
            .I(N__14495));
    CascadeMux I__2561 (
            .O(N__14498),
            .I(N__14492));
    CascadeBuf I__2560 (
            .O(N__14495),
            .I(N__14489));
    CascadeBuf I__2559 (
            .O(N__14492),
            .I(N__14486));
    CascadeMux I__2558 (
            .O(N__14489),
            .I(N__14483));
    CascadeMux I__2557 (
            .O(N__14486),
            .I(N__14480));
    CascadeBuf I__2556 (
            .O(N__14483),
            .I(N__14477));
    CascadeBuf I__2555 (
            .O(N__14480),
            .I(N__14474));
    CascadeMux I__2554 (
            .O(N__14477),
            .I(N__14471));
    CascadeMux I__2553 (
            .O(N__14474),
            .I(N__14468));
    CascadeBuf I__2552 (
            .O(N__14471),
            .I(N__14465));
    CascadeBuf I__2551 (
            .O(N__14468),
            .I(N__14462));
    CascadeMux I__2550 (
            .O(N__14465),
            .I(N__14459));
    CascadeMux I__2549 (
            .O(N__14462),
            .I(N__14456));
    CascadeBuf I__2548 (
            .O(N__14459),
            .I(N__14453));
    CascadeBuf I__2547 (
            .O(N__14456),
            .I(N__14450));
    CascadeMux I__2546 (
            .O(N__14453),
            .I(N__14447));
    CascadeMux I__2545 (
            .O(N__14450),
            .I(N__14444));
    CascadeBuf I__2544 (
            .O(N__14447),
            .I(N__14441));
    CascadeBuf I__2543 (
            .O(N__14444),
            .I(N__14438));
    CascadeMux I__2542 (
            .O(N__14441),
            .I(N__14435));
    CascadeMux I__2541 (
            .O(N__14438),
            .I(N__14432));
    CascadeBuf I__2540 (
            .O(N__14435),
            .I(N__14429));
    CascadeBuf I__2539 (
            .O(N__14432),
            .I(N__14426));
    CascadeMux I__2538 (
            .O(N__14429),
            .I(N__14423));
    CascadeMux I__2537 (
            .O(N__14426),
            .I(N__14420));
    CascadeBuf I__2536 (
            .O(N__14423),
            .I(N__14417));
    CascadeBuf I__2535 (
            .O(N__14420),
            .I(N__14414));
    CascadeMux I__2534 (
            .O(N__14417),
            .I(N__14411));
    CascadeMux I__2533 (
            .O(N__14414),
            .I(N__14408));
    CascadeBuf I__2532 (
            .O(N__14411),
            .I(N__14405));
    CascadeBuf I__2531 (
            .O(N__14408),
            .I(N__14402));
    CascadeMux I__2530 (
            .O(N__14405),
            .I(N__14399));
    CascadeMux I__2529 (
            .O(N__14402),
            .I(N__14396));
    CascadeBuf I__2528 (
            .O(N__14399),
            .I(N__14393));
    CascadeBuf I__2527 (
            .O(N__14396),
            .I(N__14390));
    CascadeMux I__2526 (
            .O(N__14393),
            .I(N__14387));
    CascadeMux I__2525 (
            .O(N__14390),
            .I(N__14384));
    CascadeBuf I__2524 (
            .O(N__14387),
            .I(N__14381));
    CascadeBuf I__2523 (
            .O(N__14384),
            .I(N__14378));
    CascadeMux I__2522 (
            .O(N__14381),
            .I(N__14375));
    CascadeMux I__2521 (
            .O(N__14378),
            .I(N__14372));
    CascadeBuf I__2520 (
            .O(N__14375),
            .I(N__14369));
    CascadeBuf I__2519 (
            .O(N__14372),
            .I(N__14366));
    CascadeMux I__2518 (
            .O(N__14369),
            .I(N__14363));
    CascadeMux I__2517 (
            .O(N__14366),
            .I(N__14360));
    CascadeBuf I__2516 (
            .O(N__14363),
            .I(N__14357));
    InMux I__2515 (
            .O(N__14360),
            .I(N__14353));
    CascadeMux I__2514 (
            .O(N__14357),
            .I(N__14350));
    InMux I__2513 (
            .O(N__14356),
            .I(N__14347));
    LocalMux I__2512 (
            .O(N__14353),
            .I(N__14344));
    InMux I__2511 (
            .O(N__14350),
            .I(N__14341));
    LocalMux I__2510 (
            .O(N__14347),
            .I(N__14338));
    Span4Mux_s1_v I__2509 (
            .O(N__14344),
            .I(N__14335));
    LocalMux I__2508 (
            .O(N__14341),
            .I(N__14332));
    Span4Mux_v I__2507 (
            .O(N__14338),
            .I(N__14329));
    Span4Mux_h I__2506 (
            .O(N__14335),
            .I(N__14325));
    Span4Mux_s1_v I__2505 (
            .O(N__14332),
            .I(N__14322));
    Sp12to4 I__2504 (
            .O(N__14329),
            .I(N__14319));
    InMux I__2503 (
            .O(N__14328),
            .I(N__14316));
    Span4Mux_h I__2502 (
            .O(N__14325),
            .I(N__14313));
    Span4Mux_h I__2501 (
            .O(N__14322),
            .I(N__14310));
    Odrv12 I__2500 (
            .O(N__14319),
            .I(RX_ADDR_2));
    LocalMux I__2499 (
            .O(N__14316),
            .I(RX_ADDR_2));
    Odrv4 I__2498 (
            .O(N__14313),
            .I(RX_ADDR_2));
    Odrv4 I__2497 (
            .O(N__14310),
            .I(RX_ADDR_2));
    InMux I__2496 (
            .O(N__14301),
            .I(\receive_module.n3149 ));
    InMux I__2495 (
            .O(N__14298),
            .I(\receive_module.n3150 ));
    InMux I__2494 (
            .O(N__14295),
            .I(\receive_module.n3151 ));
    InMux I__2493 (
            .O(N__14292),
            .I(\receive_module.n3152 ));
    InMux I__2492 (
            .O(N__14289),
            .I(bfn_15_17_0_));
    InMux I__2491 (
            .O(N__14286),
            .I(\receive_module.n3154 ));
    InMux I__2490 (
            .O(N__14283),
            .I(\receive_module.n3155 ));
    InMux I__2489 (
            .O(N__14280),
            .I(\receive_module.n3156 ));
    InMux I__2488 (
            .O(N__14277),
            .I(\receive_module.n3157 ));
    InMux I__2487 (
            .O(N__14274),
            .I(N__14271));
    LocalMux I__2486 (
            .O(N__14271),
            .I(\transmit_module.n132 ));
    CascadeMux I__2485 (
            .O(N__14268),
            .I(\transmit_module.n147_cascade_ ));
    CascadeMux I__2484 (
            .O(N__14265),
            .I(N__14262));
    CascadeBuf I__2483 (
            .O(N__14262),
            .I(N__14259));
    CascadeMux I__2482 (
            .O(N__14259),
            .I(N__14255));
    CascadeMux I__2481 (
            .O(N__14258),
            .I(N__14252));
    CascadeBuf I__2480 (
            .O(N__14255),
            .I(N__14249));
    CascadeBuf I__2479 (
            .O(N__14252),
            .I(N__14246));
    CascadeMux I__2478 (
            .O(N__14249),
            .I(N__14243));
    CascadeMux I__2477 (
            .O(N__14246),
            .I(N__14240));
    CascadeBuf I__2476 (
            .O(N__14243),
            .I(N__14237));
    CascadeBuf I__2475 (
            .O(N__14240),
            .I(N__14234));
    CascadeMux I__2474 (
            .O(N__14237),
            .I(N__14231));
    CascadeMux I__2473 (
            .O(N__14234),
            .I(N__14228));
    CascadeBuf I__2472 (
            .O(N__14231),
            .I(N__14225));
    CascadeBuf I__2471 (
            .O(N__14228),
            .I(N__14222));
    CascadeMux I__2470 (
            .O(N__14225),
            .I(N__14219));
    CascadeMux I__2469 (
            .O(N__14222),
            .I(N__14216));
    CascadeBuf I__2468 (
            .O(N__14219),
            .I(N__14213));
    CascadeBuf I__2467 (
            .O(N__14216),
            .I(N__14210));
    CascadeMux I__2466 (
            .O(N__14213),
            .I(N__14207));
    CascadeMux I__2465 (
            .O(N__14210),
            .I(N__14204));
    CascadeBuf I__2464 (
            .O(N__14207),
            .I(N__14201));
    CascadeBuf I__2463 (
            .O(N__14204),
            .I(N__14198));
    CascadeMux I__2462 (
            .O(N__14201),
            .I(N__14195));
    CascadeMux I__2461 (
            .O(N__14198),
            .I(N__14192));
    CascadeBuf I__2460 (
            .O(N__14195),
            .I(N__14189));
    CascadeBuf I__2459 (
            .O(N__14192),
            .I(N__14186));
    CascadeMux I__2458 (
            .O(N__14189),
            .I(N__14183));
    CascadeMux I__2457 (
            .O(N__14186),
            .I(N__14180));
    CascadeBuf I__2456 (
            .O(N__14183),
            .I(N__14177));
    CascadeBuf I__2455 (
            .O(N__14180),
            .I(N__14174));
    CascadeMux I__2454 (
            .O(N__14177),
            .I(N__14171));
    CascadeMux I__2453 (
            .O(N__14174),
            .I(N__14168));
    CascadeBuf I__2452 (
            .O(N__14171),
            .I(N__14165));
    CascadeBuf I__2451 (
            .O(N__14168),
            .I(N__14162));
    CascadeMux I__2450 (
            .O(N__14165),
            .I(N__14159));
    CascadeMux I__2449 (
            .O(N__14162),
            .I(N__14156));
    CascadeBuf I__2448 (
            .O(N__14159),
            .I(N__14153));
    CascadeBuf I__2447 (
            .O(N__14156),
            .I(N__14150));
    CascadeMux I__2446 (
            .O(N__14153),
            .I(N__14147));
    CascadeMux I__2445 (
            .O(N__14150),
            .I(N__14144));
    CascadeBuf I__2444 (
            .O(N__14147),
            .I(N__14141));
    CascadeBuf I__2443 (
            .O(N__14144),
            .I(N__14138));
    CascadeMux I__2442 (
            .O(N__14141),
            .I(N__14135));
    CascadeMux I__2441 (
            .O(N__14138),
            .I(N__14132));
    CascadeBuf I__2440 (
            .O(N__14135),
            .I(N__14129));
    CascadeBuf I__2439 (
            .O(N__14132),
            .I(N__14126));
    CascadeMux I__2438 (
            .O(N__14129),
            .I(N__14123));
    CascadeMux I__2437 (
            .O(N__14126),
            .I(N__14120));
    CascadeBuf I__2436 (
            .O(N__14123),
            .I(N__14117));
    CascadeBuf I__2435 (
            .O(N__14120),
            .I(N__14114));
    CascadeMux I__2434 (
            .O(N__14117),
            .I(N__14111));
    CascadeMux I__2433 (
            .O(N__14114),
            .I(N__14108));
    CascadeBuf I__2432 (
            .O(N__14111),
            .I(N__14105));
    CascadeBuf I__2431 (
            .O(N__14108),
            .I(N__14102));
    CascadeMux I__2430 (
            .O(N__14105),
            .I(N__14099));
    CascadeMux I__2429 (
            .O(N__14102),
            .I(N__14096));
    CascadeBuf I__2428 (
            .O(N__14099),
            .I(N__14093));
    CascadeBuf I__2427 (
            .O(N__14096),
            .I(N__14090));
    CascadeMux I__2426 (
            .O(N__14093),
            .I(N__14087));
    CascadeMux I__2425 (
            .O(N__14090),
            .I(N__14084));
    InMux I__2424 (
            .O(N__14087),
            .I(N__14081));
    CascadeBuf I__2423 (
            .O(N__14084),
            .I(N__14078));
    LocalMux I__2422 (
            .O(N__14081),
            .I(N__14075));
    CascadeMux I__2421 (
            .O(N__14078),
            .I(N__14072));
    Span4Mux_s2_v I__2420 (
            .O(N__14075),
            .I(N__14069));
    InMux I__2419 (
            .O(N__14072),
            .I(N__14066));
    Span4Mux_v I__2418 (
            .O(N__14069),
            .I(N__14063));
    LocalMux I__2417 (
            .O(N__14066),
            .I(N__14060));
    Sp12to4 I__2416 (
            .O(N__14063),
            .I(N__14057));
    Span12Mux_s5_v I__2415 (
            .O(N__14060),
            .I(N__14054));
    Span12Mux_h I__2414 (
            .O(N__14057),
            .I(N__14051));
    Span12Mux_v I__2413 (
            .O(N__14054),
            .I(N__14048));
    Odrv12 I__2412 (
            .O(N__14051),
            .I(n28));
    Odrv12 I__2411 (
            .O(N__14048),
            .I(n28));
    InMux I__2410 (
            .O(N__14043),
            .I(N__14036));
    InMux I__2409 (
            .O(N__14042),
            .I(N__14033));
    InMux I__2408 (
            .O(N__14041),
            .I(N__14030));
    InMux I__2407 (
            .O(N__14040),
            .I(N__14021));
    InMux I__2406 (
            .O(N__14039),
            .I(N__14018));
    LocalMux I__2405 (
            .O(N__14036),
            .I(N__14011));
    LocalMux I__2404 (
            .O(N__14033),
            .I(N__14011));
    LocalMux I__2403 (
            .O(N__14030),
            .I(N__14011));
    InMux I__2402 (
            .O(N__14029),
            .I(N__14006));
    InMux I__2401 (
            .O(N__14028),
            .I(N__14006));
    InMux I__2400 (
            .O(N__14027),
            .I(N__14003));
    InMux I__2399 (
            .O(N__14026),
            .I(N__13995));
    InMux I__2398 (
            .O(N__14025),
            .I(N__13995));
    InMux I__2397 (
            .O(N__14024),
            .I(N__13992));
    LocalMux I__2396 (
            .O(N__14021),
            .I(N__13987));
    LocalMux I__2395 (
            .O(N__14018),
            .I(N__13987));
    Span4Mux_v I__2394 (
            .O(N__14011),
            .I(N__13980));
    LocalMux I__2393 (
            .O(N__14006),
            .I(N__13980));
    LocalMux I__2392 (
            .O(N__14003),
            .I(N__13980));
    InMux I__2391 (
            .O(N__14002),
            .I(N__13973));
    InMux I__2390 (
            .O(N__14001),
            .I(N__13973));
    InMux I__2389 (
            .O(N__14000),
            .I(N__13973));
    LocalMux I__2388 (
            .O(N__13995),
            .I(\transmit_module.VGA_VISIBLE ));
    LocalMux I__2387 (
            .O(N__13992),
            .I(\transmit_module.VGA_VISIBLE ));
    Odrv12 I__2386 (
            .O(N__13987),
            .I(\transmit_module.VGA_VISIBLE ));
    Odrv4 I__2385 (
            .O(N__13980),
            .I(\transmit_module.VGA_VISIBLE ));
    LocalMux I__2384 (
            .O(N__13973),
            .I(\transmit_module.VGA_VISIBLE ));
    InMux I__2383 (
            .O(N__13962),
            .I(N__13959));
    LocalMux I__2382 (
            .O(N__13959),
            .I(\transmit_module.n128 ));
    InMux I__2381 (
            .O(N__13956),
            .I(N__13953));
    LocalMux I__2380 (
            .O(N__13953),
            .I(N__13950));
    Span4Mux_v I__2379 (
            .O(N__13950),
            .I(N__13947));
    Odrv4 I__2378 (
            .O(N__13947),
            .I(\transmit_module.n143 ));
    InMux I__2377 (
            .O(N__13944),
            .I(N__13941));
    LocalMux I__2376 (
            .O(N__13941),
            .I(N__13938));
    Span4Mux_h I__2375 (
            .O(N__13938),
            .I(N__13935));
    Odrv4 I__2374 (
            .O(N__13935),
            .I(\transmit_module.n112 ));
    CascadeMux I__2373 (
            .O(N__13932),
            .I(\transmit_module.n143_cascade_ ));
    InMux I__2372 (
            .O(N__13929),
            .I(N__13923));
    InMux I__2371 (
            .O(N__13928),
            .I(N__13923));
    LocalMux I__2370 (
            .O(N__13923),
            .I(\transmit_module.n116 ));
    InMux I__2369 (
            .O(N__13920),
            .I(N__13917));
    LocalMux I__2368 (
            .O(N__13917),
            .I(\transmit_module.n147 ));
    InMux I__2367 (
            .O(N__13914),
            .I(N__13910));
    CascadeMux I__2366 (
            .O(N__13913),
            .I(N__13905));
    LocalMux I__2365 (
            .O(N__13910),
            .I(N__13902));
    InMux I__2364 (
            .O(N__13909),
            .I(N__13899));
    InMux I__2363 (
            .O(N__13908),
            .I(N__13896));
    InMux I__2362 (
            .O(N__13905),
            .I(N__13893));
    Odrv4 I__2361 (
            .O(N__13902),
            .I(\transmit_module.TX_ADDR_0 ));
    LocalMux I__2360 (
            .O(N__13899),
            .I(\transmit_module.TX_ADDR_0 ));
    LocalMux I__2359 (
            .O(N__13896),
            .I(\transmit_module.TX_ADDR_0 ));
    LocalMux I__2358 (
            .O(N__13893),
            .I(\transmit_module.TX_ADDR_0 ));
    InMux I__2357 (
            .O(N__13884),
            .I(bfn_15_16_0_));
    InMux I__2356 (
            .O(N__13881),
            .I(\receive_module.n3146 ));
    InMux I__2355 (
            .O(N__13878),
            .I(\receive_module.n3147 ));
    InMux I__2354 (
            .O(N__13875),
            .I(\receive_module.n3148 ));
    InMux I__2353 (
            .O(N__13872),
            .I(N__13869));
    LocalMux I__2352 (
            .O(N__13869),
            .I(\transmit_module.X_DELTA_PATTERN_8 ));
    InMux I__2351 (
            .O(N__13866),
            .I(N__13863));
    LocalMux I__2350 (
            .O(N__13863),
            .I(N__13860));
    Span4Mux_v I__2349 (
            .O(N__13860),
            .I(N__13857));
    Odrv4 I__2348 (
            .O(N__13857),
            .I(\transmit_module.X_DELTA_PATTERN_7 ));
    InMux I__2347 (
            .O(N__13854),
            .I(N__13851));
    LocalMux I__2346 (
            .O(N__13851),
            .I(N__13848));
    Odrv4 I__2345 (
            .O(N__13848),
            .I(\transmit_module.X_DELTA_PATTERN_3 ));
    InMux I__2344 (
            .O(N__13845),
            .I(N__13842));
    LocalMux I__2343 (
            .O(N__13842),
            .I(\transmit_module.X_DELTA_PATTERN_9 ));
    InMux I__2342 (
            .O(N__13839),
            .I(N__13836));
    LocalMux I__2341 (
            .O(N__13836),
            .I(\transmit_module.X_DELTA_PATTERN_10 ));
    InMux I__2340 (
            .O(N__13833),
            .I(N__13830));
    LocalMux I__2339 (
            .O(N__13830),
            .I(N__13827));
    Span4Mux_v I__2338 (
            .O(N__13827),
            .I(N__13824));
    Odrv4 I__2337 (
            .O(N__13824),
            .I(\transmit_module.X_DELTA_PATTERN_12 ));
    InMux I__2336 (
            .O(N__13821),
            .I(N__13818));
    LocalMux I__2335 (
            .O(N__13818),
            .I(\transmit_module.X_DELTA_PATTERN_11 ));
    InMux I__2334 (
            .O(N__13815),
            .I(N__13812));
    LocalMux I__2333 (
            .O(N__13812),
            .I(\transmit_module.X_DELTA_PATTERN_2 ));
    InMux I__2332 (
            .O(N__13809),
            .I(N__13806));
    LocalMux I__2331 (
            .O(N__13806),
            .I(\transmit_module.X_DELTA_PATTERN_1 ));
    InMux I__2330 (
            .O(N__13803),
            .I(N__13800));
    LocalMux I__2329 (
            .O(N__13800),
            .I(\transmit_module.n126 ));
    InMux I__2328 (
            .O(N__13797),
            .I(N__13794));
    LocalMux I__2327 (
            .O(N__13794),
            .I(N__13791));
    Span4Mux_v I__2326 (
            .O(N__13791),
            .I(N__13788));
    Odrv4 I__2325 (
            .O(N__13788),
            .I(\transmit_module.n141 ));
    CascadeMux I__2324 (
            .O(N__13785),
            .I(\transmit_module.n141_cascade_ ));
    InMux I__2323 (
            .O(N__13782),
            .I(N__13779));
    LocalMux I__2322 (
            .O(N__13779),
            .I(N__13775));
    InMux I__2321 (
            .O(N__13778),
            .I(N__13772));
    Odrv4 I__2320 (
            .O(N__13775),
            .I(\transmit_module.n110 ));
    LocalMux I__2319 (
            .O(N__13772),
            .I(\transmit_module.n110 ));
    InMux I__2318 (
            .O(N__13767),
            .I(N__13764));
    LocalMux I__2317 (
            .O(N__13764),
            .I(N__13761));
    Odrv12 I__2316 (
            .O(N__13761),
            .I(\tvp_vs_buffer.BUFFER_2_0 ));
    InMux I__2315 (
            .O(N__13758),
            .I(N__13754));
    InMux I__2314 (
            .O(N__13757),
            .I(N__13750));
    LocalMux I__2313 (
            .O(N__13754),
            .I(N__13747));
    InMux I__2312 (
            .O(N__13753),
            .I(N__13744));
    LocalMux I__2311 (
            .O(N__13750),
            .I(\transmit_module.video_signal_controller.VGA_Y_11 ));
    Odrv4 I__2310 (
            .O(N__13747),
            .I(\transmit_module.video_signal_controller.VGA_Y_11 ));
    LocalMux I__2309 (
            .O(N__13744),
            .I(\transmit_module.video_signal_controller.VGA_Y_11 ));
    InMux I__2308 (
            .O(N__13737),
            .I(N__13733));
    InMux I__2307 (
            .O(N__13736),
            .I(N__13730));
    LocalMux I__2306 (
            .O(N__13733),
            .I(N__13724));
    LocalMux I__2305 (
            .O(N__13730),
            .I(N__13724));
    InMux I__2304 (
            .O(N__13729),
            .I(N__13721));
    Odrv4 I__2303 (
            .O(N__13724),
            .I(\transmit_module.video_signal_controller.VGA_Y_10 ));
    LocalMux I__2302 (
            .O(N__13721),
            .I(\transmit_module.video_signal_controller.VGA_Y_10 ));
    InMux I__2301 (
            .O(N__13716),
            .I(N__13713));
    LocalMux I__2300 (
            .O(N__13713),
            .I(\transmit_module.video_signal_controller.n3461 ));
    InMux I__2299 (
            .O(N__13710),
            .I(N__13706));
    InMux I__2298 (
            .O(N__13709),
            .I(N__13703));
    LocalMux I__2297 (
            .O(N__13706),
            .I(\transmit_module.video_signal_controller.n3375 ));
    LocalMux I__2296 (
            .O(N__13703),
            .I(\transmit_module.video_signal_controller.n3375 ));
    CascadeMux I__2295 (
            .O(N__13698),
            .I(\transmit_module.video_signal_controller.n3673_cascade_ ));
    InMux I__2294 (
            .O(N__13695),
            .I(N__13691));
    InMux I__2293 (
            .O(N__13694),
            .I(N__13687));
    LocalMux I__2292 (
            .O(N__13691),
            .I(N__13684));
    InMux I__2291 (
            .O(N__13690),
            .I(N__13681));
    LocalMux I__2290 (
            .O(N__13687),
            .I(\transmit_module.video_signal_controller.VGA_Y_9 ));
    Odrv4 I__2289 (
            .O(N__13684),
            .I(\transmit_module.video_signal_controller.VGA_Y_9 ));
    LocalMux I__2288 (
            .O(N__13681),
            .I(\transmit_module.video_signal_controller.VGA_Y_9 ));
    InMux I__2287 (
            .O(N__13674),
            .I(N__13670));
    InMux I__2286 (
            .O(N__13673),
            .I(N__13667));
    LocalMux I__2285 (
            .O(N__13670),
            .I(\transmit_module.video_signal_controller.n3379 ));
    LocalMux I__2284 (
            .O(N__13667),
            .I(\transmit_module.video_signal_controller.n3379 ));
    InMux I__2283 (
            .O(N__13662),
            .I(\receive_module.rx_counter.n3207 ));
    InMux I__2282 (
            .O(N__13659),
            .I(\receive_module.rx_counter.n3208 ));
    InMux I__2281 (
            .O(N__13656),
            .I(\receive_module.rx_counter.n3209 ));
    InMux I__2280 (
            .O(N__13653),
            .I(\receive_module.rx_counter.n3210 ));
    InMux I__2279 (
            .O(N__13650),
            .I(\receive_module.rx_counter.n3211 ));
    InMux I__2278 (
            .O(N__13647),
            .I(\receive_module.rx_counter.n3212 ));
    InMux I__2277 (
            .O(N__13644),
            .I(\receive_module.rx_counter.n3213 ));
    InMux I__2276 (
            .O(N__13641),
            .I(bfn_15_11_0_));
    InMux I__2275 (
            .O(N__13638),
            .I(\receive_module.rx_counter.n3215 ));
    InMux I__2274 (
            .O(N__13635),
            .I(N__13632));
    LocalMux I__2273 (
            .O(N__13632),
            .I(N__13629));
    Span4Mux_h I__2272 (
            .O(N__13629),
            .I(N__13626));
    Odrv4 I__2271 (
            .O(N__13626),
            .I(TVP_VIDEO_c_5));
    IoInMux I__2270 (
            .O(N__13623),
            .I(N__13620));
    LocalMux I__2269 (
            .O(N__13620),
            .I(N__13617));
    IoSpan4Mux I__2268 (
            .O(N__13617),
            .I(N__13614));
    Span4Mux_s1_h I__2267 (
            .O(N__13614),
            .I(N__13611));
    Sp12to4 I__2266 (
            .O(N__13611),
            .I(N__13607));
    InMux I__2265 (
            .O(N__13610),
            .I(N__13604));
    Span12Mux_h I__2264 (
            .O(N__13607),
            .I(N__13601));
    LocalMux I__2263 (
            .O(N__13604),
            .I(N__13598));
    Odrv12 I__2262 (
            .O(N__13601),
            .I(DEBUG_c_1_c));
    Odrv12 I__2261 (
            .O(N__13598),
            .I(DEBUG_c_1_c));
    InMux I__2260 (
            .O(N__13593),
            .I(N__13590));
    LocalMux I__2259 (
            .O(N__13590),
            .I(\tvp_vs_buffer.BUFFER_0_0 ));
    InMux I__2258 (
            .O(N__13587),
            .I(N__13584));
    LocalMux I__2257 (
            .O(N__13584),
            .I(\tvp_vs_buffer.BUFFER_1_0 ));
    InMux I__2256 (
            .O(N__13581),
            .I(N__13577));
    InMux I__2255 (
            .O(N__13580),
            .I(N__13574));
    LocalMux I__2254 (
            .O(N__13577),
            .I(N__13567));
    LocalMux I__2253 (
            .O(N__13574),
            .I(N__13564));
    InMux I__2252 (
            .O(N__13573),
            .I(N__13561));
    InMux I__2251 (
            .O(N__13572),
            .I(N__13558));
    InMux I__2250 (
            .O(N__13571),
            .I(N__13555));
    InMux I__2249 (
            .O(N__13570),
            .I(N__13550));
    Span12Mux_s8_h I__2248 (
            .O(N__13567),
            .I(N__13546));
    Span12Mux_s7_v I__2247 (
            .O(N__13564),
            .I(N__13541));
    LocalMux I__2246 (
            .O(N__13561),
            .I(N__13541));
    LocalMux I__2245 (
            .O(N__13558),
            .I(N__13536));
    LocalMux I__2244 (
            .O(N__13555),
            .I(N__13536));
    InMux I__2243 (
            .O(N__13554),
            .I(N__13533));
    InMux I__2242 (
            .O(N__13553),
            .I(N__13530));
    LocalMux I__2241 (
            .O(N__13550),
            .I(N__13527));
    InMux I__2240 (
            .O(N__13549),
            .I(N__13524));
    Span12Mux_v I__2239 (
            .O(N__13546),
            .I(N__13521));
    Span12Mux_v I__2238 (
            .O(N__13541),
            .I(N__13518));
    Span12Mux_v I__2237 (
            .O(N__13536),
            .I(N__13515));
    LocalMux I__2236 (
            .O(N__13533),
            .I(N__13512));
    LocalMux I__2235 (
            .O(N__13530),
            .I(N__13509));
    Span4Mux_h I__2234 (
            .O(N__13527),
            .I(N__13506));
    LocalMux I__2233 (
            .O(N__13524),
            .I(N__13503));
    Span12Mux_v I__2232 (
            .O(N__13521),
            .I(N__13500));
    Span12Mux_h I__2231 (
            .O(N__13518),
            .I(N__13491));
    Span12Mux_h I__2230 (
            .O(N__13515),
            .I(N__13491));
    Span12Mux_h I__2229 (
            .O(N__13512),
            .I(N__13491));
    Span12Mux_h I__2228 (
            .O(N__13509),
            .I(N__13491));
    Span4Mux_h I__2227 (
            .O(N__13506),
            .I(N__13488));
    Span4Mux_v I__2226 (
            .O(N__13503),
            .I(N__13485));
    Odrv12 I__2225 (
            .O(N__13500),
            .I(RX_DATA_5));
    Odrv12 I__2224 (
            .O(N__13491),
            .I(RX_DATA_5));
    Odrv4 I__2223 (
            .O(N__13488),
            .I(RX_DATA_5));
    Odrv4 I__2222 (
            .O(N__13485),
            .I(RX_DATA_5));
    CascadeMux I__2221 (
            .O(N__13476),
            .I(\receive_module.sync_wd.n6_cascade_ ));
    CascadeMux I__2220 (
            .O(N__13473),
            .I(\receive_module.sync_wd.n4_cascade_ ));
    InMux I__2219 (
            .O(N__13470),
            .I(N__13467));
    LocalMux I__2218 (
            .O(N__13467),
            .I(\receive_module.sync_wd.old_visible ));
    InMux I__2217 (
            .O(N__13464),
            .I(bfn_15_10_0_));
    CascadeMux I__2216 (
            .O(N__13461),
            .I(N__13457));
    CascadeMux I__2215 (
            .O(N__13460),
            .I(N__13454));
    CascadeBuf I__2214 (
            .O(N__13457),
            .I(N__13451));
    CascadeBuf I__2213 (
            .O(N__13454),
            .I(N__13448));
    CascadeMux I__2212 (
            .O(N__13451),
            .I(N__13445));
    CascadeMux I__2211 (
            .O(N__13448),
            .I(N__13442));
    CascadeBuf I__2210 (
            .O(N__13445),
            .I(N__13439));
    CascadeBuf I__2209 (
            .O(N__13442),
            .I(N__13436));
    CascadeMux I__2208 (
            .O(N__13439),
            .I(N__13433));
    CascadeMux I__2207 (
            .O(N__13436),
            .I(N__13430));
    CascadeBuf I__2206 (
            .O(N__13433),
            .I(N__13427));
    CascadeBuf I__2205 (
            .O(N__13430),
            .I(N__13424));
    CascadeMux I__2204 (
            .O(N__13427),
            .I(N__13421));
    CascadeMux I__2203 (
            .O(N__13424),
            .I(N__13418));
    CascadeBuf I__2202 (
            .O(N__13421),
            .I(N__13415));
    CascadeBuf I__2201 (
            .O(N__13418),
            .I(N__13412));
    CascadeMux I__2200 (
            .O(N__13415),
            .I(N__13409));
    CascadeMux I__2199 (
            .O(N__13412),
            .I(N__13406));
    CascadeBuf I__2198 (
            .O(N__13409),
            .I(N__13403));
    CascadeBuf I__2197 (
            .O(N__13406),
            .I(N__13400));
    CascadeMux I__2196 (
            .O(N__13403),
            .I(N__13397));
    CascadeMux I__2195 (
            .O(N__13400),
            .I(N__13394));
    CascadeBuf I__2194 (
            .O(N__13397),
            .I(N__13391));
    CascadeBuf I__2193 (
            .O(N__13394),
            .I(N__13388));
    CascadeMux I__2192 (
            .O(N__13391),
            .I(N__13385));
    CascadeMux I__2191 (
            .O(N__13388),
            .I(N__13382));
    CascadeBuf I__2190 (
            .O(N__13385),
            .I(N__13379));
    CascadeBuf I__2189 (
            .O(N__13382),
            .I(N__13376));
    CascadeMux I__2188 (
            .O(N__13379),
            .I(N__13373));
    CascadeMux I__2187 (
            .O(N__13376),
            .I(N__13370));
    CascadeBuf I__2186 (
            .O(N__13373),
            .I(N__13367));
    CascadeBuf I__2185 (
            .O(N__13370),
            .I(N__13364));
    CascadeMux I__2184 (
            .O(N__13367),
            .I(N__13361));
    CascadeMux I__2183 (
            .O(N__13364),
            .I(N__13358));
    CascadeBuf I__2182 (
            .O(N__13361),
            .I(N__13355));
    CascadeBuf I__2181 (
            .O(N__13358),
            .I(N__13352));
    CascadeMux I__2180 (
            .O(N__13355),
            .I(N__13349));
    CascadeMux I__2179 (
            .O(N__13352),
            .I(N__13346));
    CascadeBuf I__2178 (
            .O(N__13349),
            .I(N__13343));
    CascadeBuf I__2177 (
            .O(N__13346),
            .I(N__13340));
    CascadeMux I__2176 (
            .O(N__13343),
            .I(N__13337));
    CascadeMux I__2175 (
            .O(N__13340),
            .I(N__13334));
    CascadeBuf I__2174 (
            .O(N__13337),
            .I(N__13331));
    CascadeBuf I__2173 (
            .O(N__13334),
            .I(N__13328));
    CascadeMux I__2172 (
            .O(N__13331),
            .I(N__13325));
    CascadeMux I__2171 (
            .O(N__13328),
            .I(N__13322));
    CascadeBuf I__2170 (
            .O(N__13325),
            .I(N__13319));
    CascadeBuf I__2169 (
            .O(N__13322),
            .I(N__13316));
    CascadeMux I__2168 (
            .O(N__13319),
            .I(N__13313));
    CascadeMux I__2167 (
            .O(N__13316),
            .I(N__13310));
    CascadeBuf I__2166 (
            .O(N__13313),
            .I(N__13307));
    CascadeBuf I__2165 (
            .O(N__13310),
            .I(N__13304));
    CascadeMux I__2164 (
            .O(N__13307),
            .I(N__13301));
    CascadeMux I__2163 (
            .O(N__13304),
            .I(N__13298));
    CascadeBuf I__2162 (
            .O(N__13301),
            .I(N__13295));
    CascadeBuf I__2161 (
            .O(N__13298),
            .I(N__13292));
    CascadeMux I__2160 (
            .O(N__13295),
            .I(N__13289));
    CascadeMux I__2159 (
            .O(N__13292),
            .I(N__13286));
    CascadeBuf I__2158 (
            .O(N__13289),
            .I(N__13283));
    CascadeBuf I__2157 (
            .O(N__13286),
            .I(N__13280));
    CascadeMux I__2156 (
            .O(N__13283),
            .I(N__13277));
    CascadeMux I__2155 (
            .O(N__13280),
            .I(N__13274));
    InMux I__2154 (
            .O(N__13277),
            .I(N__13271));
    InMux I__2153 (
            .O(N__13274),
            .I(N__13268));
    LocalMux I__2152 (
            .O(N__13271),
            .I(N__13265));
    LocalMux I__2151 (
            .O(N__13268),
            .I(N__13262));
    Sp12to4 I__2150 (
            .O(N__13265),
            .I(N__13259));
    Span12Mux_s9_h I__2149 (
            .O(N__13262),
            .I(N__13256));
    Span12Mux_s5_v I__2148 (
            .O(N__13259),
            .I(N__13253));
    Span12Mux_v I__2147 (
            .O(N__13256),
            .I(N__13250));
    Span12Mux_h I__2146 (
            .O(N__13253),
            .I(N__13247));
    Odrv12 I__2145 (
            .O(N__13250),
            .I(n22));
    Odrv12 I__2144 (
            .O(N__13247),
            .I(n22));
    CascadeMux I__2143 (
            .O(N__13242),
            .I(\transmit_module.n112_cascade_ ));
    CascadeMux I__2142 (
            .O(N__13239),
            .I(N__13236));
    CascadeBuf I__2141 (
            .O(N__13236),
            .I(N__13232));
    CascadeMux I__2140 (
            .O(N__13235),
            .I(N__13229));
    CascadeMux I__2139 (
            .O(N__13232),
            .I(N__13226));
    CascadeBuf I__2138 (
            .O(N__13229),
            .I(N__13223));
    CascadeBuf I__2137 (
            .O(N__13226),
            .I(N__13220));
    CascadeMux I__2136 (
            .O(N__13223),
            .I(N__13217));
    CascadeMux I__2135 (
            .O(N__13220),
            .I(N__13214));
    CascadeBuf I__2134 (
            .O(N__13217),
            .I(N__13211));
    CascadeBuf I__2133 (
            .O(N__13214),
            .I(N__13208));
    CascadeMux I__2132 (
            .O(N__13211),
            .I(N__13205));
    CascadeMux I__2131 (
            .O(N__13208),
            .I(N__13202));
    CascadeBuf I__2130 (
            .O(N__13205),
            .I(N__13199));
    CascadeBuf I__2129 (
            .O(N__13202),
            .I(N__13196));
    CascadeMux I__2128 (
            .O(N__13199),
            .I(N__13193));
    CascadeMux I__2127 (
            .O(N__13196),
            .I(N__13190));
    CascadeBuf I__2126 (
            .O(N__13193),
            .I(N__13187));
    CascadeBuf I__2125 (
            .O(N__13190),
            .I(N__13184));
    CascadeMux I__2124 (
            .O(N__13187),
            .I(N__13181));
    CascadeMux I__2123 (
            .O(N__13184),
            .I(N__13178));
    CascadeBuf I__2122 (
            .O(N__13181),
            .I(N__13175));
    CascadeBuf I__2121 (
            .O(N__13178),
            .I(N__13172));
    CascadeMux I__2120 (
            .O(N__13175),
            .I(N__13169));
    CascadeMux I__2119 (
            .O(N__13172),
            .I(N__13166));
    CascadeBuf I__2118 (
            .O(N__13169),
            .I(N__13163));
    CascadeBuf I__2117 (
            .O(N__13166),
            .I(N__13160));
    CascadeMux I__2116 (
            .O(N__13163),
            .I(N__13157));
    CascadeMux I__2115 (
            .O(N__13160),
            .I(N__13154));
    CascadeBuf I__2114 (
            .O(N__13157),
            .I(N__13151));
    CascadeBuf I__2113 (
            .O(N__13154),
            .I(N__13148));
    CascadeMux I__2112 (
            .O(N__13151),
            .I(N__13145));
    CascadeMux I__2111 (
            .O(N__13148),
            .I(N__13142));
    CascadeBuf I__2110 (
            .O(N__13145),
            .I(N__13139));
    CascadeBuf I__2109 (
            .O(N__13142),
            .I(N__13136));
    CascadeMux I__2108 (
            .O(N__13139),
            .I(N__13133));
    CascadeMux I__2107 (
            .O(N__13136),
            .I(N__13130));
    CascadeBuf I__2106 (
            .O(N__13133),
            .I(N__13127));
    CascadeBuf I__2105 (
            .O(N__13130),
            .I(N__13124));
    CascadeMux I__2104 (
            .O(N__13127),
            .I(N__13121));
    CascadeMux I__2103 (
            .O(N__13124),
            .I(N__13118));
    CascadeBuf I__2102 (
            .O(N__13121),
            .I(N__13115));
    CascadeBuf I__2101 (
            .O(N__13118),
            .I(N__13112));
    CascadeMux I__2100 (
            .O(N__13115),
            .I(N__13109));
    CascadeMux I__2099 (
            .O(N__13112),
            .I(N__13106));
    CascadeBuf I__2098 (
            .O(N__13109),
            .I(N__13103));
    CascadeBuf I__2097 (
            .O(N__13106),
            .I(N__13100));
    CascadeMux I__2096 (
            .O(N__13103),
            .I(N__13097));
    CascadeMux I__2095 (
            .O(N__13100),
            .I(N__13094));
    CascadeBuf I__2094 (
            .O(N__13097),
            .I(N__13091));
    CascadeBuf I__2093 (
            .O(N__13094),
            .I(N__13088));
    CascadeMux I__2092 (
            .O(N__13091),
            .I(N__13085));
    CascadeMux I__2091 (
            .O(N__13088),
            .I(N__13082));
    CascadeBuf I__2090 (
            .O(N__13085),
            .I(N__13079));
    CascadeBuf I__2089 (
            .O(N__13082),
            .I(N__13076));
    CascadeMux I__2088 (
            .O(N__13079),
            .I(N__13073));
    CascadeMux I__2087 (
            .O(N__13076),
            .I(N__13070));
    CascadeBuf I__2086 (
            .O(N__13073),
            .I(N__13067));
    CascadeBuf I__2085 (
            .O(N__13070),
            .I(N__13064));
    CascadeMux I__2084 (
            .O(N__13067),
            .I(N__13061));
    CascadeMux I__2083 (
            .O(N__13064),
            .I(N__13058));
    CascadeBuf I__2082 (
            .O(N__13061),
            .I(N__13055));
    InMux I__2081 (
            .O(N__13058),
            .I(N__13052));
    CascadeMux I__2080 (
            .O(N__13055),
            .I(N__13049));
    LocalMux I__2079 (
            .O(N__13052),
            .I(N__13046));
    InMux I__2078 (
            .O(N__13049),
            .I(N__13043));
    Span12Mux_h I__2077 (
            .O(N__13046),
            .I(N__13040));
    LocalMux I__2076 (
            .O(N__13043),
            .I(N__13037));
    Span12Mux_v I__2075 (
            .O(N__13040),
            .I(N__13032));
    Span12Mux_v I__2074 (
            .O(N__13037),
            .I(N__13032));
    Odrv12 I__2073 (
            .O(N__13032),
            .I(n24));
    InMux I__2072 (
            .O(N__13029),
            .I(N__13026));
    LocalMux I__2071 (
            .O(N__13026),
            .I(N__13023));
    Odrv12 I__2070 (
            .O(N__13023),
            .I(\transmit_module.n125 ));
    InMux I__2069 (
            .O(N__13020),
            .I(N__13017));
    LocalMux I__2068 (
            .O(N__13017),
            .I(N__13014));
    Span4Mux_h I__2067 (
            .O(N__13014),
            .I(N__13011));
    Odrv4 I__2066 (
            .O(N__13011),
            .I(\transmit_module.n140 ));
    CascadeMux I__2065 (
            .O(N__13008),
            .I(\transmit_module.n140_cascade_ ));
    CascadeMux I__2064 (
            .O(N__13005),
            .I(N__13002));
    InMux I__2063 (
            .O(N__13002),
            .I(N__12999));
    LocalMux I__2062 (
            .O(N__12999),
            .I(N__12996));
    Span4Mux_h I__2061 (
            .O(N__12996),
            .I(N__12992));
    InMux I__2060 (
            .O(N__12995),
            .I(N__12989));
    Odrv4 I__2059 (
            .O(N__12992),
            .I(\transmit_module.n109 ));
    LocalMux I__2058 (
            .O(N__12989),
            .I(\transmit_module.n109 ));
    CascadeMux I__2057 (
            .O(N__12984),
            .I(N__12981));
    CascadeBuf I__2056 (
            .O(N__12981),
            .I(N__12977));
    CascadeMux I__2055 (
            .O(N__12980),
            .I(N__12974));
    CascadeMux I__2054 (
            .O(N__12977),
            .I(N__12971));
    CascadeBuf I__2053 (
            .O(N__12974),
            .I(N__12968));
    CascadeBuf I__2052 (
            .O(N__12971),
            .I(N__12965));
    CascadeMux I__2051 (
            .O(N__12968),
            .I(N__12962));
    CascadeMux I__2050 (
            .O(N__12965),
            .I(N__12959));
    CascadeBuf I__2049 (
            .O(N__12962),
            .I(N__12956));
    CascadeBuf I__2048 (
            .O(N__12959),
            .I(N__12953));
    CascadeMux I__2047 (
            .O(N__12956),
            .I(N__12950));
    CascadeMux I__2046 (
            .O(N__12953),
            .I(N__12947));
    CascadeBuf I__2045 (
            .O(N__12950),
            .I(N__12944));
    CascadeBuf I__2044 (
            .O(N__12947),
            .I(N__12941));
    CascadeMux I__2043 (
            .O(N__12944),
            .I(N__12938));
    CascadeMux I__2042 (
            .O(N__12941),
            .I(N__12935));
    CascadeBuf I__2041 (
            .O(N__12938),
            .I(N__12932));
    CascadeBuf I__2040 (
            .O(N__12935),
            .I(N__12929));
    CascadeMux I__2039 (
            .O(N__12932),
            .I(N__12926));
    CascadeMux I__2038 (
            .O(N__12929),
            .I(N__12923));
    CascadeBuf I__2037 (
            .O(N__12926),
            .I(N__12920));
    CascadeBuf I__2036 (
            .O(N__12923),
            .I(N__12917));
    CascadeMux I__2035 (
            .O(N__12920),
            .I(N__12914));
    CascadeMux I__2034 (
            .O(N__12917),
            .I(N__12911));
    CascadeBuf I__2033 (
            .O(N__12914),
            .I(N__12908));
    CascadeBuf I__2032 (
            .O(N__12911),
            .I(N__12905));
    CascadeMux I__2031 (
            .O(N__12908),
            .I(N__12902));
    CascadeMux I__2030 (
            .O(N__12905),
            .I(N__12899));
    CascadeBuf I__2029 (
            .O(N__12902),
            .I(N__12896));
    CascadeBuf I__2028 (
            .O(N__12899),
            .I(N__12893));
    CascadeMux I__2027 (
            .O(N__12896),
            .I(N__12890));
    CascadeMux I__2026 (
            .O(N__12893),
            .I(N__12887));
    CascadeBuf I__2025 (
            .O(N__12890),
            .I(N__12884));
    CascadeBuf I__2024 (
            .O(N__12887),
            .I(N__12881));
    CascadeMux I__2023 (
            .O(N__12884),
            .I(N__12878));
    CascadeMux I__2022 (
            .O(N__12881),
            .I(N__12875));
    CascadeBuf I__2021 (
            .O(N__12878),
            .I(N__12872));
    CascadeBuf I__2020 (
            .O(N__12875),
            .I(N__12869));
    CascadeMux I__2019 (
            .O(N__12872),
            .I(N__12866));
    CascadeMux I__2018 (
            .O(N__12869),
            .I(N__12863));
    CascadeBuf I__2017 (
            .O(N__12866),
            .I(N__12860));
    CascadeBuf I__2016 (
            .O(N__12863),
            .I(N__12857));
    CascadeMux I__2015 (
            .O(N__12860),
            .I(N__12854));
    CascadeMux I__2014 (
            .O(N__12857),
            .I(N__12851));
    CascadeBuf I__2013 (
            .O(N__12854),
            .I(N__12848));
    CascadeBuf I__2012 (
            .O(N__12851),
            .I(N__12845));
    CascadeMux I__2011 (
            .O(N__12848),
            .I(N__12842));
    CascadeMux I__2010 (
            .O(N__12845),
            .I(N__12839));
    CascadeBuf I__2009 (
            .O(N__12842),
            .I(N__12836));
    CascadeBuf I__2008 (
            .O(N__12839),
            .I(N__12833));
    CascadeMux I__2007 (
            .O(N__12836),
            .I(N__12830));
    CascadeMux I__2006 (
            .O(N__12833),
            .I(N__12827));
    CascadeBuf I__2005 (
            .O(N__12830),
            .I(N__12824));
    CascadeBuf I__2004 (
            .O(N__12827),
            .I(N__12821));
    CascadeMux I__2003 (
            .O(N__12824),
            .I(N__12818));
    CascadeMux I__2002 (
            .O(N__12821),
            .I(N__12815));
    CascadeBuf I__2001 (
            .O(N__12818),
            .I(N__12812));
    CascadeBuf I__2000 (
            .O(N__12815),
            .I(N__12809));
    CascadeMux I__1999 (
            .O(N__12812),
            .I(N__12806));
    CascadeMux I__1998 (
            .O(N__12809),
            .I(N__12803));
    CascadeBuf I__1997 (
            .O(N__12806),
            .I(N__12800));
    InMux I__1996 (
            .O(N__12803),
            .I(N__12797));
    CascadeMux I__1995 (
            .O(N__12800),
            .I(N__12794));
    LocalMux I__1994 (
            .O(N__12797),
            .I(N__12791));
    InMux I__1993 (
            .O(N__12794),
            .I(N__12788));
    Span4Mux_v I__1992 (
            .O(N__12791),
            .I(N__12785));
    LocalMux I__1991 (
            .O(N__12788),
            .I(N__12782));
    Span4Mux_v I__1990 (
            .O(N__12785),
            .I(N__12779));
    Span4Mux_v I__1989 (
            .O(N__12782),
            .I(N__12776));
    Span4Mux_v I__1988 (
            .O(N__12779),
            .I(N__12773));
    Span4Mux_v I__1987 (
            .O(N__12776),
            .I(N__12770));
    Span4Mux_h I__1986 (
            .O(N__12773),
            .I(N__12767));
    Span4Mux_v I__1985 (
            .O(N__12770),
            .I(N__12764));
    Span4Mux_h I__1984 (
            .O(N__12767),
            .I(N__12759));
    Span4Mux_h I__1983 (
            .O(N__12764),
            .I(N__12759));
    Odrv4 I__1982 (
            .O(N__12759),
            .I(n21));
    InMux I__1981 (
            .O(N__12756),
            .I(N__12752));
    InMux I__1980 (
            .O(N__12755),
            .I(N__12749));
    LocalMux I__1979 (
            .O(N__12752),
            .I(\transmit_module.n106 ));
    LocalMux I__1978 (
            .O(N__12749),
            .I(\transmit_module.n106 ));
    InMux I__1977 (
            .O(N__12744),
            .I(N__12740));
    InMux I__1976 (
            .O(N__12743),
            .I(N__12737));
    LocalMux I__1975 (
            .O(N__12740),
            .I(\transmit_module.n137 ));
    LocalMux I__1974 (
            .O(N__12737),
            .I(\transmit_module.n137 ));
    CascadeMux I__1973 (
            .O(N__12732),
            .I(N__12729));
    CascadeBuf I__1972 (
            .O(N__12729),
            .I(N__12725));
    CascadeMux I__1971 (
            .O(N__12728),
            .I(N__12722));
    CascadeMux I__1970 (
            .O(N__12725),
            .I(N__12719));
    CascadeBuf I__1969 (
            .O(N__12722),
            .I(N__12716));
    CascadeBuf I__1968 (
            .O(N__12719),
            .I(N__12713));
    CascadeMux I__1967 (
            .O(N__12716),
            .I(N__12710));
    CascadeMux I__1966 (
            .O(N__12713),
            .I(N__12707));
    CascadeBuf I__1965 (
            .O(N__12710),
            .I(N__12704));
    CascadeBuf I__1964 (
            .O(N__12707),
            .I(N__12701));
    CascadeMux I__1963 (
            .O(N__12704),
            .I(N__12698));
    CascadeMux I__1962 (
            .O(N__12701),
            .I(N__12695));
    CascadeBuf I__1961 (
            .O(N__12698),
            .I(N__12692));
    CascadeBuf I__1960 (
            .O(N__12695),
            .I(N__12689));
    CascadeMux I__1959 (
            .O(N__12692),
            .I(N__12686));
    CascadeMux I__1958 (
            .O(N__12689),
            .I(N__12683));
    CascadeBuf I__1957 (
            .O(N__12686),
            .I(N__12680));
    CascadeBuf I__1956 (
            .O(N__12683),
            .I(N__12677));
    CascadeMux I__1955 (
            .O(N__12680),
            .I(N__12674));
    CascadeMux I__1954 (
            .O(N__12677),
            .I(N__12671));
    CascadeBuf I__1953 (
            .O(N__12674),
            .I(N__12668));
    CascadeBuf I__1952 (
            .O(N__12671),
            .I(N__12665));
    CascadeMux I__1951 (
            .O(N__12668),
            .I(N__12662));
    CascadeMux I__1950 (
            .O(N__12665),
            .I(N__12659));
    CascadeBuf I__1949 (
            .O(N__12662),
            .I(N__12656));
    CascadeBuf I__1948 (
            .O(N__12659),
            .I(N__12653));
    CascadeMux I__1947 (
            .O(N__12656),
            .I(N__12650));
    CascadeMux I__1946 (
            .O(N__12653),
            .I(N__12647));
    CascadeBuf I__1945 (
            .O(N__12650),
            .I(N__12644));
    CascadeBuf I__1944 (
            .O(N__12647),
            .I(N__12641));
    CascadeMux I__1943 (
            .O(N__12644),
            .I(N__12638));
    CascadeMux I__1942 (
            .O(N__12641),
            .I(N__12635));
    CascadeBuf I__1941 (
            .O(N__12638),
            .I(N__12632));
    CascadeBuf I__1940 (
            .O(N__12635),
            .I(N__12629));
    CascadeMux I__1939 (
            .O(N__12632),
            .I(N__12626));
    CascadeMux I__1938 (
            .O(N__12629),
            .I(N__12623));
    CascadeBuf I__1937 (
            .O(N__12626),
            .I(N__12620));
    CascadeBuf I__1936 (
            .O(N__12623),
            .I(N__12617));
    CascadeMux I__1935 (
            .O(N__12620),
            .I(N__12614));
    CascadeMux I__1934 (
            .O(N__12617),
            .I(N__12611));
    CascadeBuf I__1933 (
            .O(N__12614),
            .I(N__12608));
    CascadeBuf I__1932 (
            .O(N__12611),
            .I(N__12605));
    CascadeMux I__1931 (
            .O(N__12608),
            .I(N__12602));
    CascadeMux I__1930 (
            .O(N__12605),
            .I(N__12599));
    CascadeBuf I__1929 (
            .O(N__12602),
            .I(N__12596));
    CascadeBuf I__1928 (
            .O(N__12599),
            .I(N__12593));
    CascadeMux I__1927 (
            .O(N__12596),
            .I(N__12590));
    CascadeMux I__1926 (
            .O(N__12593),
            .I(N__12587));
    CascadeBuf I__1925 (
            .O(N__12590),
            .I(N__12584));
    CascadeBuf I__1924 (
            .O(N__12587),
            .I(N__12581));
    CascadeMux I__1923 (
            .O(N__12584),
            .I(N__12578));
    CascadeMux I__1922 (
            .O(N__12581),
            .I(N__12575));
    CascadeBuf I__1921 (
            .O(N__12578),
            .I(N__12572));
    CascadeBuf I__1920 (
            .O(N__12575),
            .I(N__12569));
    CascadeMux I__1919 (
            .O(N__12572),
            .I(N__12566));
    CascadeMux I__1918 (
            .O(N__12569),
            .I(N__12563));
    CascadeBuf I__1917 (
            .O(N__12566),
            .I(N__12560));
    CascadeBuf I__1916 (
            .O(N__12563),
            .I(N__12557));
    CascadeMux I__1915 (
            .O(N__12560),
            .I(N__12554));
    CascadeMux I__1914 (
            .O(N__12557),
            .I(N__12551));
    CascadeBuf I__1913 (
            .O(N__12554),
            .I(N__12548));
    InMux I__1912 (
            .O(N__12551),
            .I(N__12545));
    CascadeMux I__1911 (
            .O(N__12548),
            .I(N__12542));
    LocalMux I__1910 (
            .O(N__12545),
            .I(N__12539));
    InMux I__1909 (
            .O(N__12542),
            .I(N__12536));
    Span4Mux_v I__1908 (
            .O(N__12539),
            .I(N__12533));
    LocalMux I__1907 (
            .O(N__12536),
            .I(N__12530));
    Span4Mux_v I__1906 (
            .O(N__12533),
            .I(N__12527));
    Span4Mux_v I__1905 (
            .O(N__12530),
            .I(N__12524));
    Span4Mux_v I__1904 (
            .O(N__12527),
            .I(N__12521));
    Span4Mux_v I__1903 (
            .O(N__12524),
            .I(N__12518));
    Span4Mux_h I__1902 (
            .O(N__12521),
            .I(N__12515));
    Span4Mux_v I__1901 (
            .O(N__12518),
            .I(N__12512));
    Span4Mux_h I__1900 (
            .O(N__12515),
            .I(N__12507));
    Span4Mux_h I__1899 (
            .O(N__12512),
            .I(N__12507));
    Odrv4 I__1898 (
            .O(N__12507),
            .I(n18));
    InMux I__1897 (
            .O(N__12504),
            .I(\transmit_module.n3171 ));
    CascadeMux I__1896 (
            .O(N__12501),
            .I(N__12495));
    InMux I__1895 (
            .O(N__12500),
            .I(N__12492));
    InMux I__1894 (
            .O(N__12499),
            .I(N__12489));
    InMux I__1893 (
            .O(N__12498),
            .I(N__12484));
    InMux I__1892 (
            .O(N__12495),
            .I(N__12484));
    LocalMux I__1891 (
            .O(N__12492),
            .I(\transmit_module.TX_ADDR_9 ));
    LocalMux I__1890 (
            .O(N__12489),
            .I(\transmit_module.TX_ADDR_9 ));
    LocalMux I__1889 (
            .O(N__12484),
            .I(\transmit_module.TX_ADDR_9 ));
    InMux I__1888 (
            .O(N__12477),
            .I(N__12474));
    LocalMux I__1887 (
            .O(N__12474),
            .I(\transmit_module.ADDR_Y_COMPONENT_9 ));
    InMux I__1886 (
            .O(N__12471),
            .I(N__12468));
    LocalMux I__1885 (
            .O(N__12468),
            .I(N__12465));
    Odrv4 I__1884 (
            .O(N__12465),
            .I(\transmit_module.ADDR_Y_COMPONENT_0 ));
    InMux I__1883 (
            .O(N__12462),
            .I(N__12457));
    InMux I__1882 (
            .O(N__12461),
            .I(N__12454));
    InMux I__1881 (
            .O(N__12460),
            .I(N__12450));
    LocalMux I__1880 (
            .O(N__12457),
            .I(N__12445));
    LocalMux I__1879 (
            .O(N__12454),
            .I(N__12445));
    InMux I__1878 (
            .O(N__12453),
            .I(N__12442));
    LocalMux I__1877 (
            .O(N__12450),
            .I(\transmit_module.TX_ADDR_1 ));
    Odrv4 I__1876 (
            .O(N__12445),
            .I(\transmit_module.TX_ADDR_1 ));
    LocalMux I__1875 (
            .O(N__12442),
            .I(\transmit_module.TX_ADDR_1 ));
    InMux I__1874 (
            .O(N__12435),
            .I(N__12432));
    LocalMux I__1873 (
            .O(N__12432),
            .I(\transmit_module.ADDR_Y_COMPONENT_1 ));
    CascadeMux I__1872 (
            .O(N__12429),
            .I(N__12423));
    InMux I__1871 (
            .O(N__12428),
            .I(N__12420));
    InMux I__1870 (
            .O(N__12427),
            .I(N__12415));
    InMux I__1869 (
            .O(N__12426),
            .I(N__12415));
    InMux I__1868 (
            .O(N__12423),
            .I(N__12412));
    LocalMux I__1867 (
            .O(N__12420),
            .I(\transmit_module.TX_ADDR_8 ));
    LocalMux I__1866 (
            .O(N__12415),
            .I(\transmit_module.TX_ADDR_8 ));
    LocalMux I__1865 (
            .O(N__12412),
            .I(\transmit_module.TX_ADDR_8 ));
    InMux I__1864 (
            .O(N__12405),
            .I(N__12402));
    LocalMux I__1863 (
            .O(N__12402),
            .I(\transmit_module.ADDR_Y_COMPONENT_8 ));
    CascadeMux I__1862 (
            .O(N__12399),
            .I(N__12393));
    InMux I__1861 (
            .O(N__12398),
            .I(N__12390));
    InMux I__1860 (
            .O(N__12397),
            .I(N__12385));
    InMux I__1859 (
            .O(N__12396),
            .I(N__12385));
    InMux I__1858 (
            .O(N__12393),
            .I(N__12382));
    LocalMux I__1857 (
            .O(N__12390),
            .I(\transmit_module.TX_ADDR_5 ));
    LocalMux I__1856 (
            .O(N__12385),
            .I(\transmit_module.TX_ADDR_5 ));
    LocalMux I__1855 (
            .O(N__12382),
            .I(\transmit_module.TX_ADDR_5 ));
    InMux I__1854 (
            .O(N__12375),
            .I(N__12372));
    LocalMux I__1853 (
            .O(N__12372),
            .I(\transmit_module.ADDR_Y_COMPONENT_5 ));
    InMux I__1852 (
            .O(N__12369),
            .I(N__12366));
    LocalMux I__1851 (
            .O(N__12366),
            .I(N__12363));
    Span4Mux_h I__1850 (
            .O(N__12363),
            .I(N__12357));
    InMux I__1849 (
            .O(N__12362),
            .I(N__12354));
    InMux I__1848 (
            .O(N__12361),
            .I(N__12351));
    InMux I__1847 (
            .O(N__12360),
            .I(N__12348));
    Odrv4 I__1846 (
            .O(N__12357),
            .I(\transmit_module.TX_ADDR_10 ));
    LocalMux I__1845 (
            .O(N__12354),
            .I(\transmit_module.TX_ADDR_10 ));
    LocalMux I__1844 (
            .O(N__12351),
            .I(\transmit_module.TX_ADDR_10 ));
    LocalMux I__1843 (
            .O(N__12348),
            .I(\transmit_module.TX_ADDR_10 ));
    InMux I__1842 (
            .O(N__12339),
            .I(N__12336));
    LocalMux I__1841 (
            .O(N__12336),
            .I(N__12333));
    Odrv4 I__1840 (
            .O(N__12333),
            .I(\transmit_module.n122 ));
    InMux I__1839 (
            .O(N__12330),
            .I(\transmit_module.n3162 ));
    CascadeMux I__1838 (
            .O(N__12327),
            .I(N__12324));
    InMux I__1837 (
            .O(N__12324),
            .I(N__12321));
    LocalMux I__1836 (
            .O(N__12321),
            .I(N__12318));
    Odrv4 I__1835 (
            .O(N__12318),
            .I(\transmit_module.n127 ));
    InMux I__1834 (
            .O(N__12315),
            .I(\transmit_module.n3163 ));
    InMux I__1833 (
            .O(N__12312),
            .I(\transmit_module.n3164 ));
    InMux I__1832 (
            .O(N__12309),
            .I(\transmit_module.n3165 ));
    InMux I__1831 (
            .O(N__12306),
            .I(N__12303));
    LocalMux I__1830 (
            .O(N__12303),
            .I(N__12300));
    Odrv4 I__1829 (
            .O(N__12300),
            .I(\transmit_module.n124 ));
    InMux I__1828 (
            .O(N__12297),
            .I(bfn_14_16_0_));
    InMux I__1827 (
            .O(N__12294),
            .I(N__12291));
    LocalMux I__1826 (
            .O(N__12291),
            .I(\transmit_module.n123 ));
    InMux I__1825 (
            .O(N__12288),
            .I(\transmit_module.n3167 ));
    InMux I__1824 (
            .O(N__12285),
            .I(\transmit_module.n3168 ));
    InMux I__1823 (
            .O(N__12282),
            .I(\transmit_module.n3169 ));
    InMux I__1822 (
            .O(N__12279),
            .I(\transmit_module.n3170 ));
    CascadeMux I__1821 (
            .O(N__12276),
            .I(\transmit_module.video_signal_controller.n6_adj_623_cascade_ ));
    InMux I__1820 (
            .O(N__12273),
            .I(N__12269));
    InMux I__1819 (
            .O(N__12272),
            .I(N__12266));
    LocalMux I__1818 (
            .O(N__12269),
            .I(N__12263));
    LocalMux I__1817 (
            .O(N__12266),
            .I(\transmit_module.video_signal_controller.VGA_VISIBLE_N_588 ));
    Odrv4 I__1816 (
            .O(N__12263),
            .I(\transmit_module.video_signal_controller.VGA_VISIBLE_N_588 ));
    InMux I__1815 (
            .O(N__12258),
            .I(N__12252));
    InMux I__1814 (
            .O(N__12257),
            .I(N__12249));
    CascadeMux I__1813 (
            .O(N__12256),
            .I(N__12246));
    InMux I__1812 (
            .O(N__12255),
            .I(N__12243));
    LocalMux I__1811 (
            .O(N__12252),
            .I(N__12237));
    LocalMux I__1810 (
            .O(N__12249),
            .I(N__12237));
    InMux I__1809 (
            .O(N__12246),
            .I(N__12234));
    LocalMux I__1808 (
            .O(N__12243),
            .I(N__12231));
    InMux I__1807 (
            .O(N__12242),
            .I(N__12228));
    Span4Mux_h I__1806 (
            .O(N__12237),
            .I(N__12225));
    LocalMux I__1805 (
            .O(N__12234),
            .I(N__12220));
    Span4Mux_h I__1804 (
            .O(N__12231),
            .I(N__12220));
    LocalMux I__1803 (
            .O(N__12228),
            .I(\transmit_module.video_signal_controller.VGA_X_11 ));
    Odrv4 I__1802 (
            .O(N__12225),
            .I(\transmit_module.video_signal_controller.VGA_X_11 ));
    Odrv4 I__1801 (
            .O(N__12220),
            .I(\transmit_module.video_signal_controller.VGA_X_11 ));
    CascadeMux I__1800 (
            .O(N__12213),
            .I(\transmit_module.video_signal_controller.n7_adj_624_cascade_ ));
    InMux I__1799 (
            .O(N__12210),
            .I(N__12204));
    InMux I__1798 (
            .O(N__12209),
            .I(N__12204));
    LocalMux I__1797 (
            .O(N__12204),
            .I(\transmit_module.video_signal_controller.n3004 ));
    InMux I__1796 (
            .O(N__12201),
            .I(N__12194));
    InMux I__1795 (
            .O(N__12200),
            .I(N__12194));
    InMux I__1794 (
            .O(N__12199),
            .I(N__12190));
    LocalMux I__1793 (
            .O(N__12194),
            .I(N__12186));
    InMux I__1792 (
            .O(N__12193),
            .I(N__12183));
    LocalMux I__1791 (
            .O(N__12190),
            .I(N__12180));
    InMux I__1790 (
            .O(N__12189),
            .I(N__12177));
    Span4Mux_h I__1789 (
            .O(N__12186),
            .I(N__12174));
    LocalMux I__1788 (
            .O(N__12183),
            .I(N__12169));
    Span4Mux_h I__1787 (
            .O(N__12180),
            .I(N__12169));
    LocalMux I__1786 (
            .O(N__12177),
            .I(\transmit_module.video_signal_controller.VGA_X_10 ));
    Odrv4 I__1785 (
            .O(N__12174),
            .I(\transmit_module.video_signal_controller.VGA_X_10 ));
    Odrv4 I__1784 (
            .O(N__12169),
            .I(\transmit_module.video_signal_controller.VGA_X_10 ));
    InMux I__1783 (
            .O(N__12162),
            .I(N__12156));
    InMux I__1782 (
            .O(N__12161),
            .I(N__12151));
    InMux I__1781 (
            .O(N__12160),
            .I(N__12151));
    InMux I__1780 (
            .O(N__12159),
            .I(N__12147));
    LocalMux I__1779 (
            .O(N__12156),
            .I(N__12144));
    LocalMux I__1778 (
            .O(N__12151),
            .I(N__12141));
    InMux I__1777 (
            .O(N__12150),
            .I(N__12138));
    LocalMux I__1776 (
            .O(N__12147),
            .I(N__12133));
    Span4Mux_h I__1775 (
            .O(N__12144),
            .I(N__12133));
    Span4Mux_h I__1774 (
            .O(N__12141),
            .I(N__12130));
    LocalMux I__1773 (
            .O(N__12138),
            .I(\transmit_module.video_signal_controller.VGA_X_9 ));
    Odrv4 I__1772 (
            .O(N__12133),
            .I(\transmit_module.video_signal_controller.VGA_X_9 ));
    Odrv4 I__1771 (
            .O(N__12130),
            .I(\transmit_module.video_signal_controller.VGA_X_9 ));
    InMux I__1770 (
            .O(N__12123),
            .I(N__12120));
    LocalMux I__1769 (
            .O(N__12120),
            .I(\transmit_module.video_signal_controller.n3014 ));
    InMux I__1768 (
            .O(N__12117),
            .I(N__12114));
    LocalMux I__1767 (
            .O(N__12114),
            .I(\transmit_module.n131 ));
    InMux I__1766 (
            .O(N__12111),
            .I(\transmit_module.n3159 ));
    InMux I__1765 (
            .O(N__12108),
            .I(N__12101));
    InMux I__1764 (
            .O(N__12107),
            .I(N__12101));
    InMux I__1763 (
            .O(N__12106),
            .I(N__12097));
    LocalMux I__1762 (
            .O(N__12101),
            .I(N__12094));
    InMux I__1761 (
            .O(N__12100),
            .I(N__12091));
    LocalMux I__1760 (
            .O(N__12097),
            .I(\transmit_module.TX_ADDR_2 ));
    Odrv4 I__1759 (
            .O(N__12094),
            .I(\transmit_module.TX_ADDR_2 ));
    LocalMux I__1758 (
            .O(N__12091),
            .I(\transmit_module.TX_ADDR_2 ));
    InMux I__1757 (
            .O(N__12084),
            .I(N__12081));
    LocalMux I__1756 (
            .O(N__12081),
            .I(\transmit_module.n130 ));
    InMux I__1755 (
            .O(N__12078),
            .I(\transmit_module.n3160 ));
    InMux I__1754 (
            .O(N__12075),
            .I(N__12070));
    InMux I__1753 (
            .O(N__12074),
            .I(N__12065));
    InMux I__1752 (
            .O(N__12073),
            .I(N__12065));
    LocalMux I__1751 (
            .O(N__12070),
            .I(N__12061));
    LocalMux I__1750 (
            .O(N__12065),
            .I(N__12058));
    InMux I__1749 (
            .O(N__12064),
            .I(N__12055));
    Odrv12 I__1748 (
            .O(N__12061),
            .I(\transmit_module.TX_ADDR_3 ));
    Odrv4 I__1747 (
            .O(N__12058),
            .I(\transmit_module.TX_ADDR_3 ));
    LocalMux I__1746 (
            .O(N__12055),
            .I(\transmit_module.TX_ADDR_3 ));
    InMux I__1745 (
            .O(N__12048),
            .I(N__12045));
    LocalMux I__1744 (
            .O(N__12045),
            .I(N__12042));
    Span4Mux_v I__1743 (
            .O(N__12042),
            .I(N__12039));
    Odrv4 I__1742 (
            .O(N__12039),
            .I(\transmit_module.n129 ));
    InMux I__1741 (
            .O(N__12036),
            .I(\transmit_module.n3161 ));
    InMux I__1740 (
            .O(N__12033),
            .I(N__12030));
    LocalMux I__1739 (
            .O(N__12030),
            .I(N__12027));
    Span4Mux_v I__1738 (
            .O(N__12027),
            .I(N__12021));
    InMux I__1737 (
            .O(N__12026),
            .I(N__12018));
    InMux I__1736 (
            .O(N__12025),
            .I(N__12013));
    InMux I__1735 (
            .O(N__12024),
            .I(N__12013));
    Odrv4 I__1734 (
            .O(N__12021),
            .I(\transmit_module.video_signal_controller.VGA_Y_2 ));
    LocalMux I__1733 (
            .O(N__12018),
            .I(\transmit_module.video_signal_controller.VGA_Y_2 ));
    LocalMux I__1732 (
            .O(N__12013),
            .I(\transmit_module.video_signal_controller.VGA_Y_2 ));
    InMux I__1731 (
            .O(N__12006),
            .I(N__12003));
    LocalMux I__1730 (
            .O(N__12003),
            .I(\transmit_module.video_signal_controller.n3517 ));
    CascadeMux I__1729 (
            .O(N__12000),
            .I(N__11997));
    InMux I__1728 (
            .O(N__11997),
            .I(N__11994));
    LocalMux I__1727 (
            .O(N__11994),
            .I(N__11988));
    InMux I__1726 (
            .O(N__11993),
            .I(N__11985));
    InMux I__1725 (
            .O(N__11992),
            .I(N__11980));
    InMux I__1724 (
            .O(N__11991),
            .I(N__11980));
    Odrv4 I__1723 (
            .O(N__11988),
            .I(\transmit_module.video_signal_controller.VGA_Y_1 ));
    LocalMux I__1722 (
            .O(N__11985),
            .I(\transmit_module.video_signal_controller.VGA_Y_1 ));
    LocalMux I__1721 (
            .O(N__11980),
            .I(\transmit_module.video_signal_controller.VGA_Y_1 ));
    InMux I__1720 (
            .O(N__11973),
            .I(N__11969));
    InMux I__1719 (
            .O(N__11972),
            .I(N__11966));
    LocalMux I__1718 (
            .O(N__11969),
            .I(\transmit_module.video_signal_controller.VGA_Y_0 ));
    LocalMux I__1717 (
            .O(N__11966),
            .I(\transmit_module.video_signal_controller.VGA_Y_0 ));
    InMux I__1716 (
            .O(N__11961),
            .I(N__11958));
    LocalMux I__1715 (
            .O(N__11958),
            .I(\transmit_module.video_signal_controller.n2955 ));
    InMux I__1714 (
            .O(N__11955),
            .I(N__11950));
    InMux I__1713 (
            .O(N__11954),
            .I(N__11944));
    InMux I__1712 (
            .O(N__11953),
            .I(N__11944));
    LocalMux I__1711 (
            .O(N__11950),
            .I(N__11941));
    InMux I__1710 (
            .O(N__11949),
            .I(N__11938));
    LocalMux I__1709 (
            .O(N__11944),
            .I(N__11933));
    Span4Mux_h I__1708 (
            .O(N__11941),
            .I(N__11933));
    LocalMux I__1707 (
            .O(N__11938),
            .I(\transmit_module.video_signal_controller.VGA_X_8 ));
    Odrv4 I__1706 (
            .O(N__11933),
            .I(\transmit_module.video_signal_controller.VGA_X_8 ));
    CascadeMux I__1705 (
            .O(N__11928),
            .I(N__11924));
    InMux I__1704 (
            .O(N__11927),
            .I(N__11921));
    InMux I__1703 (
            .O(N__11924),
            .I(N__11918));
    LocalMux I__1702 (
            .O(N__11921),
            .I(\transmit_module.video_signal_controller.n3363 ));
    LocalMux I__1701 (
            .O(N__11918),
            .I(\transmit_module.video_signal_controller.n3363 ));
    InMux I__1700 (
            .O(N__11913),
            .I(N__11910));
    LocalMux I__1699 (
            .O(N__11910),
            .I(\transmit_module.video_signal_controller.n2014 ));
    CascadeMux I__1698 (
            .O(N__11907),
            .I(\transmit_module.video_signal_controller.n2972_cascade_ ));
    SRMux I__1697 (
            .O(N__11904),
            .I(N__11901));
    LocalMux I__1696 (
            .O(N__11901),
            .I(N__11895));
    SRMux I__1695 (
            .O(N__11900),
            .I(N__11892));
    CEMux I__1694 (
            .O(N__11899),
            .I(N__11888));
    CEMux I__1693 (
            .O(N__11898),
            .I(N__11885));
    Span4Mux_h I__1692 (
            .O(N__11895),
            .I(N__11882));
    LocalMux I__1691 (
            .O(N__11892),
            .I(N__11879));
    InMux I__1690 (
            .O(N__11891),
            .I(N__11876));
    LocalMux I__1689 (
            .O(N__11888),
            .I(N__11873));
    LocalMux I__1688 (
            .O(N__11885),
            .I(N__11864));
    Span4Mux_v I__1687 (
            .O(N__11882),
            .I(N__11864));
    Span4Mux_v I__1686 (
            .O(N__11879),
            .I(N__11864));
    LocalMux I__1685 (
            .O(N__11876),
            .I(N__11864));
    Odrv4 I__1684 (
            .O(N__11873),
            .I(\transmit_module.video_signal_controller.n2047 ));
    Odrv4 I__1683 (
            .O(N__11864),
            .I(\transmit_module.video_signal_controller.n2047 ));
    CascadeMux I__1682 (
            .O(N__11859),
            .I(N__11854));
    CascadeMux I__1681 (
            .O(N__11858),
            .I(N__11851));
    InMux I__1680 (
            .O(N__11857),
            .I(N__11847));
    InMux I__1679 (
            .O(N__11854),
            .I(N__11842));
    InMux I__1678 (
            .O(N__11851),
            .I(N__11842));
    InMux I__1677 (
            .O(N__11850),
            .I(N__11839));
    LocalMux I__1676 (
            .O(N__11847),
            .I(\transmit_module.VGA_VISIBLE_Y ));
    LocalMux I__1675 (
            .O(N__11842),
            .I(\transmit_module.VGA_VISIBLE_Y ));
    LocalMux I__1674 (
            .O(N__11839),
            .I(\transmit_module.VGA_VISIBLE_Y ));
    IoInMux I__1673 (
            .O(N__11832),
            .I(N__11829));
    LocalMux I__1672 (
            .O(N__11829),
            .I(N__11826));
    IoSpan4Mux I__1671 (
            .O(N__11826),
            .I(N__11823));
    IoSpan4Mux I__1670 (
            .O(N__11823),
            .I(N__11820));
    Sp12to4 I__1669 (
            .O(N__11820),
            .I(N__11817));
    Span12Mux_h I__1668 (
            .O(N__11817),
            .I(N__11809));
    InMux I__1667 (
            .O(N__11816),
            .I(N__11804));
    InMux I__1666 (
            .O(N__11815),
            .I(N__11804));
    InMux I__1665 (
            .O(N__11814),
            .I(N__11799));
    InMux I__1664 (
            .O(N__11813),
            .I(N__11799));
    InMux I__1663 (
            .O(N__11812),
            .I(N__11796));
    Odrv12 I__1662 (
            .O(N__11809),
            .I(ADV_HSYNC_c));
    LocalMux I__1661 (
            .O(N__11804),
            .I(ADV_HSYNC_c));
    LocalMux I__1660 (
            .O(N__11799),
            .I(ADV_HSYNC_c));
    LocalMux I__1659 (
            .O(N__11796),
            .I(ADV_HSYNC_c));
    InMux I__1658 (
            .O(N__11787),
            .I(N__11781));
    InMux I__1657 (
            .O(N__11786),
            .I(N__11776));
    InMux I__1656 (
            .O(N__11785),
            .I(N__11776));
    InMux I__1655 (
            .O(N__11784),
            .I(N__11773));
    LocalMux I__1654 (
            .O(N__11781),
            .I(\transmit_module.old_VGA_HS ));
    LocalMux I__1653 (
            .O(N__11776),
            .I(\transmit_module.old_VGA_HS ));
    LocalMux I__1652 (
            .O(N__11773),
            .I(\transmit_module.old_VGA_HS ));
    CascadeMux I__1651 (
            .O(N__11766),
            .I(\transmit_module.n3675_cascade_ ));
    CascadeMux I__1650 (
            .O(N__11763),
            .I(\transmit_module.video_signal_controller.n6_adj_622_cascade_ ));
    InMux I__1649 (
            .O(N__11760),
            .I(N__11754));
    InMux I__1648 (
            .O(N__11759),
            .I(N__11747));
    InMux I__1647 (
            .O(N__11758),
            .I(N__11747));
    InMux I__1646 (
            .O(N__11757),
            .I(N__11747));
    LocalMux I__1645 (
            .O(N__11754),
            .I(\transmit_module.video_signal_controller.VGA_Y_3 ));
    LocalMux I__1644 (
            .O(N__11747),
            .I(\transmit_module.video_signal_controller.VGA_Y_3 ));
    InMux I__1643 (
            .O(N__11742),
            .I(N__11736));
    InMux I__1642 (
            .O(N__11741),
            .I(N__11733));
    InMux I__1641 (
            .O(N__11740),
            .I(N__11728));
    InMux I__1640 (
            .O(N__11739),
            .I(N__11728));
    LocalMux I__1639 (
            .O(N__11736),
            .I(\transmit_module.video_signal_controller.VGA_Y_4 ));
    LocalMux I__1638 (
            .O(N__11733),
            .I(\transmit_module.video_signal_controller.VGA_Y_4 ));
    LocalMux I__1637 (
            .O(N__11728),
            .I(\transmit_module.video_signal_controller.VGA_Y_4 ));
    CascadeMux I__1636 (
            .O(N__11721),
            .I(\transmit_module.video_signal_controller.n3482_cascade_ ));
    InMux I__1635 (
            .O(N__11718),
            .I(N__11713));
    InMux I__1634 (
            .O(N__11717),
            .I(N__11708));
    InMux I__1633 (
            .O(N__11716),
            .I(N__11708));
    LocalMux I__1632 (
            .O(N__11713),
            .I(\transmit_module.video_signal_controller.VGA_Y_6 ));
    LocalMux I__1631 (
            .O(N__11708),
            .I(\transmit_module.video_signal_controller.VGA_Y_6 ));
    InMux I__1630 (
            .O(N__11703),
            .I(N__11698));
    InMux I__1629 (
            .O(N__11702),
            .I(N__11693));
    InMux I__1628 (
            .O(N__11701),
            .I(N__11693));
    LocalMux I__1627 (
            .O(N__11698),
            .I(\transmit_module.video_signal_controller.VGA_Y_5 ));
    LocalMux I__1626 (
            .O(N__11693),
            .I(\transmit_module.video_signal_controller.VGA_Y_5 ));
    CascadeMux I__1625 (
            .O(N__11688),
            .I(\transmit_module.video_signal_controller.n6_cascade_ ));
    InMux I__1624 (
            .O(N__11685),
            .I(N__11679));
    InMux I__1623 (
            .O(N__11684),
            .I(N__11679));
    LocalMux I__1622 (
            .O(N__11679),
            .I(\transmit_module.video_signal_controller.n2016 ));
    InMux I__1621 (
            .O(N__11676),
            .I(N__11672));
    InMux I__1620 (
            .O(N__11675),
            .I(N__11669));
    LocalMux I__1619 (
            .O(N__11672),
            .I(\transmit_module.video_signal_controller.VGA_Y_8 ));
    LocalMux I__1618 (
            .O(N__11669),
            .I(\transmit_module.video_signal_controller.VGA_Y_8 ));
    InMux I__1617 (
            .O(N__11664),
            .I(N__11660));
    InMux I__1616 (
            .O(N__11663),
            .I(N__11657));
    LocalMux I__1615 (
            .O(N__11660),
            .I(\transmit_module.video_signal_controller.VGA_Y_7 ));
    LocalMux I__1614 (
            .O(N__11657),
            .I(\transmit_module.video_signal_controller.VGA_Y_7 ));
    InMux I__1613 (
            .O(N__11652),
            .I(N__11649));
    LocalMux I__1612 (
            .O(N__11649),
            .I(\transmit_module.Y_DELTA_PATTERN_20 ));
    InMux I__1611 (
            .O(N__11646),
            .I(N__11643));
    LocalMux I__1610 (
            .O(N__11643),
            .I(\transmit_module.Y_DELTA_PATTERN_21 ));
    InMux I__1609 (
            .O(N__11640),
            .I(N__11637));
    LocalMux I__1608 (
            .O(N__11637),
            .I(\transmit_module.Y_DELTA_PATTERN_22 ));
    InMux I__1607 (
            .O(N__11634),
            .I(N__11631));
    LocalMux I__1606 (
            .O(N__11631),
            .I(\transmit_module.Y_DELTA_PATTERN_24 ));
    InMux I__1605 (
            .O(N__11628),
            .I(N__11625));
    LocalMux I__1604 (
            .O(N__11625),
            .I(\transmit_module.Y_DELTA_PATTERN_23 ));
    InMux I__1603 (
            .O(N__11622),
            .I(N__11619));
    LocalMux I__1602 (
            .O(N__11619),
            .I(N__11616));
    Odrv4 I__1601 (
            .O(N__11616),
            .I(\transmit_module.X_DELTA_PATTERN_13 ));
    InMux I__1600 (
            .O(N__11613),
            .I(N__11610));
    LocalMux I__1599 (
            .O(N__11610),
            .I(\transmit_module.X_DELTA_PATTERN_14 ));
    InMux I__1598 (
            .O(N__11607),
            .I(N__11604));
    LocalMux I__1597 (
            .O(N__11604),
            .I(N__11601));
    Odrv12 I__1596 (
            .O(N__11601),
            .I(\transmit_module.X_DELTA_PATTERN_6 ));
    InMux I__1595 (
            .O(N__11598),
            .I(N__11595));
    LocalMux I__1594 (
            .O(N__11595),
            .I(\transmit_module.X_DELTA_PATTERN_5 ));
    InMux I__1593 (
            .O(N__11592),
            .I(N__11589));
    LocalMux I__1592 (
            .O(N__11589),
            .I(\transmit_module.X_DELTA_PATTERN_4 ));
    InMux I__1591 (
            .O(N__11586),
            .I(N__11583));
    LocalMux I__1590 (
            .O(N__11583),
            .I(\transmit_module.ADDR_Y_COMPONENT_3 ));
    InMux I__1589 (
            .O(N__11580),
            .I(N__11577));
    LocalMux I__1588 (
            .O(N__11577),
            .I(N__11574));
    Span4Mux_h I__1587 (
            .O(N__11574),
            .I(N__11571));
    Span4Mux_h I__1586 (
            .O(N__11571),
            .I(N__11568));
    Odrv4 I__1585 (
            .O(N__11568),
            .I(\line_buffer.n568 ));
    InMux I__1584 (
            .O(N__11565),
            .I(N__11562));
    LocalMux I__1583 (
            .O(N__11562),
            .I(N__11559));
    Span12Mux_v I__1582 (
            .O(N__11559),
            .I(N__11556));
    Span12Mux_v I__1581 (
            .O(N__11556),
            .I(N__11553));
    Span12Mux_h I__1580 (
            .O(N__11553),
            .I(N__11550));
    Odrv12 I__1579 (
            .O(N__11550),
            .I(\line_buffer.n560 ));
    InMux I__1578 (
            .O(N__11547),
            .I(N__11544));
    LocalMux I__1577 (
            .O(N__11544),
            .I(N__11541));
    Span4Mux_h I__1576 (
            .O(N__11541),
            .I(N__11538));
    Odrv4 I__1575 (
            .O(N__11538),
            .I(\line_buffer.n3530 ));
    CascadeMux I__1574 (
            .O(N__11535),
            .I(\line_buffer.n3531_cascade_ ));
    InMux I__1573 (
            .O(N__11532),
            .I(N__11529));
    LocalMux I__1572 (
            .O(N__11529),
            .I(\line_buffer.n3617 ));
    InMux I__1571 (
            .O(N__11526),
            .I(N__11523));
    LocalMux I__1570 (
            .O(N__11523),
            .I(TX_DATA_7));
    IoInMux I__1569 (
            .O(N__11520),
            .I(N__11515));
    IoInMux I__1568 (
            .O(N__11519),
            .I(N__11512));
    IoInMux I__1567 (
            .O(N__11518),
            .I(N__11509));
    LocalMux I__1566 (
            .O(N__11515),
            .I(N__11506));
    LocalMux I__1565 (
            .O(N__11512),
            .I(N__11503));
    LocalMux I__1564 (
            .O(N__11509),
            .I(N__11500));
    IoSpan4Mux I__1563 (
            .O(N__11506),
            .I(N__11497));
    IoSpan4Mux I__1562 (
            .O(N__11503),
            .I(N__11494));
    Span12Mux_s10_v I__1561 (
            .O(N__11500),
            .I(N__11491));
    Sp12to4 I__1560 (
            .O(N__11497),
            .I(N__11488));
    Span4Mux_s3_v I__1559 (
            .O(N__11494),
            .I(N__11485));
    Span12Mux_h I__1558 (
            .O(N__11491),
            .I(N__11482));
    Span12Mux_h I__1557 (
            .O(N__11488),
            .I(N__11479));
    Span4Mux_v I__1556 (
            .O(N__11485),
            .I(N__11476));
    Odrv12 I__1555 (
            .O(N__11482),
            .I(ADV_B_c));
    Odrv12 I__1554 (
            .O(N__11479),
            .I(ADV_B_c));
    Odrv4 I__1553 (
            .O(N__11476),
            .I(ADV_B_c));
    InMux I__1552 (
            .O(N__11469),
            .I(N__11466));
    LocalMux I__1551 (
            .O(N__11466),
            .I(N__11463));
    Span12Mux_h I__1550 (
            .O(N__11463),
            .I(N__11460));
    Odrv12 I__1549 (
            .O(N__11460),
            .I(\transmit_module.Y_DELTA_PATTERN_26 ));
    InMux I__1548 (
            .O(N__11457),
            .I(N__11454));
    LocalMux I__1547 (
            .O(N__11454),
            .I(\transmit_module.Y_DELTA_PATTERN_25 ));
    InMux I__1546 (
            .O(N__11451),
            .I(N__11448));
    LocalMux I__1545 (
            .O(N__11448),
            .I(\transmit_module.Y_DELTA_PATTERN_19 ));
    InMux I__1544 (
            .O(N__11445),
            .I(N__11442));
    LocalMux I__1543 (
            .O(N__11442),
            .I(\transmit_module.n139 ));
    InMux I__1542 (
            .O(N__11439),
            .I(N__11435));
    InMux I__1541 (
            .O(N__11438),
            .I(N__11432));
    LocalMux I__1540 (
            .O(N__11435),
            .I(\transmit_module.n108 ));
    LocalMux I__1539 (
            .O(N__11432),
            .I(\transmit_module.n108 ));
    CascadeMux I__1538 (
            .O(N__11427),
            .I(\transmit_module.n139_cascade_ ));
    CascadeMux I__1537 (
            .O(N__11424),
            .I(N__11421));
    CascadeBuf I__1536 (
            .O(N__11421),
            .I(N__11417));
    CascadeMux I__1535 (
            .O(N__11420),
            .I(N__11414));
    CascadeMux I__1534 (
            .O(N__11417),
            .I(N__11411));
    CascadeBuf I__1533 (
            .O(N__11414),
            .I(N__11408));
    CascadeBuf I__1532 (
            .O(N__11411),
            .I(N__11405));
    CascadeMux I__1531 (
            .O(N__11408),
            .I(N__11402));
    CascadeMux I__1530 (
            .O(N__11405),
            .I(N__11399));
    CascadeBuf I__1529 (
            .O(N__11402),
            .I(N__11396));
    CascadeBuf I__1528 (
            .O(N__11399),
            .I(N__11393));
    CascadeMux I__1527 (
            .O(N__11396),
            .I(N__11390));
    CascadeMux I__1526 (
            .O(N__11393),
            .I(N__11387));
    CascadeBuf I__1525 (
            .O(N__11390),
            .I(N__11384));
    CascadeBuf I__1524 (
            .O(N__11387),
            .I(N__11381));
    CascadeMux I__1523 (
            .O(N__11384),
            .I(N__11378));
    CascadeMux I__1522 (
            .O(N__11381),
            .I(N__11375));
    CascadeBuf I__1521 (
            .O(N__11378),
            .I(N__11372));
    CascadeBuf I__1520 (
            .O(N__11375),
            .I(N__11369));
    CascadeMux I__1519 (
            .O(N__11372),
            .I(N__11366));
    CascadeMux I__1518 (
            .O(N__11369),
            .I(N__11363));
    CascadeBuf I__1517 (
            .O(N__11366),
            .I(N__11360));
    CascadeBuf I__1516 (
            .O(N__11363),
            .I(N__11357));
    CascadeMux I__1515 (
            .O(N__11360),
            .I(N__11354));
    CascadeMux I__1514 (
            .O(N__11357),
            .I(N__11351));
    CascadeBuf I__1513 (
            .O(N__11354),
            .I(N__11348));
    CascadeBuf I__1512 (
            .O(N__11351),
            .I(N__11345));
    CascadeMux I__1511 (
            .O(N__11348),
            .I(N__11342));
    CascadeMux I__1510 (
            .O(N__11345),
            .I(N__11339));
    CascadeBuf I__1509 (
            .O(N__11342),
            .I(N__11336));
    CascadeBuf I__1508 (
            .O(N__11339),
            .I(N__11333));
    CascadeMux I__1507 (
            .O(N__11336),
            .I(N__11330));
    CascadeMux I__1506 (
            .O(N__11333),
            .I(N__11327));
    CascadeBuf I__1505 (
            .O(N__11330),
            .I(N__11324));
    CascadeBuf I__1504 (
            .O(N__11327),
            .I(N__11321));
    CascadeMux I__1503 (
            .O(N__11324),
            .I(N__11318));
    CascadeMux I__1502 (
            .O(N__11321),
            .I(N__11315));
    CascadeBuf I__1501 (
            .O(N__11318),
            .I(N__11312));
    CascadeBuf I__1500 (
            .O(N__11315),
            .I(N__11309));
    CascadeMux I__1499 (
            .O(N__11312),
            .I(N__11306));
    CascadeMux I__1498 (
            .O(N__11309),
            .I(N__11303));
    CascadeBuf I__1497 (
            .O(N__11306),
            .I(N__11300));
    CascadeBuf I__1496 (
            .O(N__11303),
            .I(N__11297));
    CascadeMux I__1495 (
            .O(N__11300),
            .I(N__11294));
    CascadeMux I__1494 (
            .O(N__11297),
            .I(N__11291));
    CascadeBuf I__1493 (
            .O(N__11294),
            .I(N__11288));
    CascadeBuf I__1492 (
            .O(N__11291),
            .I(N__11285));
    CascadeMux I__1491 (
            .O(N__11288),
            .I(N__11282));
    CascadeMux I__1490 (
            .O(N__11285),
            .I(N__11279));
    CascadeBuf I__1489 (
            .O(N__11282),
            .I(N__11276));
    CascadeBuf I__1488 (
            .O(N__11279),
            .I(N__11273));
    CascadeMux I__1487 (
            .O(N__11276),
            .I(N__11270));
    CascadeMux I__1486 (
            .O(N__11273),
            .I(N__11267));
    CascadeBuf I__1485 (
            .O(N__11270),
            .I(N__11264));
    CascadeBuf I__1484 (
            .O(N__11267),
            .I(N__11261));
    CascadeMux I__1483 (
            .O(N__11264),
            .I(N__11258));
    CascadeMux I__1482 (
            .O(N__11261),
            .I(N__11255));
    CascadeBuf I__1481 (
            .O(N__11258),
            .I(N__11252));
    CascadeBuf I__1480 (
            .O(N__11255),
            .I(N__11249));
    CascadeMux I__1479 (
            .O(N__11252),
            .I(N__11246));
    CascadeMux I__1478 (
            .O(N__11249),
            .I(N__11243));
    CascadeBuf I__1477 (
            .O(N__11246),
            .I(N__11240));
    InMux I__1476 (
            .O(N__11243),
            .I(N__11237));
    CascadeMux I__1475 (
            .O(N__11240),
            .I(N__11234));
    LocalMux I__1474 (
            .O(N__11237),
            .I(N__11231));
    InMux I__1473 (
            .O(N__11234),
            .I(N__11228));
    Span4Mux_s3_v I__1472 (
            .O(N__11231),
            .I(N__11225));
    LocalMux I__1471 (
            .O(N__11228),
            .I(N__11222));
    Span4Mux_v I__1470 (
            .O(N__11225),
            .I(N__11219));
    Span12Mux_s10_v I__1469 (
            .O(N__11222),
            .I(N__11216));
    Span4Mux_v I__1468 (
            .O(N__11219),
            .I(N__11213));
    Span12Mux_h I__1467 (
            .O(N__11216),
            .I(N__11210));
    Span4Mux_h I__1466 (
            .O(N__11213),
            .I(N__11207));
    Odrv12 I__1465 (
            .O(N__11210),
            .I(n20));
    Odrv4 I__1464 (
            .O(N__11207),
            .I(n20));
    InMux I__1463 (
            .O(N__11202),
            .I(N__11199));
    LocalMux I__1462 (
            .O(N__11199),
            .I(N__11196));
    Span4Mux_h I__1461 (
            .O(N__11196),
            .I(N__11193));
    Odrv4 I__1460 (
            .O(N__11193),
            .I(\transmit_module.ADDR_Y_COMPONENT_10 ));
    InMux I__1459 (
            .O(N__11190),
            .I(N__11187));
    LocalMux I__1458 (
            .O(N__11187),
            .I(N__11184));
    Odrv4 I__1457 (
            .O(N__11184),
            .I(\transmit_module.n145 ));
    CascadeMux I__1456 (
            .O(N__11181),
            .I(N__11178));
    CascadeBuf I__1455 (
            .O(N__11178),
            .I(N__11175));
    CascadeMux I__1454 (
            .O(N__11175),
            .I(N__11172));
    CascadeBuf I__1453 (
            .O(N__11172),
            .I(N__11168));
    CascadeMux I__1452 (
            .O(N__11171),
            .I(N__11165));
    CascadeMux I__1451 (
            .O(N__11168),
            .I(N__11162));
    CascadeBuf I__1450 (
            .O(N__11165),
            .I(N__11159));
    CascadeBuf I__1449 (
            .O(N__11162),
            .I(N__11156));
    CascadeMux I__1448 (
            .O(N__11159),
            .I(N__11153));
    CascadeMux I__1447 (
            .O(N__11156),
            .I(N__11150));
    CascadeBuf I__1446 (
            .O(N__11153),
            .I(N__11147));
    CascadeBuf I__1445 (
            .O(N__11150),
            .I(N__11144));
    CascadeMux I__1444 (
            .O(N__11147),
            .I(N__11141));
    CascadeMux I__1443 (
            .O(N__11144),
            .I(N__11138));
    CascadeBuf I__1442 (
            .O(N__11141),
            .I(N__11135));
    CascadeBuf I__1441 (
            .O(N__11138),
            .I(N__11132));
    CascadeMux I__1440 (
            .O(N__11135),
            .I(N__11129));
    CascadeMux I__1439 (
            .O(N__11132),
            .I(N__11126));
    CascadeBuf I__1438 (
            .O(N__11129),
            .I(N__11123));
    CascadeBuf I__1437 (
            .O(N__11126),
            .I(N__11120));
    CascadeMux I__1436 (
            .O(N__11123),
            .I(N__11117));
    CascadeMux I__1435 (
            .O(N__11120),
            .I(N__11114));
    CascadeBuf I__1434 (
            .O(N__11117),
            .I(N__11111));
    CascadeBuf I__1433 (
            .O(N__11114),
            .I(N__11108));
    CascadeMux I__1432 (
            .O(N__11111),
            .I(N__11105));
    CascadeMux I__1431 (
            .O(N__11108),
            .I(N__11102));
    CascadeBuf I__1430 (
            .O(N__11105),
            .I(N__11099));
    CascadeBuf I__1429 (
            .O(N__11102),
            .I(N__11096));
    CascadeMux I__1428 (
            .O(N__11099),
            .I(N__11093));
    CascadeMux I__1427 (
            .O(N__11096),
            .I(N__11090));
    CascadeBuf I__1426 (
            .O(N__11093),
            .I(N__11087));
    CascadeBuf I__1425 (
            .O(N__11090),
            .I(N__11084));
    CascadeMux I__1424 (
            .O(N__11087),
            .I(N__11081));
    CascadeMux I__1423 (
            .O(N__11084),
            .I(N__11078));
    CascadeBuf I__1422 (
            .O(N__11081),
            .I(N__11075));
    CascadeBuf I__1421 (
            .O(N__11078),
            .I(N__11072));
    CascadeMux I__1420 (
            .O(N__11075),
            .I(N__11069));
    CascadeMux I__1419 (
            .O(N__11072),
            .I(N__11066));
    CascadeBuf I__1418 (
            .O(N__11069),
            .I(N__11063));
    CascadeBuf I__1417 (
            .O(N__11066),
            .I(N__11060));
    CascadeMux I__1416 (
            .O(N__11063),
            .I(N__11057));
    CascadeMux I__1415 (
            .O(N__11060),
            .I(N__11054));
    CascadeBuf I__1414 (
            .O(N__11057),
            .I(N__11051));
    CascadeBuf I__1413 (
            .O(N__11054),
            .I(N__11048));
    CascadeMux I__1412 (
            .O(N__11051),
            .I(N__11045));
    CascadeMux I__1411 (
            .O(N__11048),
            .I(N__11042));
    CascadeBuf I__1410 (
            .O(N__11045),
            .I(N__11039));
    CascadeBuf I__1409 (
            .O(N__11042),
            .I(N__11036));
    CascadeMux I__1408 (
            .O(N__11039),
            .I(N__11033));
    CascadeMux I__1407 (
            .O(N__11036),
            .I(N__11030));
    CascadeBuf I__1406 (
            .O(N__11033),
            .I(N__11027));
    CascadeBuf I__1405 (
            .O(N__11030),
            .I(N__11024));
    CascadeMux I__1404 (
            .O(N__11027),
            .I(N__11021));
    CascadeMux I__1403 (
            .O(N__11024),
            .I(N__11018));
    CascadeBuf I__1402 (
            .O(N__11021),
            .I(N__11015));
    CascadeBuf I__1401 (
            .O(N__11018),
            .I(N__11012));
    CascadeMux I__1400 (
            .O(N__11015),
            .I(N__11009));
    CascadeMux I__1399 (
            .O(N__11012),
            .I(N__11006));
    CascadeBuf I__1398 (
            .O(N__11009),
            .I(N__11003));
    InMux I__1397 (
            .O(N__11006),
            .I(N__11000));
    CascadeMux I__1396 (
            .O(N__11003),
            .I(N__10997));
    LocalMux I__1395 (
            .O(N__11000),
            .I(N__10994));
    CascadeBuf I__1394 (
            .O(N__10997),
            .I(N__10991));
    Span4Mux_v I__1393 (
            .O(N__10994),
            .I(N__10988));
    CascadeMux I__1392 (
            .O(N__10991),
            .I(N__10985));
    Span4Mux_v I__1391 (
            .O(N__10988),
            .I(N__10982));
    InMux I__1390 (
            .O(N__10985),
            .I(N__10979));
    Span4Mux_v I__1389 (
            .O(N__10982),
            .I(N__10976));
    LocalMux I__1388 (
            .O(N__10979),
            .I(N__10973));
    Span4Mux_h I__1387 (
            .O(N__10976),
            .I(N__10970));
    Sp12to4 I__1386 (
            .O(N__10973),
            .I(N__10967));
    Span4Mux_h I__1385 (
            .O(N__10970),
            .I(N__10964));
    Span12Mux_v I__1384 (
            .O(N__10967),
            .I(N__10961));
    Odrv4 I__1383 (
            .O(N__10964),
            .I(n26));
    Odrv12 I__1382 (
            .O(N__10961),
            .I(n26));
    InMux I__1381 (
            .O(N__10956),
            .I(N__10953));
    LocalMux I__1380 (
            .O(N__10953),
            .I(N__10949));
    InMux I__1379 (
            .O(N__10952),
            .I(N__10946));
    Odrv4 I__1378 (
            .O(N__10949),
            .I(\transmit_module.n114 ));
    LocalMux I__1377 (
            .O(N__10946),
            .I(\transmit_module.n114 ));
    InMux I__1376 (
            .O(N__10941),
            .I(N__10938));
    LocalMux I__1375 (
            .O(N__10938),
            .I(N__10935));
    Odrv4 I__1374 (
            .O(N__10935),
            .I(\transmit_module.n144 ));
    CascadeMux I__1373 (
            .O(N__10932),
            .I(\transmit_module.n144_cascade_ ));
    CascadeMux I__1372 (
            .O(N__10929),
            .I(N__10926));
    CascadeBuf I__1371 (
            .O(N__10926),
            .I(N__10923));
    CascadeMux I__1370 (
            .O(N__10923),
            .I(N__10920));
    CascadeBuf I__1369 (
            .O(N__10920),
            .I(N__10916));
    CascadeMux I__1368 (
            .O(N__10919),
            .I(N__10913));
    CascadeMux I__1367 (
            .O(N__10916),
            .I(N__10910));
    CascadeBuf I__1366 (
            .O(N__10913),
            .I(N__10907));
    CascadeBuf I__1365 (
            .O(N__10910),
            .I(N__10904));
    CascadeMux I__1364 (
            .O(N__10907),
            .I(N__10901));
    CascadeMux I__1363 (
            .O(N__10904),
            .I(N__10898));
    CascadeBuf I__1362 (
            .O(N__10901),
            .I(N__10895));
    CascadeBuf I__1361 (
            .O(N__10898),
            .I(N__10892));
    CascadeMux I__1360 (
            .O(N__10895),
            .I(N__10889));
    CascadeMux I__1359 (
            .O(N__10892),
            .I(N__10886));
    CascadeBuf I__1358 (
            .O(N__10889),
            .I(N__10883));
    CascadeBuf I__1357 (
            .O(N__10886),
            .I(N__10880));
    CascadeMux I__1356 (
            .O(N__10883),
            .I(N__10877));
    CascadeMux I__1355 (
            .O(N__10880),
            .I(N__10874));
    CascadeBuf I__1354 (
            .O(N__10877),
            .I(N__10871));
    CascadeBuf I__1353 (
            .O(N__10874),
            .I(N__10868));
    CascadeMux I__1352 (
            .O(N__10871),
            .I(N__10865));
    CascadeMux I__1351 (
            .O(N__10868),
            .I(N__10862));
    CascadeBuf I__1350 (
            .O(N__10865),
            .I(N__10859));
    CascadeBuf I__1349 (
            .O(N__10862),
            .I(N__10856));
    CascadeMux I__1348 (
            .O(N__10859),
            .I(N__10853));
    CascadeMux I__1347 (
            .O(N__10856),
            .I(N__10850));
    CascadeBuf I__1346 (
            .O(N__10853),
            .I(N__10847));
    CascadeBuf I__1345 (
            .O(N__10850),
            .I(N__10844));
    CascadeMux I__1344 (
            .O(N__10847),
            .I(N__10841));
    CascadeMux I__1343 (
            .O(N__10844),
            .I(N__10838));
    CascadeBuf I__1342 (
            .O(N__10841),
            .I(N__10835));
    CascadeBuf I__1341 (
            .O(N__10838),
            .I(N__10832));
    CascadeMux I__1340 (
            .O(N__10835),
            .I(N__10829));
    CascadeMux I__1339 (
            .O(N__10832),
            .I(N__10826));
    CascadeBuf I__1338 (
            .O(N__10829),
            .I(N__10823));
    CascadeBuf I__1337 (
            .O(N__10826),
            .I(N__10820));
    CascadeMux I__1336 (
            .O(N__10823),
            .I(N__10817));
    CascadeMux I__1335 (
            .O(N__10820),
            .I(N__10814));
    CascadeBuf I__1334 (
            .O(N__10817),
            .I(N__10811));
    CascadeBuf I__1333 (
            .O(N__10814),
            .I(N__10808));
    CascadeMux I__1332 (
            .O(N__10811),
            .I(N__10805));
    CascadeMux I__1331 (
            .O(N__10808),
            .I(N__10802));
    CascadeBuf I__1330 (
            .O(N__10805),
            .I(N__10799));
    CascadeBuf I__1329 (
            .O(N__10802),
            .I(N__10796));
    CascadeMux I__1328 (
            .O(N__10799),
            .I(N__10793));
    CascadeMux I__1327 (
            .O(N__10796),
            .I(N__10790));
    CascadeBuf I__1326 (
            .O(N__10793),
            .I(N__10787));
    CascadeBuf I__1325 (
            .O(N__10790),
            .I(N__10784));
    CascadeMux I__1324 (
            .O(N__10787),
            .I(N__10781));
    CascadeMux I__1323 (
            .O(N__10784),
            .I(N__10778));
    CascadeBuf I__1322 (
            .O(N__10781),
            .I(N__10775));
    CascadeBuf I__1321 (
            .O(N__10778),
            .I(N__10772));
    CascadeMux I__1320 (
            .O(N__10775),
            .I(N__10769));
    CascadeMux I__1319 (
            .O(N__10772),
            .I(N__10766));
    CascadeBuf I__1318 (
            .O(N__10769),
            .I(N__10763));
    CascadeBuf I__1317 (
            .O(N__10766),
            .I(N__10760));
    CascadeMux I__1316 (
            .O(N__10763),
            .I(N__10757));
    CascadeMux I__1315 (
            .O(N__10760),
            .I(N__10754));
    CascadeBuf I__1314 (
            .O(N__10757),
            .I(N__10751));
    InMux I__1313 (
            .O(N__10754),
            .I(N__10748));
    CascadeMux I__1312 (
            .O(N__10751),
            .I(N__10745));
    LocalMux I__1311 (
            .O(N__10748),
            .I(N__10742));
    CascadeBuf I__1310 (
            .O(N__10745),
            .I(N__10739));
    Span4Mux_v I__1309 (
            .O(N__10742),
            .I(N__10736));
    CascadeMux I__1308 (
            .O(N__10739),
            .I(N__10733));
    Span4Mux_v I__1307 (
            .O(N__10736),
            .I(N__10730));
    InMux I__1306 (
            .O(N__10733),
            .I(N__10727));
    Span4Mux_h I__1305 (
            .O(N__10730),
            .I(N__10724));
    LocalMux I__1304 (
            .O(N__10727),
            .I(N__10721));
    Span4Mux_h I__1303 (
            .O(N__10724),
            .I(N__10718));
    Span4Mux_v I__1302 (
            .O(N__10721),
            .I(N__10715));
    Span4Mux_h I__1301 (
            .O(N__10718),
            .I(N__10710));
    Span4Mux_h I__1300 (
            .O(N__10715),
            .I(N__10710));
    Sp12to4 I__1299 (
            .O(N__10710),
            .I(N__10707));
    Odrv12 I__1298 (
            .O(N__10707),
            .I(n25));
    InMux I__1297 (
            .O(N__10704),
            .I(N__10701));
    LocalMux I__1296 (
            .O(N__10701),
            .I(N__10697));
    InMux I__1295 (
            .O(N__10700),
            .I(N__10694));
    Odrv4 I__1294 (
            .O(N__10697),
            .I(\transmit_module.n113 ));
    LocalMux I__1293 (
            .O(N__10694),
            .I(\transmit_module.n113 ));
    InMux I__1292 (
            .O(N__10689),
            .I(N__10686));
    LocalMux I__1291 (
            .O(N__10686),
            .I(\transmit_module.ADDR_Y_COMPONENT_2 ));
    InMux I__1290 (
            .O(N__10683),
            .I(N__10677));
    InMux I__1289 (
            .O(N__10682),
            .I(N__10677));
    LocalMux I__1288 (
            .O(N__10677),
            .I(\transmit_module.n115 ));
    InMux I__1287 (
            .O(N__10674),
            .I(N__10671));
    LocalMux I__1286 (
            .O(N__10671),
            .I(\transmit_module.n142 ));
    CascadeMux I__1285 (
            .O(N__10668),
            .I(\transmit_module.n142_cascade_ ));
    CascadeMux I__1284 (
            .O(N__10665),
            .I(N__10662));
    CascadeBuf I__1283 (
            .O(N__10662),
            .I(N__10659));
    CascadeMux I__1282 (
            .O(N__10659),
            .I(N__10656));
    CascadeBuf I__1281 (
            .O(N__10656),
            .I(N__10652));
    CascadeMux I__1280 (
            .O(N__10655),
            .I(N__10649));
    CascadeMux I__1279 (
            .O(N__10652),
            .I(N__10646));
    CascadeBuf I__1278 (
            .O(N__10649),
            .I(N__10643));
    CascadeBuf I__1277 (
            .O(N__10646),
            .I(N__10640));
    CascadeMux I__1276 (
            .O(N__10643),
            .I(N__10637));
    CascadeMux I__1275 (
            .O(N__10640),
            .I(N__10634));
    CascadeBuf I__1274 (
            .O(N__10637),
            .I(N__10631));
    CascadeBuf I__1273 (
            .O(N__10634),
            .I(N__10628));
    CascadeMux I__1272 (
            .O(N__10631),
            .I(N__10625));
    CascadeMux I__1271 (
            .O(N__10628),
            .I(N__10622));
    CascadeBuf I__1270 (
            .O(N__10625),
            .I(N__10619));
    CascadeBuf I__1269 (
            .O(N__10622),
            .I(N__10616));
    CascadeMux I__1268 (
            .O(N__10619),
            .I(N__10613));
    CascadeMux I__1267 (
            .O(N__10616),
            .I(N__10610));
    CascadeBuf I__1266 (
            .O(N__10613),
            .I(N__10607));
    CascadeBuf I__1265 (
            .O(N__10610),
            .I(N__10604));
    CascadeMux I__1264 (
            .O(N__10607),
            .I(N__10601));
    CascadeMux I__1263 (
            .O(N__10604),
            .I(N__10598));
    CascadeBuf I__1262 (
            .O(N__10601),
            .I(N__10595));
    CascadeBuf I__1261 (
            .O(N__10598),
            .I(N__10592));
    CascadeMux I__1260 (
            .O(N__10595),
            .I(N__10589));
    CascadeMux I__1259 (
            .O(N__10592),
            .I(N__10586));
    CascadeBuf I__1258 (
            .O(N__10589),
            .I(N__10583));
    CascadeBuf I__1257 (
            .O(N__10586),
            .I(N__10580));
    CascadeMux I__1256 (
            .O(N__10583),
            .I(N__10577));
    CascadeMux I__1255 (
            .O(N__10580),
            .I(N__10574));
    CascadeBuf I__1254 (
            .O(N__10577),
            .I(N__10571));
    CascadeBuf I__1253 (
            .O(N__10574),
            .I(N__10568));
    CascadeMux I__1252 (
            .O(N__10571),
            .I(N__10565));
    CascadeMux I__1251 (
            .O(N__10568),
            .I(N__10562));
    CascadeBuf I__1250 (
            .O(N__10565),
            .I(N__10559));
    CascadeBuf I__1249 (
            .O(N__10562),
            .I(N__10556));
    CascadeMux I__1248 (
            .O(N__10559),
            .I(N__10553));
    CascadeMux I__1247 (
            .O(N__10556),
            .I(N__10550));
    CascadeBuf I__1246 (
            .O(N__10553),
            .I(N__10547));
    CascadeBuf I__1245 (
            .O(N__10550),
            .I(N__10544));
    CascadeMux I__1244 (
            .O(N__10547),
            .I(N__10541));
    CascadeMux I__1243 (
            .O(N__10544),
            .I(N__10538));
    CascadeBuf I__1242 (
            .O(N__10541),
            .I(N__10535));
    CascadeBuf I__1241 (
            .O(N__10538),
            .I(N__10532));
    CascadeMux I__1240 (
            .O(N__10535),
            .I(N__10529));
    CascadeMux I__1239 (
            .O(N__10532),
            .I(N__10526));
    CascadeBuf I__1238 (
            .O(N__10529),
            .I(N__10523));
    CascadeBuf I__1237 (
            .O(N__10526),
            .I(N__10520));
    CascadeMux I__1236 (
            .O(N__10523),
            .I(N__10517));
    CascadeMux I__1235 (
            .O(N__10520),
            .I(N__10514));
    CascadeBuf I__1234 (
            .O(N__10517),
            .I(N__10511));
    CascadeBuf I__1233 (
            .O(N__10514),
            .I(N__10508));
    CascadeMux I__1232 (
            .O(N__10511),
            .I(N__10505));
    CascadeMux I__1231 (
            .O(N__10508),
            .I(N__10502));
    CascadeBuf I__1230 (
            .O(N__10505),
            .I(N__10499));
    CascadeBuf I__1229 (
            .O(N__10502),
            .I(N__10496));
    CascadeMux I__1228 (
            .O(N__10499),
            .I(N__10493));
    CascadeMux I__1227 (
            .O(N__10496),
            .I(N__10490));
    CascadeBuf I__1226 (
            .O(N__10493),
            .I(N__10487));
    InMux I__1225 (
            .O(N__10490),
            .I(N__10484));
    CascadeMux I__1224 (
            .O(N__10487),
            .I(N__10481));
    LocalMux I__1223 (
            .O(N__10484),
            .I(N__10478));
    CascadeBuf I__1222 (
            .O(N__10481),
            .I(N__10475));
    Span4Mux_v I__1221 (
            .O(N__10478),
            .I(N__10472));
    CascadeMux I__1220 (
            .O(N__10475),
            .I(N__10469));
    Span4Mux_v I__1219 (
            .O(N__10472),
            .I(N__10466));
    InMux I__1218 (
            .O(N__10469),
            .I(N__10463));
    Span4Mux_h I__1217 (
            .O(N__10466),
            .I(N__10460));
    LocalMux I__1216 (
            .O(N__10463),
            .I(N__10457));
    Span4Mux_h I__1215 (
            .O(N__10460),
            .I(N__10454));
    Span4Mux_v I__1214 (
            .O(N__10457),
            .I(N__10451));
    Span4Mux_h I__1213 (
            .O(N__10454),
            .I(N__10446));
    Span4Mux_h I__1212 (
            .O(N__10451),
            .I(N__10446));
    Sp12to4 I__1211 (
            .O(N__10446),
            .I(N__10443));
    Odrv12 I__1210 (
            .O(N__10443),
            .I(n23));
    InMux I__1209 (
            .O(N__10440),
            .I(N__10436));
    InMux I__1208 (
            .O(N__10439),
            .I(N__10433));
    LocalMux I__1207 (
            .O(N__10436),
            .I(\transmit_module.n111 ));
    LocalMux I__1206 (
            .O(N__10433),
            .I(\transmit_module.n111 ));
    InMux I__1205 (
            .O(N__10428),
            .I(N__10425));
    LocalMux I__1204 (
            .O(N__10425),
            .I(\transmit_module.n138 ));
    CascadeMux I__1203 (
            .O(N__10422),
            .I(\transmit_module.n138_cascade_ ));
    InMux I__1202 (
            .O(N__10419),
            .I(N__10416));
    LocalMux I__1201 (
            .O(N__10416),
            .I(\transmit_module.n107 ));
    CascadeMux I__1200 (
            .O(N__10413),
            .I(N__10410));
    CascadeBuf I__1199 (
            .O(N__10410),
            .I(N__10407));
    CascadeMux I__1198 (
            .O(N__10407),
            .I(N__10403));
    CascadeMux I__1197 (
            .O(N__10406),
            .I(N__10400));
    CascadeBuf I__1196 (
            .O(N__10403),
            .I(N__10397));
    CascadeBuf I__1195 (
            .O(N__10400),
            .I(N__10394));
    CascadeMux I__1194 (
            .O(N__10397),
            .I(N__10391));
    CascadeMux I__1193 (
            .O(N__10394),
            .I(N__10388));
    CascadeBuf I__1192 (
            .O(N__10391),
            .I(N__10385));
    CascadeBuf I__1191 (
            .O(N__10388),
            .I(N__10382));
    CascadeMux I__1190 (
            .O(N__10385),
            .I(N__10379));
    CascadeMux I__1189 (
            .O(N__10382),
            .I(N__10376));
    CascadeBuf I__1188 (
            .O(N__10379),
            .I(N__10373));
    CascadeBuf I__1187 (
            .O(N__10376),
            .I(N__10370));
    CascadeMux I__1186 (
            .O(N__10373),
            .I(N__10367));
    CascadeMux I__1185 (
            .O(N__10370),
            .I(N__10364));
    CascadeBuf I__1184 (
            .O(N__10367),
            .I(N__10361));
    CascadeBuf I__1183 (
            .O(N__10364),
            .I(N__10358));
    CascadeMux I__1182 (
            .O(N__10361),
            .I(N__10355));
    CascadeMux I__1181 (
            .O(N__10358),
            .I(N__10352));
    CascadeBuf I__1180 (
            .O(N__10355),
            .I(N__10349));
    CascadeBuf I__1179 (
            .O(N__10352),
            .I(N__10346));
    CascadeMux I__1178 (
            .O(N__10349),
            .I(N__10343));
    CascadeMux I__1177 (
            .O(N__10346),
            .I(N__10340));
    CascadeBuf I__1176 (
            .O(N__10343),
            .I(N__10337));
    CascadeBuf I__1175 (
            .O(N__10340),
            .I(N__10334));
    CascadeMux I__1174 (
            .O(N__10337),
            .I(N__10331));
    CascadeMux I__1173 (
            .O(N__10334),
            .I(N__10328));
    CascadeBuf I__1172 (
            .O(N__10331),
            .I(N__10325));
    CascadeBuf I__1171 (
            .O(N__10328),
            .I(N__10322));
    CascadeMux I__1170 (
            .O(N__10325),
            .I(N__10319));
    CascadeMux I__1169 (
            .O(N__10322),
            .I(N__10316));
    CascadeBuf I__1168 (
            .O(N__10319),
            .I(N__10313));
    CascadeBuf I__1167 (
            .O(N__10316),
            .I(N__10310));
    CascadeMux I__1166 (
            .O(N__10313),
            .I(N__10307));
    CascadeMux I__1165 (
            .O(N__10310),
            .I(N__10304));
    CascadeBuf I__1164 (
            .O(N__10307),
            .I(N__10301));
    CascadeBuf I__1163 (
            .O(N__10304),
            .I(N__10298));
    CascadeMux I__1162 (
            .O(N__10301),
            .I(N__10295));
    CascadeMux I__1161 (
            .O(N__10298),
            .I(N__10292));
    CascadeBuf I__1160 (
            .O(N__10295),
            .I(N__10289));
    CascadeBuf I__1159 (
            .O(N__10292),
            .I(N__10286));
    CascadeMux I__1158 (
            .O(N__10289),
            .I(N__10283));
    CascadeMux I__1157 (
            .O(N__10286),
            .I(N__10280));
    CascadeBuf I__1156 (
            .O(N__10283),
            .I(N__10277));
    CascadeBuf I__1155 (
            .O(N__10280),
            .I(N__10274));
    CascadeMux I__1154 (
            .O(N__10277),
            .I(N__10271));
    CascadeMux I__1153 (
            .O(N__10274),
            .I(N__10268));
    CascadeBuf I__1152 (
            .O(N__10271),
            .I(N__10265));
    CascadeBuf I__1151 (
            .O(N__10268),
            .I(N__10262));
    CascadeMux I__1150 (
            .O(N__10265),
            .I(N__10259));
    CascadeMux I__1149 (
            .O(N__10262),
            .I(N__10256));
    CascadeBuf I__1148 (
            .O(N__10259),
            .I(N__10253));
    CascadeBuf I__1147 (
            .O(N__10256),
            .I(N__10250));
    CascadeMux I__1146 (
            .O(N__10253),
            .I(N__10247));
    CascadeMux I__1145 (
            .O(N__10250),
            .I(N__10244));
    CascadeBuf I__1144 (
            .O(N__10247),
            .I(N__10241));
    CascadeBuf I__1143 (
            .O(N__10244),
            .I(N__10238));
    CascadeMux I__1142 (
            .O(N__10241),
            .I(N__10235));
    CascadeMux I__1141 (
            .O(N__10238),
            .I(N__10232));
    InMux I__1140 (
            .O(N__10235),
            .I(N__10229));
    CascadeBuf I__1139 (
            .O(N__10232),
            .I(N__10226));
    LocalMux I__1138 (
            .O(N__10229),
            .I(N__10223));
    CascadeMux I__1137 (
            .O(N__10226),
            .I(N__10220));
    Span4Mux_v I__1136 (
            .O(N__10223),
            .I(N__10217));
    InMux I__1135 (
            .O(N__10220),
            .I(N__10214));
    Span4Mux_v I__1134 (
            .O(N__10217),
            .I(N__10211));
    LocalMux I__1133 (
            .O(N__10214),
            .I(N__10208));
    Span4Mux_v I__1132 (
            .O(N__10211),
            .I(N__10205));
    Span4Mux_v I__1131 (
            .O(N__10208),
            .I(N__10202));
    Span4Mux_h I__1130 (
            .O(N__10205),
            .I(N__10199));
    Span4Mux_v I__1129 (
            .O(N__10202),
            .I(N__10196));
    Span4Mux_h I__1128 (
            .O(N__10199),
            .I(N__10193));
    Span4Mux_v I__1127 (
            .O(N__10196),
            .I(N__10190));
    Span4Mux_h I__1126 (
            .O(N__10193),
            .I(N__10185));
    Span4Mux_h I__1125 (
            .O(N__10190),
            .I(N__10185));
    Odrv4 I__1124 (
            .O(N__10185),
            .I(n19));
    InMux I__1123 (
            .O(N__10182),
            .I(N__10179));
    LocalMux I__1122 (
            .O(N__10179),
            .I(\transmit_module.n146 ));
    CascadeMux I__1121 (
            .O(N__10176),
            .I(\transmit_module.n146_cascade_ ));
    CascadeMux I__1120 (
            .O(N__10173),
            .I(N__10169));
    CascadeMux I__1119 (
            .O(N__10172),
            .I(N__10166));
    CascadeBuf I__1118 (
            .O(N__10169),
            .I(N__10163));
    CascadeBuf I__1117 (
            .O(N__10166),
            .I(N__10160));
    CascadeMux I__1116 (
            .O(N__10163),
            .I(N__10157));
    CascadeMux I__1115 (
            .O(N__10160),
            .I(N__10154));
    CascadeBuf I__1114 (
            .O(N__10157),
            .I(N__10151));
    CascadeBuf I__1113 (
            .O(N__10154),
            .I(N__10148));
    CascadeMux I__1112 (
            .O(N__10151),
            .I(N__10145));
    CascadeMux I__1111 (
            .O(N__10148),
            .I(N__10142));
    CascadeBuf I__1110 (
            .O(N__10145),
            .I(N__10139));
    CascadeBuf I__1109 (
            .O(N__10142),
            .I(N__10136));
    CascadeMux I__1108 (
            .O(N__10139),
            .I(N__10133));
    CascadeMux I__1107 (
            .O(N__10136),
            .I(N__10130));
    CascadeBuf I__1106 (
            .O(N__10133),
            .I(N__10127));
    CascadeBuf I__1105 (
            .O(N__10130),
            .I(N__10124));
    CascadeMux I__1104 (
            .O(N__10127),
            .I(N__10121));
    CascadeMux I__1103 (
            .O(N__10124),
            .I(N__10118));
    CascadeBuf I__1102 (
            .O(N__10121),
            .I(N__10115));
    CascadeBuf I__1101 (
            .O(N__10118),
            .I(N__10112));
    CascadeMux I__1100 (
            .O(N__10115),
            .I(N__10109));
    CascadeMux I__1099 (
            .O(N__10112),
            .I(N__10106));
    CascadeBuf I__1098 (
            .O(N__10109),
            .I(N__10103));
    CascadeBuf I__1097 (
            .O(N__10106),
            .I(N__10100));
    CascadeMux I__1096 (
            .O(N__10103),
            .I(N__10097));
    CascadeMux I__1095 (
            .O(N__10100),
            .I(N__10094));
    CascadeBuf I__1094 (
            .O(N__10097),
            .I(N__10091));
    CascadeBuf I__1093 (
            .O(N__10094),
            .I(N__10088));
    CascadeMux I__1092 (
            .O(N__10091),
            .I(N__10085));
    CascadeMux I__1091 (
            .O(N__10088),
            .I(N__10082));
    CascadeBuf I__1090 (
            .O(N__10085),
            .I(N__10079));
    CascadeBuf I__1089 (
            .O(N__10082),
            .I(N__10076));
    CascadeMux I__1088 (
            .O(N__10079),
            .I(N__10073));
    CascadeMux I__1087 (
            .O(N__10076),
            .I(N__10070));
    CascadeBuf I__1086 (
            .O(N__10073),
            .I(N__10067));
    CascadeBuf I__1085 (
            .O(N__10070),
            .I(N__10064));
    CascadeMux I__1084 (
            .O(N__10067),
            .I(N__10061));
    CascadeMux I__1083 (
            .O(N__10064),
            .I(N__10058));
    CascadeBuf I__1082 (
            .O(N__10061),
            .I(N__10055));
    CascadeBuf I__1081 (
            .O(N__10058),
            .I(N__10052));
    CascadeMux I__1080 (
            .O(N__10055),
            .I(N__10049));
    CascadeMux I__1079 (
            .O(N__10052),
            .I(N__10046));
    CascadeBuf I__1078 (
            .O(N__10049),
            .I(N__10043));
    CascadeBuf I__1077 (
            .O(N__10046),
            .I(N__10040));
    CascadeMux I__1076 (
            .O(N__10043),
            .I(N__10037));
    CascadeMux I__1075 (
            .O(N__10040),
            .I(N__10034));
    CascadeBuf I__1074 (
            .O(N__10037),
            .I(N__10031));
    CascadeBuf I__1073 (
            .O(N__10034),
            .I(N__10028));
    CascadeMux I__1072 (
            .O(N__10031),
            .I(N__10025));
    CascadeMux I__1071 (
            .O(N__10028),
            .I(N__10022));
    CascadeBuf I__1070 (
            .O(N__10025),
            .I(N__10019));
    CascadeBuf I__1069 (
            .O(N__10022),
            .I(N__10016));
    CascadeMux I__1068 (
            .O(N__10019),
            .I(N__10013));
    CascadeMux I__1067 (
            .O(N__10016),
            .I(N__10010));
    CascadeBuf I__1066 (
            .O(N__10013),
            .I(N__10007));
    CascadeBuf I__1065 (
            .O(N__10010),
            .I(N__10004));
    CascadeMux I__1064 (
            .O(N__10007),
            .I(N__10001));
    CascadeMux I__1063 (
            .O(N__10004),
            .I(N__9998));
    CascadeBuf I__1062 (
            .O(N__10001),
            .I(N__9995));
    CascadeBuf I__1061 (
            .O(N__9998),
            .I(N__9992));
    CascadeMux I__1060 (
            .O(N__9995),
            .I(N__9989));
    CascadeMux I__1059 (
            .O(N__9992),
            .I(N__9986));
    InMux I__1058 (
            .O(N__9989),
            .I(N__9983));
    InMux I__1057 (
            .O(N__9986),
            .I(N__9980));
    LocalMux I__1056 (
            .O(N__9983),
            .I(N__9977));
    LocalMux I__1055 (
            .O(N__9980),
            .I(N__9974));
    Span4Mux_v I__1054 (
            .O(N__9977),
            .I(N__9971));
    Sp12to4 I__1053 (
            .O(N__9974),
            .I(N__9968));
    Span4Mux_v I__1052 (
            .O(N__9971),
            .I(N__9965));
    Span12Mux_s10_v I__1051 (
            .O(N__9968),
            .I(N__9962));
    Span4Mux_h I__1050 (
            .O(N__9965),
            .I(N__9959));
    Span12Mux_h I__1049 (
            .O(N__9962),
            .I(N__9954));
    Sp12to4 I__1048 (
            .O(N__9959),
            .I(N__9954));
    Odrv12 I__1047 (
            .O(N__9954),
            .I(n27));
    CascadeMux I__1046 (
            .O(N__9951),
            .I(\transmit_module.n107_cascade_ ));
    CascadeMux I__1045 (
            .O(N__9948),
            .I(\transmit_module.n145_cascade_ ));
    InMux I__1044 (
            .O(N__9945),
            .I(N__9942));
    LocalMux I__1043 (
            .O(N__9942),
            .I(\transmit_module.video_signal_controller.n7 ));
    InMux I__1042 (
            .O(N__9939),
            .I(N__9934));
    InMux I__1041 (
            .O(N__9938),
            .I(N__9931));
    InMux I__1040 (
            .O(N__9937),
            .I(N__9928));
    LocalMux I__1039 (
            .O(N__9934),
            .I(N__9925));
    LocalMux I__1038 (
            .O(N__9931),
            .I(N__9922));
    LocalMux I__1037 (
            .O(N__9928),
            .I(\transmit_module.video_signal_controller.VGA_X_0 ));
    Odrv4 I__1036 (
            .O(N__9925),
            .I(\transmit_module.video_signal_controller.VGA_X_0 ));
    Odrv4 I__1035 (
            .O(N__9922),
            .I(\transmit_module.video_signal_controller.VGA_X_0 ));
    CEMux I__1034 (
            .O(N__9915),
            .I(N__9909));
    CEMux I__1033 (
            .O(N__9914),
            .I(N__9905));
    CEMux I__1032 (
            .O(N__9913),
            .I(N__9901));
    CEMux I__1031 (
            .O(N__9912),
            .I(N__9896));
    LocalMux I__1030 (
            .O(N__9909),
            .I(N__9891));
    CEMux I__1029 (
            .O(N__9908),
            .I(N__9888));
    LocalMux I__1028 (
            .O(N__9905),
            .I(N__9885));
    CEMux I__1027 (
            .O(N__9904),
            .I(N__9882));
    LocalMux I__1026 (
            .O(N__9901),
            .I(N__9879));
    CEMux I__1025 (
            .O(N__9900),
            .I(N__9876));
    CEMux I__1024 (
            .O(N__9899),
            .I(N__9873));
    LocalMux I__1023 (
            .O(N__9896),
            .I(N__9869));
    CEMux I__1022 (
            .O(N__9895),
            .I(N__9866));
    CEMux I__1021 (
            .O(N__9894),
            .I(N__9863));
    Span4Mux_v I__1020 (
            .O(N__9891),
            .I(N__9854));
    LocalMux I__1019 (
            .O(N__9888),
            .I(N__9854));
    Span4Mux_v I__1018 (
            .O(N__9885),
            .I(N__9854));
    LocalMux I__1017 (
            .O(N__9882),
            .I(N__9854));
    Span4Mux_v I__1016 (
            .O(N__9879),
            .I(N__9847));
    LocalMux I__1015 (
            .O(N__9876),
            .I(N__9847));
    LocalMux I__1014 (
            .O(N__9873),
            .I(N__9847));
    CEMux I__1013 (
            .O(N__9872),
            .I(N__9844));
    Span4Mux_v I__1012 (
            .O(N__9869),
            .I(N__9837));
    LocalMux I__1011 (
            .O(N__9866),
            .I(N__9837));
    LocalMux I__1010 (
            .O(N__9863),
            .I(N__9837));
    Span4Mux_v I__1009 (
            .O(N__9854),
            .I(N__9834));
    Span4Mux_h I__1008 (
            .O(N__9847),
            .I(N__9831));
    LocalMux I__1007 (
            .O(N__9844),
            .I(N__9828));
    Span4Mux_h I__1006 (
            .O(N__9837),
            .I(N__9825));
    Odrv4 I__1005 (
            .O(N__9834),
            .I(\transmit_module.n3680 ));
    Odrv4 I__1004 (
            .O(N__9831),
            .I(\transmit_module.n3680 ));
    Odrv12 I__1003 (
            .O(N__9828),
            .I(\transmit_module.n3680 ));
    Odrv4 I__1002 (
            .O(N__9825),
            .I(\transmit_module.n3680 ));
    CascadeMux I__1001 (
            .O(N__9816),
            .I(N__9812));
    InMux I__1000 (
            .O(N__9815),
            .I(N__9807));
    InMux I__999 (
            .O(N__9812),
            .I(N__9804));
    InMux I__998 (
            .O(N__9811),
            .I(N__9801));
    InMux I__997 (
            .O(N__9810),
            .I(N__9798));
    LocalMux I__996 (
            .O(N__9807),
            .I(N__9791));
    LocalMux I__995 (
            .O(N__9804),
            .I(N__9791));
    LocalMux I__994 (
            .O(N__9801),
            .I(N__9791));
    LocalMux I__993 (
            .O(N__9798),
            .I(\transmit_module.video_signal_controller.VGA_X_4 ));
    Odrv4 I__992 (
            .O(N__9791),
            .I(\transmit_module.video_signal_controller.VGA_X_4 ));
    CascadeMux I__991 (
            .O(N__9786),
            .I(N__9782));
    InMux I__990 (
            .O(N__9785),
            .I(N__9775));
    InMux I__989 (
            .O(N__9782),
            .I(N__9775));
    InMux I__988 (
            .O(N__9781),
            .I(N__9772));
    InMux I__987 (
            .O(N__9780),
            .I(N__9769));
    LocalMux I__986 (
            .O(N__9775),
            .I(N__9764));
    LocalMux I__985 (
            .O(N__9772),
            .I(N__9764));
    LocalMux I__984 (
            .O(N__9769),
            .I(\transmit_module.video_signal_controller.VGA_X_3 ));
    Odrv4 I__983 (
            .O(N__9764),
            .I(\transmit_module.video_signal_controller.VGA_X_3 ));
    InMux I__982 (
            .O(N__9759),
            .I(N__9751));
    InMux I__981 (
            .O(N__9758),
            .I(N__9751));
    InMux I__980 (
            .O(N__9757),
            .I(N__9748));
    InMux I__979 (
            .O(N__9756),
            .I(N__9745));
    LocalMux I__978 (
            .O(N__9751),
            .I(N__9740));
    LocalMux I__977 (
            .O(N__9748),
            .I(N__9740));
    LocalMux I__976 (
            .O(N__9745),
            .I(\transmit_module.video_signal_controller.VGA_X_5 ));
    Odrv4 I__975 (
            .O(N__9740),
            .I(\transmit_module.video_signal_controller.VGA_X_5 ));
    InMux I__974 (
            .O(N__9735),
            .I(N__9727));
    InMux I__973 (
            .O(N__9734),
            .I(N__9727));
    InMux I__972 (
            .O(N__9733),
            .I(N__9724));
    InMux I__971 (
            .O(N__9732),
            .I(N__9721));
    LocalMux I__970 (
            .O(N__9727),
            .I(N__9716));
    LocalMux I__969 (
            .O(N__9724),
            .I(N__9716));
    LocalMux I__968 (
            .O(N__9721),
            .I(\transmit_module.video_signal_controller.VGA_X_6 ));
    Odrv4 I__967 (
            .O(N__9716),
            .I(\transmit_module.video_signal_controller.VGA_X_6 ));
    InMux I__966 (
            .O(N__9711),
            .I(N__9706));
    InMux I__965 (
            .O(N__9710),
            .I(N__9703));
    InMux I__964 (
            .O(N__9709),
            .I(N__9700));
    LocalMux I__963 (
            .O(N__9706),
            .I(N__9695));
    LocalMux I__962 (
            .O(N__9703),
            .I(N__9695));
    LocalMux I__961 (
            .O(N__9700),
            .I(\transmit_module.video_signal_controller.VGA_X_7 ));
    Odrv4 I__960 (
            .O(N__9695),
            .I(\transmit_module.video_signal_controller.VGA_X_7 ));
    CascadeMux I__959 (
            .O(N__9690),
            .I(\transmit_module.video_signal_controller.n2014_cascade_ ));
    InMux I__958 (
            .O(N__9687),
            .I(N__9681));
    InMux I__957 (
            .O(N__9686),
            .I(N__9678));
    InMux I__956 (
            .O(N__9685),
            .I(N__9675));
    InMux I__955 (
            .O(N__9684),
            .I(N__9672));
    LocalMux I__954 (
            .O(N__9681),
            .I(N__9667));
    LocalMux I__953 (
            .O(N__9678),
            .I(N__9667));
    LocalMux I__952 (
            .O(N__9675),
            .I(\transmit_module.video_signal_controller.VGA_X_2 ));
    LocalMux I__951 (
            .O(N__9672),
            .I(\transmit_module.video_signal_controller.VGA_X_2 ));
    Odrv4 I__950 (
            .O(N__9667),
            .I(\transmit_module.video_signal_controller.VGA_X_2 ));
    InMux I__949 (
            .O(N__9660),
            .I(N__9656));
    InMux I__948 (
            .O(N__9659),
            .I(N__9651));
    LocalMux I__947 (
            .O(N__9656),
            .I(N__9648));
    InMux I__946 (
            .O(N__9655),
            .I(N__9645));
    InMux I__945 (
            .O(N__9654),
            .I(N__9642));
    LocalMux I__944 (
            .O(N__9651),
            .I(N__9639));
    Odrv4 I__943 (
            .O(N__9648),
            .I(\transmit_module.video_signal_controller.VGA_X_1 ));
    LocalMux I__942 (
            .O(N__9645),
            .I(\transmit_module.video_signal_controller.VGA_X_1 ));
    LocalMux I__941 (
            .O(N__9642),
            .I(\transmit_module.video_signal_controller.VGA_X_1 ));
    Odrv4 I__940 (
            .O(N__9639),
            .I(\transmit_module.video_signal_controller.VGA_X_1 ));
    InMux I__939 (
            .O(N__9630),
            .I(N__9627));
    LocalMux I__938 (
            .O(N__9627),
            .I(\transmit_module.video_signal_controller.n3676 ));
    InMux I__937 (
            .O(N__9624),
            .I(\transmit_module.video_signal_controller.n3193 ));
    InMux I__936 (
            .O(N__9621),
            .I(\transmit_module.video_signal_controller.n3194 ));
    InMux I__935 (
            .O(N__9618),
            .I(\transmit_module.video_signal_controller.n3195 ));
    InMux I__934 (
            .O(N__9615),
            .I(\transmit_module.video_signal_controller.n3196 ));
    InMux I__933 (
            .O(N__9612),
            .I(\transmit_module.video_signal_controller.n3197 ));
    InMux I__932 (
            .O(N__9609),
            .I(bfn_13_13_0_));
    InMux I__931 (
            .O(N__9606),
            .I(\transmit_module.video_signal_controller.n3199 ));
    InMux I__930 (
            .O(N__9603),
            .I(\transmit_module.video_signal_controller.n3200 ));
    InMux I__929 (
            .O(N__9600),
            .I(\transmit_module.video_signal_controller.n3201 ));
    SRMux I__928 (
            .O(N__9597),
            .I(N__9594));
    LocalMux I__927 (
            .O(N__9594),
            .I(N__9590));
    SRMux I__926 (
            .O(N__9593),
            .I(N__9587));
    Span4Mux_v I__925 (
            .O(N__9590),
            .I(N__9582));
    LocalMux I__924 (
            .O(N__9587),
            .I(N__9582));
    Odrv4 I__923 (
            .O(N__9582),
            .I(\transmit_module.video_signal_controller.n2395 ));
    InMux I__922 (
            .O(N__9579),
            .I(N__9576));
    LocalMux I__921 (
            .O(N__9576),
            .I(\transmit_module.Y_DELTA_PATTERN_17 ));
    InMux I__920 (
            .O(N__9573),
            .I(N__9570));
    LocalMux I__919 (
            .O(N__9570),
            .I(\transmit_module.Y_DELTA_PATTERN_16 ));
    InMux I__918 (
            .O(N__9567),
            .I(N__9564));
    LocalMux I__917 (
            .O(N__9564),
            .I(\transmit_module.Y_DELTA_PATTERN_13 ));
    InMux I__916 (
            .O(N__9561),
            .I(N__9558));
    LocalMux I__915 (
            .O(N__9558),
            .I(\transmit_module.Y_DELTA_PATTERN_15 ));
    InMux I__914 (
            .O(N__9555),
            .I(N__9552));
    LocalMux I__913 (
            .O(N__9552),
            .I(\transmit_module.Y_DELTA_PATTERN_14 ));
    InMux I__912 (
            .O(N__9549),
            .I(N__9546));
    LocalMux I__911 (
            .O(N__9546),
            .I(\transmit_module.Y_DELTA_PATTERN_18 ));
    InMux I__910 (
            .O(N__9543),
            .I(N__9540));
    LocalMux I__909 (
            .O(N__9540),
            .I(N__9537));
    Odrv4 I__908 (
            .O(N__9537),
            .I(\tvp_video_buffer.BUFFER_1_4 ));
    InMux I__907 (
            .O(N__9534),
            .I(N__9531));
    LocalMux I__906 (
            .O(N__9531),
            .I(N__9528));
    Span4Mux_s1_v I__905 (
            .O(N__9528),
            .I(N__9525));
    Span4Mux_v I__904 (
            .O(N__9525),
            .I(N__9521));
    InMux I__903 (
            .O(N__9524),
            .I(N__9516));
    Span4Mux_v I__902 (
            .O(N__9521),
            .I(N__9510));
    InMux I__901 (
            .O(N__9520),
            .I(N__9507));
    InMux I__900 (
            .O(N__9519),
            .I(N__9504));
    LocalMux I__899 (
            .O(N__9516),
            .I(N__9500));
    InMux I__898 (
            .O(N__9515),
            .I(N__9497));
    InMux I__897 (
            .O(N__9514),
            .I(N__9494));
    InMux I__896 (
            .O(N__9513),
            .I(N__9491));
    Span4Mux_v I__895 (
            .O(N__9510),
            .I(N__9486));
    LocalMux I__894 (
            .O(N__9507),
            .I(N__9486));
    LocalMux I__893 (
            .O(N__9504),
            .I(N__9483));
    InMux I__892 (
            .O(N__9503),
            .I(N__9480));
    Span12Mux_s9_v I__891 (
            .O(N__9500),
            .I(N__9473));
    LocalMux I__890 (
            .O(N__9497),
            .I(N__9473));
    LocalMux I__889 (
            .O(N__9494),
            .I(N__9473));
    LocalMux I__888 (
            .O(N__9491),
            .I(N__9470));
    Span4Mux_v I__887 (
            .O(N__9486),
            .I(N__9467));
    Span4Mux_v I__886 (
            .O(N__9483),
            .I(N__9462));
    LocalMux I__885 (
            .O(N__9480),
            .I(N__9462));
    Span12Mux_v I__884 (
            .O(N__9473),
            .I(N__9457));
    Span12Mux_s10_v I__883 (
            .O(N__9470),
            .I(N__9457));
    Span4Mux_v I__882 (
            .O(N__9467),
            .I(N__9452));
    Span4Mux_v I__881 (
            .O(N__9462),
            .I(N__9452));
    Span12Mux_h I__880 (
            .O(N__9457),
            .I(N__9449));
    Span4Mux_h I__879 (
            .O(N__9452),
            .I(N__9446));
    Odrv12 I__878 (
            .O(N__9449),
            .I(RX_DATA_2));
    Odrv4 I__877 (
            .O(N__9446),
            .I(RX_DATA_2));
    InMux I__876 (
            .O(N__9441),
            .I(bfn_13_12_0_));
    InMux I__875 (
            .O(N__9438),
            .I(\transmit_module.video_signal_controller.n3191 ));
    InMux I__874 (
            .O(N__9435),
            .I(\transmit_module.video_signal_controller.n3192 ));
    InMux I__873 (
            .O(N__9432),
            .I(N__9429));
    LocalMux I__872 (
            .O(N__9429),
            .I(\line_buffer.n3527 ));
    InMux I__871 (
            .O(N__9426),
            .I(N__9423));
    LocalMux I__870 (
            .O(N__9423),
            .I(TX_DATA_2));
    IoInMux I__869 (
            .O(N__9420),
            .I(N__9416));
    IoInMux I__868 (
            .O(N__9419),
            .I(N__9413));
    LocalMux I__867 (
            .O(N__9416),
            .I(N__9410));
    LocalMux I__866 (
            .O(N__9413),
            .I(N__9407));
    IoSpan4Mux I__865 (
            .O(N__9410),
            .I(N__9404));
    IoSpan4Mux I__864 (
            .O(N__9407),
            .I(N__9401));
    Span4Mux_s2_v I__863 (
            .O(N__9404),
            .I(N__9397));
    Span4Mux_s2_v I__862 (
            .O(N__9401),
            .I(N__9394));
    IoInMux I__861 (
            .O(N__9400),
            .I(N__9391));
    Sp12to4 I__860 (
            .O(N__9397),
            .I(N__9388));
    Sp12to4 I__859 (
            .O(N__9394),
            .I(N__9385));
    LocalMux I__858 (
            .O(N__9391),
            .I(N__9382));
    Span12Mux_s10_v I__857 (
            .O(N__9388),
            .I(N__9379));
    Span12Mux_s10_v I__856 (
            .O(N__9385),
            .I(N__9374));
    Span12Mux_s9_h I__855 (
            .O(N__9382),
            .I(N__9374));
    Odrv12 I__854 (
            .O(N__9379),
            .I(n1816));
    Odrv12 I__853 (
            .O(N__9374),
            .I(n1816));
    InMux I__852 (
            .O(N__9369),
            .I(N__9366));
    LocalMux I__851 (
            .O(N__9366),
            .I(N__9363));
    Span12Mux_h I__850 (
            .O(N__9363),
            .I(N__9360));
    Odrv12 I__849 (
            .O(N__9360),
            .I(\line_buffer.n471 ));
    InMux I__848 (
            .O(N__9357),
            .I(N__9354));
    LocalMux I__847 (
            .O(N__9354),
            .I(N__9351));
    Span4Mux_h I__846 (
            .O(N__9351),
            .I(N__9348));
    Odrv4 I__845 (
            .O(N__9348),
            .I(\line_buffer.n463 ));
    InMux I__844 (
            .O(N__9345),
            .I(N__9342));
    LocalMux I__843 (
            .O(N__9342),
            .I(\tvp_video_buffer.BUFFER_1_3 ));
    InMux I__842 (
            .O(N__9339),
            .I(N__9336));
    LocalMux I__841 (
            .O(N__9336),
            .I(N__9332));
    InMux I__840 (
            .O(N__9335),
            .I(N__9328));
    Span4Mux_v I__839 (
            .O(N__9332),
            .I(N__9325));
    InMux I__838 (
            .O(N__9331),
            .I(N__9322));
    LocalMux I__837 (
            .O(N__9328),
            .I(N__9319));
    Span4Mux_v I__836 (
            .O(N__9325),
            .I(N__9313));
    LocalMux I__835 (
            .O(N__9322),
            .I(N__9313));
    Span4Mux_v I__834 (
            .O(N__9319),
            .I(N__9307));
    InMux I__833 (
            .O(N__9318),
            .I(N__9304));
    Span4Mux_v I__832 (
            .O(N__9313),
            .I(N__9300));
    InMux I__831 (
            .O(N__9312),
            .I(N__9297));
    InMux I__830 (
            .O(N__9311),
            .I(N__9294));
    InMux I__829 (
            .O(N__9310),
            .I(N__9291));
    Span4Mux_v I__828 (
            .O(N__9307),
            .I(N__9286));
    LocalMux I__827 (
            .O(N__9304),
            .I(N__9286));
    InMux I__826 (
            .O(N__9303),
            .I(N__9283));
    Sp12to4 I__825 (
            .O(N__9300),
            .I(N__9276));
    LocalMux I__824 (
            .O(N__9297),
            .I(N__9276));
    LocalMux I__823 (
            .O(N__9294),
            .I(N__9276));
    LocalMux I__822 (
            .O(N__9291),
            .I(N__9273));
    Span4Mux_v I__821 (
            .O(N__9286),
            .I(N__9270));
    LocalMux I__820 (
            .O(N__9283),
            .I(N__9267));
    Span12Mux_v I__819 (
            .O(N__9276),
            .I(N__9262));
    Span12Mux_s9_v I__818 (
            .O(N__9273),
            .I(N__9262));
    Span4Mux_v I__817 (
            .O(N__9270),
            .I(N__9257));
    Span4Mux_h I__816 (
            .O(N__9267),
            .I(N__9257));
    Span12Mux_h I__815 (
            .O(N__9262),
            .I(N__9254));
    Span4Mux_h I__814 (
            .O(N__9257),
            .I(N__9251));
    Odrv12 I__813 (
            .O(N__9254),
            .I(RX_DATA_1));
    Odrv4 I__812 (
            .O(N__9251),
            .I(RX_DATA_1));
    InMux I__811 (
            .O(N__9246),
            .I(N__9243));
    LocalMux I__810 (
            .O(N__9243),
            .I(\tvp_video_buffer.BUFFER_1_7 ));
    IoInMux I__809 (
            .O(N__9240),
            .I(N__9237));
    LocalMux I__808 (
            .O(N__9237),
            .I(N__9234));
    IoSpan4Mux I__807 (
            .O(N__9234),
            .I(N__9231));
    Span4Mux_s2_h I__806 (
            .O(N__9231),
            .I(N__9227));
    InMux I__805 (
            .O(N__9230),
            .I(N__9224));
    Sp12to4 I__804 (
            .O(N__9227),
            .I(N__9221));
    LocalMux I__803 (
            .O(N__9224),
            .I(N__9218));
    Span12Mux_v I__802 (
            .O(N__9221),
            .I(N__9215));
    Span4Mux_h I__801 (
            .O(N__9218),
            .I(N__9212));
    Span12Mux_h I__800 (
            .O(N__9215),
            .I(N__9207));
    Sp12to4 I__799 (
            .O(N__9212),
            .I(N__9207));
    Odrv12 I__798 (
            .O(N__9207),
            .I(DEBUG_c_6_c));
    InMux I__797 (
            .O(N__9204),
            .I(N__9201));
    LocalMux I__796 (
            .O(N__9201),
            .I(\tvp_video_buffer.BUFFER_0_7 ));
    InMux I__795 (
            .O(N__9198),
            .I(N__9195));
    LocalMux I__794 (
            .O(N__9195),
            .I(N__9192));
    Odrv4 I__793 (
            .O(N__9192),
            .I(\tvp_video_buffer.BUFFER_0_4 ));
    InMux I__792 (
            .O(N__9189),
            .I(bfn_12_17_0_));
    InMux I__791 (
            .O(N__9186),
            .I(\transmit_module.video_signal_controller.n3188 ));
    InMux I__790 (
            .O(N__9183),
            .I(\transmit_module.video_signal_controller.n3189 ));
    InMux I__789 (
            .O(N__9180),
            .I(\transmit_module.video_signal_controller.n3190 ));
    InMux I__788 (
            .O(N__9177),
            .I(N__9174));
    LocalMux I__787 (
            .O(N__9174),
            .I(N__9171));
    Odrv4 I__786 (
            .O(N__9171),
            .I(\transmit_module.Y_DELTA_PATTERN_3 ));
    InMux I__785 (
            .O(N__9168),
            .I(N__9165));
    LocalMux I__784 (
            .O(N__9165),
            .I(\transmit_module.Y_DELTA_PATTERN_2 ));
    InMux I__783 (
            .O(N__9162),
            .I(N__9159));
    LocalMux I__782 (
            .O(N__9159),
            .I(\transmit_module.Y_DELTA_PATTERN_1 ));
    InMux I__781 (
            .O(N__9156),
            .I(N__9153));
    LocalMux I__780 (
            .O(N__9153),
            .I(N__9150));
    Span4Mux_v I__779 (
            .O(N__9150),
            .I(N__9147));
    Odrv4 I__778 (
            .O(N__9147),
            .I(\line_buffer.n536 ));
    InMux I__777 (
            .O(N__9144),
            .I(N__9141));
    LocalMux I__776 (
            .O(N__9141),
            .I(N__9138));
    Span4Mux_v I__775 (
            .O(N__9138),
            .I(N__9135));
    Sp12to4 I__774 (
            .O(N__9135),
            .I(N__9132));
    Span12Mux_v I__773 (
            .O(N__9132),
            .I(N__9129));
    Span12Mux_h I__772 (
            .O(N__9129),
            .I(N__9126));
    Odrv12 I__771 (
            .O(N__9126),
            .I(\line_buffer.n528 ));
    InMux I__770 (
            .O(N__9123),
            .I(N__9120));
    LocalMux I__769 (
            .O(N__9120),
            .I(N__9117));
    Odrv4 I__768 (
            .O(N__9117),
            .I(\line_buffer.n3528 ));
    InMux I__767 (
            .O(N__9114),
            .I(N__9111));
    LocalMux I__766 (
            .O(N__9111),
            .I(N__9108));
    Span12Mux_v I__765 (
            .O(N__9108),
            .I(N__9105));
    Odrv12 I__764 (
            .O(N__9105),
            .I(\line_buffer.n563 ));
    InMux I__763 (
            .O(N__9102),
            .I(N__9099));
    LocalMux I__762 (
            .O(N__9099),
            .I(N__9096));
    Span4Mux_v I__761 (
            .O(N__9096),
            .I(N__9093));
    Span4Mux_h I__760 (
            .O(N__9093),
            .I(N__9090));
    Sp12to4 I__759 (
            .O(N__9090),
            .I(N__9087));
    Odrv12 I__758 (
            .O(N__9087),
            .I(\line_buffer.n555 ));
    InMux I__757 (
            .O(N__9084),
            .I(N__9081));
    LocalMux I__756 (
            .O(N__9081),
            .I(N__9078));
    Span4Mux_v I__755 (
            .O(N__9078),
            .I(N__9075));
    Odrv4 I__754 (
            .O(N__9075),
            .I(\line_buffer.n3567 ));
    InMux I__753 (
            .O(N__9072),
            .I(bfn_12_16_0_));
    InMux I__752 (
            .O(N__9069),
            .I(\transmit_module.video_signal_controller.n3180 ));
    InMux I__751 (
            .O(N__9066),
            .I(\transmit_module.video_signal_controller.n3181 ));
    InMux I__750 (
            .O(N__9063),
            .I(\transmit_module.video_signal_controller.n3182 ));
    InMux I__749 (
            .O(N__9060),
            .I(\transmit_module.video_signal_controller.n3183 ));
    InMux I__748 (
            .O(N__9057),
            .I(\transmit_module.video_signal_controller.n3184 ));
    InMux I__747 (
            .O(N__9054),
            .I(\transmit_module.video_signal_controller.n3185 ));
    InMux I__746 (
            .O(N__9051),
            .I(\transmit_module.video_signal_controller.n3186 ));
    InMux I__745 (
            .O(N__9048),
            .I(N__9045));
    LocalMux I__744 (
            .O(N__9045),
            .I(\transmit_module.Y_DELTA_PATTERN_12 ));
    InMux I__743 (
            .O(N__9042),
            .I(N__9039));
    LocalMux I__742 (
            .O(N__9039),
            .I(\transmit_module.Y_DELTA_PATTERN_11 ));
    InMux I__741 (
            .O(N__9036),
            .I(N__9033));
    LocalMux I__740 (
            .O(N__9033),
            .I(\transmit_module.Y_DELTA_PATTERN_10 ));
    InMux I__739 (
            .O(N__9030),
            .I(N__9027));
    LocalMux I__738 (
            .O(N__9027),
            .I(\sync_buffer.BUFFER_0_0 ));
    InMux I__737 (
            .O(N__9024),
            .I(N__9021));
    LocalMux I__736 (
            .O(N__9021),
            .I(\sync_buffer.BUFFER_1_0 ));
    InMux I__735 (
            .O(N__9018),
            .I(N__9015));
    LocalMux I__734 (
            .O(N__9015),
            .I(RX_TX_SYNC_BUFF));
    CascadeMux I__733 (
            .O(N__9012),
            .I(\transmit_module.video_signal_controller.n3479_cascade_ ));
    CascadeMux I__732 (
            .O(N__9009),
            .I(\transmit_module.video_signal_controller.n3475_cascade_ ));
    InMux I__731 (
            .O(N__9006),
            .I(N__9003));
    LocalMux I__730 (
            .O(N__9003),
            .I(\transmit_module.video_signal_controller.n55 ));
    InMux I__729 (
            .O(N__9000),
            .I(N__8997));
    LocalMux I__728 (
            .O(N__8997),
            .I(\transmit_module.Y_DELTA_PATTERN_63 ));
    InMux I__727 (
            .O(N__8994),
            .I(N__8991));
    LocalMux I__726 (
            .O(N__8991),
            .I(\transmit_module.Y_DELTA_PATTERN_62 ));
    InMux I__725 (
            .O(N__8988),
            .I(N__8985));
    LocalMux I__724 (
            .O(N__8985),
            .I(N__8982));
    Span12Mux_v I__723 (
            .O(N__8982),
            .I(N__8979));
    Odrv12 I__722 (
            .O(N__8979),
            .I(\line_buffer.n3569 ));
    InMux I__721 (
            .O(N__8976),
            .I(N__8973));
    LocalMux I__720 (
            .O(N__8973),
            .I(\line_buffer.n3566 ));
    CascadeMux I__719 (
            .O(N__8970),
            .I(\line_buffer.n3599_cascade_ ));
    InMux I__718 (
            .O(N__8967),
            .I(N__8964));
    LocalMux I__717 (
            .O(N__8964),
            .I(N__8961));
    Span4Mux_v I__716 (
            .O(N__8961),
            .I(N__8958));
    Odrv4 I__715 (
            .O(N__8958),
            .I(\line_buffer.n595 ));
    InMux I__714 (
            .O(N__8955),
            .I(N__8952));
    LocalMux I__713 (
            .O(N__8952),
            .I(N__8949));
    Span4Mux_h I__712 (
            .O(N__8949),
            .I(N__8946));
    Span4Mux_v I__711 (
            .O(N__8946),
            .I(N__8943));
    Span4Mux_h I__710 (
            .O(N__8943),
            .I(N__8940));
    Span4Mux_h I__709 (
            .O(N__8940),
            .I(N__8937));
    Span4Mux_h I__708 (
            .O(N__8937),
            .I(N__8934));
    Odrv4 I__707 (
            .O(N__8934),
            .I(\line_buffer.n587 ));
    InMux I__706 (
            .O(N__8931),
            .I(N__8928));
    LocalMux I__705 (
            .O(N__8928),
            .I(\line_buffer.n3570 ));
    InMux I__704 (
            .O(N__8925),
            .I(N__8922));
    LocalMux I__703 (
            .O(N__8922),
            .I(N__8919));
    Span4Mux_h I__702 (
            .O(N__8919),
            .I(N__8916));
    IoSpan4Mux I__701 (
            .O(N__8916),
            .I(N__8913));
    Odrv4 I__700 (
            .O(N__8913),
            .I(TVP_VIDEO_c_3));
    InMux I__699 (
            .O(N__8910),
            .I(N__8907));
    LocalMux I__698 (
            .O(N__8907),
            .I(\tvp_video_buffer.BUFFER_0_3 ));
    InMux I__697 (
            .O(N__8904),
            .I(N__8901));
    LocalMux I__696 (
            .O(N__8901),
            .I(\transmit_module.Y_DELTA_PATTERN_71 ));
    InMux I__695 (
            .O(N__8898),
            .I(N__8895));
    LocalMux I__694 (
            .O(N__8895),
            .I(\transmit_module.Y_DELTA_PATTERN_79 ));
    InMux I__693 (
            .O(N__8892),
            .I(N__8889));
    LocalMux I__692 (
            .O(N__8889),
            .I(\transmit_module.Y_DELTA_PATTERN_78 ));
    InMux I__691 (
            .O(N__8886),
            .I(N__8883));
    LocalMux I__690 (
            .O(N__8883),
            .I(\transmit_module.Y_DELTA_PATTERN_72 ));
    InMux I__689 (
            .O(N__8880),
            .I(N__8877));
    LocalMux I__688 (
            .O(N__8877),
            .I(\transmit_module.Y_DELTA_PATTERN_75 ));
    InMux I__687 (
            .O(N__8874),
            .I(N__8871));
    LocalMux I__686 (
            .O(N__8871),
            .I(\transmit_module.Y_DELTA_PATTERN_53 ));
    InMux I__685 (
            .O(N__8868),
            .I(N__8865));
    LocalMux I__684 (
            .O(N__8865),
            .I(\transmit_module.Y_DELTA_PATTERN_52 ));
    InMux I__683 (
            .O(N__8862),
            .I(N__8859));
    LocalMux I__682 (
            .O(N__8859),
            .I(\transmit_module.Y_DELTA_PATTERN_74 ));
    InMux I__681 (
            .O(N__8856),
            .I(N__8853));
    LocalMux I__680 (
            .O(N__8853),
            .I(\transmit_module.Y_DELTA_PATTERN_73 ));
    InMux I__679 (
            .O(N__8850),
            .I(N__8847));
    LocalMux I__678 (
            .O(N__8847),
            .I(\transmit_module.Y_DELTA_PATTERN_61 ));
    InMux I__677 (
            .O(N__8844),
            .I(N__8841));
    LocalMux I__676 (
            .O(N__8841),
            .I(\transmit_module.Y_DELTA_PATTERN_65 ));
    InMux I__675 (
            .O(N__8838),
            .I(N__8835));
    LocalMux I__674 (
            .O(N__8835),
            .I(\transmit_module.Y_DELTA_PATTERN_64 ));
    InMux I__673 (
            .O(N__8832),
            .I(N__8829));
    LocalMux I__672 (
            .O(N__8829),
            .I(\transmit_module.Y_DELTA_PATTERN_33 ));
    InMux I__671 (
            .O(N__8826),
            .I(N__8823));
    LocalMux I__670 (
            .O(N__8823),
            .I(N__8820));
    Odrv4 I__669 (
            .O(N__8820),
            .I(\transmit_module.Y_DELTA_PATTERN_37 ));
    InMux I__668 (
            .O(N__8817),
            .I(N__8814));
    LocalMux I__667 (
            .O(N__8814),
            .I(\transmit_module.Y_DELTA_PATTERN_36 ));
    InMux I__666 (
            .O(N__8811),
            .I(N__8808));
    LocalMux I__665 (
            .O(N__8808),
            .I(\transmit_module.Y_DELTA_PATTERN_35 ));
    InMux I__664 (
            .O(N__8805),
            .I(N__8802));
    LocalMux I__663 (
            .O(N__8802),
            .I(\transmit_module.Y_DELTA_PATTERN_34 ));
    InMux I__662 (
            .O(N__8799),
            .I(N__8796));
    LocalMux I__661 (
            .O(N__8796),
            .I(\transmit_module.Y_DELTA_PATTERN_81 ));
    InMux I__660 (
            .O(N__8793),
            .I(N__8790));
    LocalMux I__659 (
            .O(N__8790),
            .I(\transmit_module.Y_DELTA_PATTERN_82 ));
    InMux I__658 (
            .O(N__8787),
            .I(N__8784));
    LocalMux I__657 (
            .O(N__8784),
            .I(\transmit_module.Y_DELTA_PATTERN_80 ));
    InMux I__656 (
            .O(N__8781),
            .I(N__8778));
    LocalMux I__655 (
            .O(N__8778),
            .I(\transmit_module.Y_DELTA_PATTERN_51 ));
    InMux I__654 (
            .O(N__8775),
            .I(N__8772));
    LocalMux I__653 (
            .O(N__8772),
            .I(\transmit_module.Y_DELTA_PATTERN_70 ));
    InMux I__652 (
            .O(N__8769),
            .I(N__8766));
    LocalMux I__651 (
            .O(N__8766),
            .I(N__8763));
    Span4Mux_v I__650 (
            .O(N__8763),
            .I(N__8760));
    Sp12to4 I__649 (
            .O(N__8760),
            .I(N__8757));
    Span12Mux_h I__648 (
            .O(N__8757),
            .I(N__8754));
    Odrv12 I__647 (
            .O(N__8754),
            .I(\line_buffer.n466 ));
    InMux I__646 (
            .O(N__8751),
            .I(N__8748));
    LocalMux I__645 (
            .O(N__8748),
            .I(N__8745));
    Span4Mux_v I__644 (
            .O(N__8745),
            .I(N__8742));
    Span4Mux_v I__643 (
            .O(N__8742),
            .I(N__8739));
    Span4Mux_v I__642 (
            .O(N__8739),
            .I(N__8736));
    Odrv4 I__641 (
            .O(N__8736),
            .I(\line_buffer.n458 ));
    InMux I__640 (
            .O(N__8733),
            .I(N__8730));
    LocalMux I__639 (
            .O(N__8730),
            .I(N__8727));
    Span4Mux_v I__638 (
            .O(N__8727),
            .I(N__8724));
    Span4Mux_h I__637 (
            .O(N__8724),
            .I(N__8721));
    Odrv4 I__636 (
            .O(N__8721),
            .I(\line_buffer.n531 ));
    InMux I__635 (
            .O(N__8718),
            .I(N__8715));
    LocalMux I__634 (
            .O(N__8715),
            .I(N__8712));
    Span4Mux_v I__633 (
            .O(N__8712),
            .I(N__8709));
    Span4Mux_h I__632 (
            .O(N__8709),
            .I(N__8706));
    Sp12to4 I__631 (
            .O(N__8706),
            .I(N__8703));
    Odrv12 I__630 (
            .O(N__8703),
            .I(\line_buffer.n523 ));
    InMux I__629 (
            .O(N__8700),
            .I(N__8697));
    LocalMux I__628 (
            .O(N__8697),
            .I(N__8694));
    Odrv12 I__627 (
            .O(N__8694),
            .I(TVP_VIDEO_c_4));
    InMux I__626 (
            .O(N__8691),
            .I(N__8688));
    LocalMux I__625 (
            .O(N__8688),
            .I(\transmit_module.Y_DELTA_PATTERN_9 ));
    InMux I__624 (
            .O(N__8685),
            .I(N__8682));
    LocalMux I__623 (
            .O(N__8682),
            .I(\transmit_module.Y_DELTA_PATTERN_29 ));
    InMux I__622 (
            .O(N__8679),
            .I(N__8676));
    LocalMux I__621 (
            .O(N__8676),
            .I(\transmit_module.Y_DELTA_PATTERN_30 ));
    InMux I__620 (
            .O(N__8673),
            .I(N__8670));
    LocalMux I__619 (
            .O(N__8670),
            .I(\transmit_module.Y_DELTA_PATTERN_32 ));
    InMux I__618 (
            .O(N__8667),
            .I(N__8664));
    LocalMux I__617 (
            .O(N__8664),
            .I(\transmit_module.Y_DELTA_PATTERN_31 ));
    InMux I__616 (
            .O(N__8661),
            .I(N__8658));
    LocalMux I__615 (
            .O(N__8658),
            .I(\transmit_module.Y_DELTA_PATTERN_66 ));
    InMux I__614 (
            .O(N__8655),
            .I(N__8652));
    LocalMux I__613 (
            .O(N__8652),
            .I(\transmit_module.Y_DELTA_PATTERN_44 ));
    InMux I__612 (
            .O(N__8649),
            .I(N__8646));
    LocalMux I__611 (
            .O(N__8646),
            .I(\transmit_module.Y_DELTA_PATTERN_43 ));
    InMux I__610 (
            .O(N__8643),
            .I(N__8640));
    LocalMux I__609 (
            .O(N__8640),
            .I(\transmit_module.Y_DELTA_PATTERN_42 ));
    InMux I__608 (
            .O(N__8637),
            .I(N__8634));
    LocalMux I__607 (
            .O(N__8634),
            .I(\transmit_module.Y_DELTA_PATTERN_41 ));
    InMux I__606 (
            .O(N__8631),
            .I(N__8628));
    LocalMux I__605 (
            .O(N__8628),
            .I(\transmit_module.Y_DELTA_PATTERN_40 ));
    InMux I__604 (
            .O(N__8625),
            .I(N__8622));
    LocalMux I__603 (
            .O(N__8622),
            .I(\transmit_module.Y_DELTA_PATTERN_60 ));
    InMux I__602 (
            .O(N__8619),
            .I(N__8616));
    LocalMux I__601 (
            .O(N__8616),
            .I(N__8613));
    Odrv12 I__600 (
            .O(N__8613),
            .I(\transmit_module.Y_DELTA_PATTERN_7 ));
    InMux I__599 (
            .O(N__8610),
            .I(N__8607));
    LocalMux I__598 (
            .O(N__8607),
            .I(N__8604));
    Odrv4 I__597 (
            .O(N__8604),
            .I(\transmit_module.Y_DELTA_PATTERN_6 ));
    InMux I__596 (
            .O(N__8601),
            .I(N__8598));
    LocalMux I__595 (
            .O(N__8598),
            .I(\transmit_module.Y_DELTA_PATTERN_5 ));
    InMux I__594 (
            .O(N__8595),
            .I(N__8592));
    LocalMux I__593 (
            .O(N__8592),
            .I(\transmit_module.Y_DELTA_PATTERN_4 ));
    InMux I__592 (
            .O(N__8589),
            .I(N__8586));
    LocalMux I__591 (
            .O(N__8586),
            .I(\transmit_module.Y_DELTA_PATTERN_50 ));
    InMux I__590 (
            .O(N__8583),
            .I(N__8580));
    LocalMux I__589 (
            .O(N__8580),
            .I(\transmit_module.Y_DELTA_PATTERN_49 ));
    InMux I__588 (
            .O(N__8577),
            .I(N__8574));
    LocalMux I__587 (
            .O(N__8574),
            .I(\transmit_module.Y_DELTA_PATTERN_54 ));
    InMux I__586 (
            .O(N__8571),
            .I(N__8568));
    LocalMux I__585 (
            .O(N__8568),
            .I(\transmit_module.Y_DELTA_PATTERN_67 ));
    InMux I__584 (
            .O(N__8565),
            .I(N__8562));
    LocalMux I__583 (
            .O(N__8562),
            .I(\transmit_module.Y_DELTA_PATTERN_77 ));
    InMux I__582 (
            .O(N__8559),
            .I(N__8556));
    LocalMux I__581 (
            .O(N__8556),
            .I(\transmit_module.Y_DELTA_PATTERN_69 ));
    InMux I__580 (
            .O(N__8553),
            .I(N__8550));
    LocalMux I__579 (
            .O(N__8550),
            .I(\transmit_module.Y_DELTA_PATTERN_68 ));
    InMux I__578 (
            .O(N__8547),
            .I(N__8544));
    LocalMux I__577 (
            .O(N__8544),
            .I(\transmit_module.Y_DELTA_PATTERN_76 ));
    InMux I__576 (
            .O(N__8541),
            .I(N__8538));
    LocalMux I__575 (
            .O(N__8538),
            .I(N__8535));
    Span4Mux_v I__574 (
            .O(N__8535),
            .I(N__8532));
    Odrv4 I__573 (
            .O(N__8532),
            .I(\line_buffer.n600 ));
    InMux I__572 (
            .O(N__8529),
            .I(N__8526));
    LocalMux I__571 (
            .O(N__8526),
            .I(N__8523));
    Span4Mux_v I__570 (
            .O(N__8523),
            .I(N__8520));
    Odrv4 I__569 (
            .O(N__8520),
            .I(\line_buffer.n592 ));
    InMux I__568 (
            .O(N__8517),
            .I(N__8514));
    LocalMux I__567 (
            .O(N__8514),
            .I(\transmit_module.Y_DELTA_PATTERN_28 ));
    InMux I__566 (
            .O(N__8511),
            .I(N__8508));
    LocalMux I__565 (
            .O(N__8508),
            .I(\transmit_module.Y_DELTA_PATTERN_27 ));
    InMux I__564 (
            .O(N__8505),
            .I(N__8502));
    LocalMux I__563 (
            .O(N__8502),
            .I(\transmit_module.Y_DELTA_PATTERN_8 ));
    InMux I__562 (
            .O(N__8499),
            .I(N__8496));
    LocalMux I__561 (
            .O(N__8496),
            .I(\transmit_module.Y_DELTA_PATTERN_48 ));
    InMux I__560 (
            .O(N__8493),
            .I(N__8490));
    LocalMux I__559 (
            .O(N__8490),
            .I(\transmit_module.Y_DELTA_PATTERN_47 ));
    InMux I__558 (
            .O(N__8487),
            .I(N__8484));
    LocalMux I__557 (
            .O(N__8484),
            .I(\transmit_module.Y_DELTA_PATTERN_55 ));
    InMux I__556 (
            .O(N__8481),
            .I(N__8478));
    LocalMux I__555 (
            .O(N__8478),
            .I(\transmit_module.Y_DELTA_PATTERN_46 ));
    InMux I__554 (
            .O(N__8475),
            .I(N__8472));
    LocalMux I__553 (
            .O(N__8472),
            .I(\transmit_module.Y_DELTA_PATTERN_58 ));
    InMux I__552 (
            .O(N__8469),
            .I(N__8466));
    LocalMux I__551 (
            .O(N__8466),
            .I(\transmit_module.Y_DELTA_PATTERN_59 ));
    InMux I__550 (
            .O(N__8463),
            .I(N__8460));
    LocalMux I__549 (
            .O(N__8460),
            .I(\transmit_module.Y_DELTA_PATTERN_57 ));
    InMux I__548 (
            .O(N__8457),
            .I(N__8454));
    LocalMux I__547 (
            .O(N__8454),
            .I(\transmit_module.Y_DELTA_PATTERN_56 ));
    InMux I__546 (
            .O(N__8451),
            .I(N__8448));
    LocalMux I__545 (
            .O(N__8448),
            .I(N__8445));
    Odrv4 I__544 (
            .O(N__8445),
            .I(\transmit_module.Y_DELTA_PATTERN_39 ));
    InMux I__543 (
            .O(N__8442),
            .I(N__8439));
    LocalMux I__542 (
            .O(N__8439),
            .I(\transmit_module.Y_DELTA_PATTERN_45 ));
    InMux I__541 (
            .O(N__8436),
            .I(N__8433));
    LocalMux I__540 (
            .O(N__8433),
            .I(N__8430));
    Span4Mux_v I__539 (
            .O(N__8430),
            .I(N__8427));
    Odrv4 I__538 (
            .O(N__8427),
            .I(\line_buffer.n599 ));
    InMux I__537 (
            .O(N__8424),
            .I(N__8421));
    LocalMux I__536 (
            .O(N__8421),
            .I(N__8418));
    Span4Mux_v I__535 (
            .O(N__8418),
            .I(N__8415));
    Odrv4 I__534 (
            .O(N__8415),
            .I(\line_buffer.n591 ));
    InMux I__533 (
            .O(N__8412),
            .I(N__8409));
    LocalMux I__532 (
            .O(N__8409),
            .I(\transmit_module.Y_DELTA_PATTERN_38 ));
    defparam IN_MUX_bfv_13_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_12_0_));
    defparam IN_MUX_bfv_13_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_13_0_ (
            .carryinitin(\transmit_module.video_signal_controller.n3198 ),
            .carryinitout(bfn_13_13_0_));
    defparam IN_MUX_bfv_12_16_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_16_0_));
    defparam IN_MUX_bfv_12_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_17_0_ (
            .carryinitin(\transmit_module.video_signal_controller.n3187 ),
            .carryinitout(bfn_12_17_0_));
    defparam IN_MUX_bfv_14_15_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_15_0_));
    defparam IN_MUX_bfv_14_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_16_0_ (
            .carryinitin(\transmit_module.n3166 ),
            .carryinitout(bfn_14_16_0_));
    defparam IN_MUX_bfv_17_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_9_0_));
    defparam IN_MUX_bfv_17_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_10_0_ (
            .carryinitin(\receive_module.rx_counter.n3179 ),
            .carryinitout(bfn_17_10_0_));
    defparam IN_MUX_bfv_15_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_10_0_));
    defparam IN_MUX_bfv_15_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_11_0_ (
            .carryinitin(\receive_module.rx_counter.n3214 ),
            .carryinitout(bfn_15_11_0_));
    defparam IN_MUX_bfv_16_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_12_0_));
    defparam IN_MUX_bfv_15_16_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_16_0_));
    defparam IN_MUX_bfv_15_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_17_0_ (
            .carryinitin(\receive_module.n3153 ),
            .carryinitout(bfn_15_17_0_));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \transmit_module.Y_DELTA_PATTERN_i26_LC_9_11_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i26_LC_9_11_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i26_LC_9_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i26_LC_9_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8511),
            .lcout(\transmit_module.Y_DELTA_PATTERN_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24301),
            .ce(N__20514),
            .sr(N__23331));
    defparam \transmit_module.Y_DELTA_PATTERN_i37_LC_9_12_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i37_LC_9_12_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i37_LC_9_12_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i37_LC_9_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8412),
            .lcout(\transmit_module.Y_DELTA_PATTERN_37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24335),
            .ce(N__9912),
            .sr(N__23335));
    defparam \transmit_module.Y_DELTA_PATTERN_i46_LC_9_13_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i46_LC_9_13_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i46_LC_9_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i46_LC_9_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8493),
            .lcout(\transmit_module.Y_DELTA_PATTERN_46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24312),
            .ce(N__9900),
            .sr(N__23274));
    defparam \transmit_module.Y_DELTA_PATTERN_i38_LC_9_13_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i38_LC_9_13_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i38_LC_9_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i38_LC_9_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8451),
            .lcout(\transmit_module.Y_DELTA_PATTERN_38 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24312),
            .ce(N__9900),
            .sr(N__23274));
    defparam \transmit_module.Y_DELTA_PATTERN_i54_LC_9_14_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i54_LC_9_14_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i54_LC_9_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i54_LC_9_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8487),
            .lcout(\transmit_module.Y_DELTA_PATTERN_54 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24299),
            .ce(N__9895),
            .sr(N__23303));
    defparam \transmit_module.Y_DELTA_PATTERN_i55_LC_9_14_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i55_LC_9_14_2 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i55_LC_9_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i55_LC_9_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8457),
            .lcout(\transmit_module.Y_DELTA_PATTERN_55 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24299),
            .ce(N__9895),
            .sr(N__23303));
    defparam \transmit_module.Y_DELTA_PATTERN_i45_LC_9_14_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i45_LC_9_14_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i45_LC_9_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i45_LC_9_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8481),
            .lcout(\transmit_module.Y_DELTA_PATTERN_45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24299),
            .ce(N__9895),
            .sr(N__23303));
    defparam \transmit_module.Y_DELTA_PATTERN_i58_LC_9_14_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i58_LC_9_14_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i58_LC_9_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i58_LC_9_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8469),
            .lcout(\transmit_module.Y_DELTA_PATTERN_58 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24299),
            .ce(N__9895),
            .sr(N__23303));
    defparam \transmit_module.Y_DELTA_PATTERN_i57_LC_9_14_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i57_LC_9_14_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i57_LC_9_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i57_LC_9_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8475),
            .lcout(\transmit_module.Y_DELTA_PATTERN_57 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24299),
            .ce(N__9895),
            .sr(N__23303));
    defparam \transmit_module.Y_DELTA_PATTERN_i59_LC_9_14_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i59_LC_9_14_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i59_LC_9_14_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i59_LC_9_14_6  (
            .in0(N__8625),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.Y_DELTA_PATTERN_59 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24299),
            .ce(N__9895),
            .sr(N__23303));
    defparam \transmit_module.Y_DELTA_PATTERN_i56_LC_9_14_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i56_LC_9_14_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i56_LC_9_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i56_LC_9_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8463),
            .lcout(\transmit_module.Y_DELTA_PATTERN_56 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24299),
            .ce(N__9895),
            .sr(N__23303));
    defparam \transmit_module.Y_DELTA_PATTERN_i39_LC_9_15_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i39_LC_9_15_2 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i39_LC_9_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i39_LC_9_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8631),
            .lcout(\transmit_module.Y_DELTA_PATTERN_39 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24241),
            .ce(N__9913),
            .sr(N__23300));
    defparam \transmit_module.Y_DELTA_PATTERN_i44_LC_9_15_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i44_LC_9_15_7 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i44_LC_9_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i44_LC_9_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8442),
            .lcout(\transmit_module.Y_DELTA_PATTERN_44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24241),
            .ce(N__9913),
            .sr(N__23300));
    defparam \line_buffer.i2203_3_lut_LC_9_20_2 .C_ON=1'b0;
    defparam \line_buffer.i2203_3_lut_LC_9_20_2 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2203_3_lut_LC_9_20_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \line_buffer.i2203_3_lut_LC_9_20_2  (
            .in0(N__22827),
            .in1(N__8436),
            .in2(_gnd_net_),
            .in3(N__8424),
            .lcout(\line_buffer.n3540 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2191_3_lut_LC_9_20_4 .C_ON=1'b0;
    defparam \line_buffer.i2191_3_lut_LC_9_20_4 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2191_3_lut_LC_9_20_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \line_buffer.i2191_3_lut_LC_9_20_4  (
            .in0(N__22826),
            .in1(N__8541),
            .in2(_gnd_net_),
            .in3(N__8529),
            .lcout(\line_buffer.n3528 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.Y_DELTA_PATTERN_i28_LC_10_10_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i28_LC_10_10_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i28_LC_10_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i28_LC_10_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8685),
            .lcout(\transmit_module.Y_DELTA_PATTERN_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24334),
            .ce(N__20517),
            .sr(N__23333));
    defparam \transmit_module.Y_DELTA_PATTERN_i27_LC_10_11_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i27_LC_10_11_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i27_LC_10_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i27_LC_10_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8517),
            .lcout(\transmit_module.Y_DELTA_PATTERN_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24352),
            .ce(N__20499),
            .sr(N__23332));
    defparam \transmit_module.Y_DELTA_PATTERN_i8_LC_10_11_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i8_LC_10_11_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i8_LC_10_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i8_LC_10_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8691),
            .lcout(\transmit_module.Y_DELTA_PATTERN_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24352),
            .ce(N__20499),
            .sr(N__23332));
    defparam \transmit_module.Y_DELTA_PATTERN_i7_LC_10_11_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i7_LC_10_11_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i7_LC_10_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i7_LC_10_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8505),
            .lcout(\transmit_module.Y_DELTA_PATTERN_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24352),
            .ce(N__20499),
            .sr(N__23332));
    defparam \transmit_module.Y_DELTA_PATTERN_i48_LC_10_13_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i48_LC_10_13_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i48_LC_10_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i48_LC_10_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8583),
            .lcout(\transmit_module.Y_DELTA_PATTERN_48 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24350),
            .ce(N__9914),
            .sr(N__23284));
    defparam \transmit_module.Y_DELTA_PATTERN_i69_LC_10_13_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i69_LC_10_13_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i69_LC_10_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i69_LC_10_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8775),
            .lcout(\transmit_module.Y_DELTA_PATTERN_69 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24350),
            .ce(N__9914),
            .sr(N__23284));
    defparam \transmit_module.Y_DELTA_PATTERN_i47_LC_10_13_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i47_LC_10_13_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i47_LC_10_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i47_LC_10_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8499),
            .lcout(\transmit_module.Y_DELTA_PATTERN_47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24350),
            .ce(N__9914),
            .sr(N__23284));
    defparam \transmit_module.Y_DELTA_PATTERN_i50_LC_10_13_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i50_LC_10_13_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i50_LC_10_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i50_LC_10_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8781),
            .lcout(\transmit_module.Y_DELTA_PATTERN_50 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24350),
            .ce(N__9914),
            .sr(N__23284));
    defparam \transmit_module.Y_DELTA_PATTERN_i49_LC_10_13_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i49_LC_10_13_7 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i49_LC_10_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i49_LC_10_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8589),
            .lcout(\transmit_module.Y_DELTA_PATTERN_49 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24350),
            .ce(N__9914),
            .sr(N__23284));
    defparam \transmit_module.Y_DELTA_PATTERN_i53_LC_10_14_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i53_LC_10_14_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i53_LC_10_14_0 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i53_LC_10_14_0  (
            .in0(_gnd_net_),
            .in1(N__8577),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.Y_DELTA_PATTERN_53 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24287),
            .ce(N__9872),
            .sr(N__23310));
    defparam \transmit_module.Y_DELTA_PATTERN_i76_LC_10_14_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i76_LC_10_14_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i76_LC_10_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i76_LC_10_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8565),
            .lcout(\transmit_module.Y_DELTA_PATTERN_76 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24287),
            .ce(N__9872),
            .sr(N__23310));
    defparam \transmit_module.Y_DELTA_PATTERN_i67_LC_10_14_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i67_LC_10_14_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i67_LC_10_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i67_LC_10_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8553),
            .lcout(\transmit_module.Y_DELTA_PATTERN_67 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24287),
            .ce(N__9872),
            .sr(N__23310));
    defparam \transmit_module.Y_DELTA_PATTERN_i66_LC_10_14_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i66_LC_10_14_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i66_LC_10_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i66_LC_10_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8571),
            .lcout(\transmit_module.Y_DELTA_PATTERN_66 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24287),
            .ce(N__9872),
            .sr(N__23310));
    defparam \transmit_module.Y_DELTA_PATTERN_i77_LC_10_14_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i77_LC_10_14_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i77_LC_10_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i77_LC_10_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8892),
            .lcout(\transmit_module.Y_DELTA_PATTERN_77 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24287),
            .ce(N__9872),
            .sr(N__23310));
    defparam \transmit_module.Y_DELTA_PATTERN_i68_LC_10_14_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i68_LC_10_14_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i68_LC_10_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i68_LC_10_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8559),
            .lcout(\transmit_module.Y_DELTA_PATTERN_68 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24287),
            .ce(N__9872),
            .sr(N__23310));
    defparam \transmit_module.Y_DELTA_PATTERN_i75_LC_10_14_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i75_LC_10_14_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i75_LC_10_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i75_LC_10_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8547),
            .lcout(\transmit_module.Y_DELTA_PATTERN_75 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24287),
            .ce(N__9872),
            .sr(N__23310));
    defparam \transmit_module.Y_DELTA_PATTERN_i41_LC_10_15_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i41_LC_10_15_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i41_LC_10_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i41_LC_10_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8643),
            .lcout(\transmit_module.Y_DELTA_PATTERN_41 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24292),
            .ce(N__9908),
            .sr(N__23228));
    defparam \transmit_module.Y_DELTA_PATTERN_i65_LC_10_15_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i65_LC_10_15_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i65_LC_10_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i65_LC_10_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8661),
            .lcout(\transmit_module.Y_DELTA_PATTERN_65 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24292),
            .ce(N__9908),
            .sr(N__23228));
    defparam \transmit_module.Y_DELTA_PATTERN_i43_LC_10_15_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i43_LC_10_15_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i43_LC_10_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i43_LC_10_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8655),
            .lcout(\transmit_module.Y_DELTA_PATTERN_43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24292),
            .ce(N__9908),
            .sr(N__23228));
    defparam \transmit_module.Y_DELTA_PATTERN_i42_LC_10_15_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i42_LC_10_15_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i42_LC_10_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i42_LC_10_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8649),
            .lcout(\transmit_module.Y_DELTA_PATTERN_42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24292),
            .ce(N__9908),
            .sr(N__23228));
    defparam \transmit_module.Y_DELTA_PATTERN_i40_LC_10_15_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i40_LC_10_15_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i40_LC_10_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i40_LC_10_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8637),
            .lcout(\transmit_module.Y_DELTA_PATTERN_40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24292),
            .ce(N__9908),
            .sr(N__23228));
    defparam \transmit_module.Y_DELTA_PATTERN_i60_LC_10_15_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i60_LC_10_15_7 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i60_LC_10_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i60_LC_10_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8850),
            .lcout(\transmit_module.Y_DELTA_PATTERN_60 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24292),
            .ce(N__9908),
            .sr(N__23228));
    defparam \transmit_module.Y_DELTA_PATTERN_i6_LC_10_16_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i6_LC_10_16_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i6_LC_10_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i6_LC_10_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8619),
            .lcout(\transmit_module.Y_DELTA_PATTERN_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24291),
            .ce(N__20518),
            .sr(N__23327));
    defparam \transmit_module.Y_DELTA_PATTERN_i5_LC_10_18_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i5_LC_10_18_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i5_LC_10_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i5_LC_10_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8610),
            .lcout(\transmit_module.Y_DELTA_PATTERN_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24197),
            .ce(N__20525),
            .sr(N__23326));
    defparam \transmit_module.Y_DELTA_PATTERN_i4_LC_10_18_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i4_LC_10_18_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i4_LC_10_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i4_LC_10_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8601),
            .lcout(\transmit_module.Y_DELTA_PATTERN_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24197),
            .ce(N__20525),
            .sr(N__23326));
    defparam \transmit_module.Y_DELTA_PATTERN_i3_LC_10_18_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i3_LC_10_18_7 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i3_LC_10_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i3_LC_10_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8595),
            .lcout(\transmit_module.Y_DELTA_PATTERN_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24197),
            .ce(N__20525),
            .sr(N__23326));
    defparam \line_buffer.i2229_3_lut_LC_10_21_6 .C_ON=1'b0;
    defparam \line_buffer.i2229_3_lut_LC_10_21_6 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2229_3_lut_LC_10_21_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \line_buffer.i2229_3_lut_LC_10_21_6  (
            .in0(N__8769),
            .in1(N__8751),
            .in2(_gnd_net_),
            .in3(N__22831),
            .lcout(\line_buffer.n3566 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2232_3_lut_LC_11_9_4 .C_ON=1'b0;
    defparam \line_buffer.i2232_3_lut_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2232_3_lut_LC_11_9_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \line_buffer.i2232_3_lut_LC_11_9_4  (
            .in0(N__22828),
            .in1(N__8733),
            .in2(_gnd_net_),
            .in3(N__8718),
            .lcout(\line_buffer.n3569 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.BUFFER_0__i3_LC_11_9_5 .C_ON=1'b0;
    defparam \tvp_video_buffer.BUFFER_0__i3_LC_11_9_5 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.BUFFER_0__i3_LC_11_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.BUFFER_0__i3_LC_11_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8700),
            .lcout(\tvp_video_buffer.BUFFER_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21958),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.Y_DELTA_PATTERN_i32_LC_11_11_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i32_LC_11_11_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i32_LC_11_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i32_LC_11_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8832),
            .lcout(\transmit_module.Y_DELTA_PATTERN_32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24351),
            .ce(N__20488),
            .sr(N__23276));
    defparam \transmit_module.Y_DELTA_PATTERN_i9_LC_11_11_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i9_LC_11_11_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i9_LC_11_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i9_LC_11_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9036),
            .lcout(\transmit_module.Y_DELTA_PATTERN_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24351),
            .ce(N__20488),
            .sr(N__23276));
    defparam \transmit_module.Y_DELTA_PATTERN_i29_LC_11_11_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i29_LC_11_11_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i29_LC_11_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i29_LC_11_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8679),
            .lcout(\transmit_module.Y_DELTA_PATTERN_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24351),
            .ce(N__20488),
            .sr(N__23276));
    defparam \transmit_module.Y_DELTA_PATTERN_i30_LC_11_11_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i30_LC_11_11_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i30_LC_11_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i30_LC_11_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8667),
            .lcout(\transmit_module.Y_DELTA_PATTERN_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24351),
            .ce(N__20488),
            .sr(N__23276));
    defparam \transmit_module.Y_DELTA_PATTERN_i31_LC_11_11_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i31_LC_11_11_7 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i31_LC_11_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i31_LC_11_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8673),
            .lcout(\transmit_module.Y_DELTA_PATTERN_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24351),
            .ce(N__20488),
            .sr(N__23276));
    defparam \transmit_module.Y_DELTA_PATTERN_i35_LC_11_12_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i35_LC_11_12_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i35_LC_11_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i35_LC_11_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8817),
            .lcout(\transmit_module.Y_DELTA_PATTERN_35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24353),
            .ce(N__9915),
            .sr(N__23334));
    defparam \transmit_module.Y_DELTA_PATTERN_i33_LC_11_12_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i33_LC_11_12_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i33_LC_11_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i33_LC_11_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8805),
            .lcout(\transmit_module.Y_DELTA_PATTERN_33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24353),
            .ce(N__9915),
            .sr(N__23334));
    defparam \transmit_module.Y_DELTA_PATTERN_i36_LC_11_12_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i36_LC_11_12_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i36_LC_11_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i36_LC_11_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8826),
            .lcout(\transmit_module.Y_DELTA_PATTERN_36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24353),
            .ce(N__9915),
            .sr(N__23334));
    defparam \transmit_module.Y_DELTA_PATTERN_i34_LC_11_12_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i34_LC_11_12_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i34_LC_11_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i34_LC_11_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8811),
            .lcout(\transmit_module.Y_DELTA_PATTERN_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24353),
            .ce(N__9915),
            .sr(N__23334));
    defparam \transmit_module.Y_DELTA_PATTERN_i80_LC_11_13_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i80_LC_11_13_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i80_LC_11_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i80_LC_11_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8799),
            .lcout(\transmit_module.Y_DELTA_PATTERN_80 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24349),
            .ce(N__9899),
            .sr(N__23196));
    defparam \transmit_module.Y_DELTA_PATTERN_i81_LC_11_13_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i81_LC_11_13_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i81_LC_11_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i81_LC_11_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8793),
            .lcout(\transmit_module.Y_DELTA_PATTERN_81 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24349),
            .ce(N__9899),
            .sr(N__23196));
    defparam \transmit_module.Y_DELTA_PATTERN_i82_LC_11_13_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i82_LC_11_13_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i82_LC_11_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i82_LC_11_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21135),
            .lcout(\transmit_module.Y_DELTA_PATTERN_82 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24349),
            .ce(N__9899),
            .sr(N__23196));
    defparam \transmit_module.Y_DELTA_PATTERN_i79_LC_11_13_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i79_LC_11_13_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i79_LC_11_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i79_LC_11_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8787),
            .lcout(\transmit_module.Y_DELTA_PATTERN_79 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24349),
            .ce(N__9899),
            .sr(N__23196));
    defparam \transmit_module.Y_DELTA_PATTERN_i51_LC_11_13_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i51_LC_11_13_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i51_LC_11_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i51_LC_11_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8868),
            .lcout(\transmit_module.Y_DELTA_PATTERN_51 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24349),
            .ce(N__9899),
            .sr(N__23196));
    defparam \transmit_module.Y_DELTA_PATTERN_i70_LC_11_14_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i70_LC_11_14_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i70_LC_11_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i70_LC_11_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8904),
            .lcout(\transmit_module.Y_DELTA_PATTERN_70 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24271),
            .ce(N__9894),
            .sr(N__23323));
    defparam \transmit_module.Y_DELTA_PATTERN_i71_LC_11_14_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i71_LC_11_14_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i71_LC_11_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i71_LC_11_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8886),
            .lcout(\transmit_module.Y_DELTA_PATTERN_71 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24271),
            .ce(N__9894),
            .sr(N__23323));
    defparam \transmit_module.Y_DELTA_PATTERN_i78_LC_11_14_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i78_LC_11_14_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i78_LC_11_14_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i78_LC_11_14_3  (
            .in0(N__8898),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.Y_DELTA_PATTERN_78 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24271),
            .ce(N__9894),
            .sr(N__23323));
    defparam \transmit_module.Y_DELTA_PATTERN_i72_LC_11_14_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i72_LC_11_14_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i72_LC_11_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i72_LC_11_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8856),
            .lcout(\transmit_module.Y_DELTA_PATTERN_72 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24271),
            .ce(N__9894),
            .sr(N__23323));
    defparam \transmit_module.Y_DELTA_PATTERN_i74_LC_11_14_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i74_LC_11_14_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i74_LC_11_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i74_LC_11_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8880),
            .lcout(\transmit_module.Y_DELTA_PATTERN_74 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24271),
            .ce(N__9894),
            .sr(N__23323));
    defparam \transmit_module.Y_DELTA_PATTERN_i52_LC_11_14_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i52_LC_11_14_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i52_LC_11_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i52_LC_11_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8874),
            .lcout(\transmit_module.Y_DELTA_PATTERN_52 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24271),
            .ce(N__9894),
            .sr(N__23323));
    defparam \transmit_module.Y_DELTA_PATTERN_i73_LC_11_14_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i73_LC_11_14_7 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i73_LC_11_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i73_LC_11_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8862),
            .lcout(\transmit_module.Y_DELTA_PATTERN_73 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24271),
            .ce(N__9894),
            .sr(N__23323));
    defparam \transmit_module.Y_DELTA_PATTERN_i61_LC_11_15_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i61_LC_11_15_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i61_LC_11_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i61_LC_11_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8994),
            .lcout(\transmit_module.Y_DELTA_PATTERN_61 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24113),
            .ce(N__9904),
            .sr(N__23224));
    defparam \transmit_module.Y_DELTA_PATTERN_i63_LC_11_15_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i63_LC_11_15_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i63_LC_11_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i63_LC_11_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8838),
            .lcout(\transmit_module.Y_DELTA_PATTERN_63 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24113),
            .ce(N__9904),
            .sr(N__23224));
    defparam \transmit_module.Y_DELTA_PATTERN_i64_LC_11_15_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i64_LC_11_15_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i64_LC_11_15_4 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i64_LC_11_15_4  (
            .in0(_gnd_net_),
            .in1(N__8844),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.Y_DELTA_PATTERN_64 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24113),
            .ce(N__9904),
            .sr(N__23224));
    defparam \transmit_module.Y_DELTA_PATTERN_i62_LC_11_15_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i62_LC_11_15_7 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i62_LC_11_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i62_LC_11_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9000),
            .lcout(\transmit_module.Y_DELTA_PATTERN_62 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24113),
            .ce(N__9904),
            .sr(N__23224));
    defparam \transmit_module.ADDR_Y_COMPONENT__i11_LC_11_16_4 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i11_LC_11_16_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i11_LC_11_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i11_LC_11_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22767),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24222),
            .ce(N__15388),
            .sr(N__23324));
    defparam \transmit_module.ADDR_Y_COMPONENT__i10_LC_11_19_4 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i10_LC_11_19_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i10_LC_11_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i10_LC_11_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12369),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23973),
            .ce(N__15401),
            .sr(N__23296));
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_2266_LC_11_21_2 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_2266_LC_11_21_2 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_2266_LC_11_21_2 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \line_buffer.TX_ADDR_12__bdd_4_lut_2266_LC_11_21_2  (
            .in0(N__21507),
            .in1(N__8931),
            .in2(N__21306),
            .in3(N__8988),
            .lcout(),
            .ltout(\line_buffer.n3599_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i2_LC_11_21_3 .C_ON=1'b0;
    defparam \line_buffer.dout_i2_LC_11_21_3 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i2_LC_11_21_3 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \line_buffer.dout_i2_LC_11_21_3  (
            .in0(N__21304),
            .in1(N__8976),
            .in2(N__8970),
            .in3(N__9084),
            .lcout(TX_DATA_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23972),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2233_3_lut_LC_11_22_4 .C_ON=1'b0;
    defparam \line_buffer.i2233_3_lut_LC_11_22_4 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2233_3_lut_LC_11_22_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \line_buffer.i2233_3_lut_LC_11_22_4  (
            .in0(N__8967),
            .in1(N__22829),
            .in2(_gnd_net_),
            .in3(N__8955),
            .lcout(\line_buffer.n3570 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.BUFFER_0__i2_LC_12_4_1 .C_ON=1'b0;
    defparam \tvp_video_buffer.BUFFER_0__i2_LC_12_4_1 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.BUFFER_0__i2_LC_12_4_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.BUFFER_0__i2_LC_12_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8925),
            .lcout(\tvp_video_buffer.BUFFER_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21931),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.BUFFER_0__i10_LC_12_4_2 .C_ON=1'b0;
    defparam \tvp_video_buffer.BUFFER_0__i10_LC_12_4_2 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.BUFFER_0__i10_LC_12_4_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.BUFFER_0__i10_LC_12_4_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8910),
            .lcout(\tvp_video_buffer.BUFFER_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21931),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.Y_DELTA_PATTERN_i12_LC_12_10_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i12_LC_12_10_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i12_LC_12_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i12_LC_12_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9567),
            .lcout(\transmit_module.Y_DELTA_PATTERN_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24332),
            .ce(N__20510),
            .sr(N__23275));
    defparam \transmit_module.Y_DELTA_PATTERN_i11_LC_12_10_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i11_LC_12_10_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i11_LC_12_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i11_LC_12_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9048),
            .lcout(\transmit_module.Y_DELTA_PATTERN_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24332),
            .ce(N__20510),
            .sr(N__23275));
    defparam \transmit_module.Y_DELTA_PATTERN_i10_LC_12_10_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i10_LC_12_10_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i10_LC_12_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i10_LC_12_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9042),
            .lcout(\transmit_module.Y_DELTA_PATTERN_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24332),
            .ce(N__20510),
            .sr(N__23275));
    defparam \sync_buffer.BUFFER_0__i1_LC_12_13_1 .C_ON=1'b0;
    defparam \sync_buffer.BUFFER_0__i1_LC_12_13_1 .SEQ_MODE=4'b1000;
    defparam \sync_buffer.BUFFER_0__i1_LC_12_13_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \sync_buffer.BUFFER_0__i1_LC_12_13_1  (
            .in0(N__15540),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\sync_buffer.BUFFER_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24229),
            .ce(),
            .sr(_gnd_net_));
    defparam \sync_buffer.WIRE_OUT_0__9_LC_12_13_3 .C_ON=1'b0;
    defparam \sync_buffer.WIRE_OUT_0__9_LC_12_13_3 .SEQ_MODE=4'b1000;
    defparam \sync_buffer.WIRE_OUT_0__9_LC_12_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sync_buffer.WIRE_OUT_0__9_LC_12_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9024),
            .lcout(RX_TX_SYNC_BUFF),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24229),
            .ce(),
            .sr(_gnd_net_));
    defparam \sync_buffer.BUFFER_0__i2_LC_12_13_5 .C_ON=1'b0;
    defparam \sync_buffer.BUFFER_0__i2_LC_12_13_5 .SEQ_MODE=4'b1000;
    defparam \sync_buffer.BUFFER_0__i2_LC_12_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \sync_buffer.BUFFER_0__i2_LC_12_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9030),
            .lcout(\sync_buffer.BUFFER_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24229),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1160_2_lut_LC_12_13_6 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1160_2_lut_LC_12_13_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1160_2_lut_LC_12_13_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \transmit_module.video_signal_controller.i1160_2_lut_LC_12_13_6  (
            .in0(_gnd_net_),
            .in1(N__9018),
            .in2(_gnd_net_),
            .in3(N__11891),
            .lcout(\transmit_module.video_signal_controller.n2395 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i2_4_lut_adj_30_LC_12_14_4 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i2_4_lut_adj_30_LC_12_14_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i2_4_lut_adj_30_LC_12_14_4 .LUT_INIT=16'b1010000010000000;
    LogicCell40 \transmit_module.video_signal_controller.i2_4_lut_adj_30_LC_12_14_4  (
            .in0(N__9687),
            .in1(N__9939),
            .in2(N__9786),
            .in3(N__9660),
            .lcout(),
            .ltout(\transmit_module.video_signal_controller.n3479_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i3_4_lut_LC_12_14_5 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i3_4_lut_LC_12_14_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i3_4_lut_LC_12_14_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \transmit_module.video_signal_controller.i3_4_lut_LC_12_14_5  (
            .in0(N__9735),
            .in1(N__9759),
            .in2(N__9012),
            .in3(N__9815),
            .lcout(),
            .ltout(\transmit_module.video_signal_controller.n3475_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i2_4_lut_adj_32_LC_12_14_6 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i2_4_lut_adj_32_LC_12_14_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i2_4_lut_adj_32_LC_12_14_6 .LUT_INIT=16'b0000010101000100;
    LogicCell40 \transmit_module.video_signal_controller.i2_4_lut_adj_32_LC_12_14_6  (
            .in0(N__12193),
            .in1(N__9006),
            .in2(N__9009),
            .in3(N__9711),
            .lcout(\transmit_module.video_signal_controller.n7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_4_lut_adj_31_LC_12_14_7 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_4_lut_adj_31_LC_12_14_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_4_lut_adj_31_LC_12_14_7 .LUT_INIT=16'b1110111011101010;
    LogicCell40 \transmit_module.video_signal_controller.i1_4_lut_adj_31_LC_12_14_7  (
            .in0(N__9734),
            .in1(N__9758),
            .in2(N__9816),
            .in3(N__9785),
            .lcout(\transmit_module.video_signal_controller.n55 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2230_3_lut_LC_12_15_3 .C_ON=1'b0;
    defparam \line_buffer.i2230_3_lut_LC_12_15_3 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2230_3_lut_LC_12_15_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \line_buffer.i2230_3_lut_LC_12_15_3  (
            .in0(N__9114),
            .in1(N__9102),
            .in2(_gnd_net_),
            .in3(N__22821),
            .lcout(\line_buffer.n3567 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.VGA_X_i0_LC_12_16_0 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i0_LC_12_16_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i0_LC_12_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i0_LC_12_16_0  (
            .in0(_gnd_net_),
            .in1(N__9937),
            .in2(_gnd_net_),
            .in3(N__9072),
            .lcout(\transmit_module.video_signal_controller.VGA_X_0 ),
            .ltout(),
            .carryin(bfn_12_16_0_),
            .carryout(\transmit_module.video_signal_controller.n3180 ),
            .clk(N__24221),
            .ce(),
            .sr(N__11900));
    defparam \transmit_module.video_signal_controller.VGA_X_i1_LC_12_16_1 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i1_LC_12_16_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i1_LC_12_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i1_LC_12_16_1  (
            .in0(_gnd_net_),
            .in1(N__9655),
            .in2(_gnd_net_),
            .in3(N__9069),
            .lcout(\transmit_module.video_signal_controller.VGA_X_1 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3180 ),
            .carryout(\transmit_module.video_signal_controller.n3181 ),
            .clk(N__24221),
            .ce(),
            .sr(N__11900));
    defparam \transmit_module.video_signal_controller.VGA_X_i2_LC_12_16_2 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i2_LC_12_16_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i2_LC_12_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i2_LC_12_16_2  (
            .in0(_gnd_net_),
            .in1(N__9685),
            .in2(_gnd_net_),
            .in3(N__9066),
            .lcout(\transmit_module.video_signal_controller.VGA_X_2 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3181 ),
            .carryout(\transmit_module.video_signal_controller.n3182 ),
            .clk(N__24221),
            .ce(),
            .sr(N__11900));
    defparam \transmit_module.video_signal_controller.VGA_X_i3_LC_12_16_3 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i3_LC_12_16_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i3_LC_12_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i3_LC_12_16_3  (
            .in0(_gnd_net_),
            .in1(N__9780),
            .in2(_gnd_net_),
            .in3(N__9063),
            .lcout(\transmit_module.video_signal_controller.VGA_X_3 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3182 ),
            .carryout(\transmit_module.video_signal_controller.n3183 ),
            .clk(N__24221),
            .ce(),
            .sr(N__11900));
    defparam \transmit_module.video_signal_controller.VGA_X_i4_LC_12_16_4 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i4_LC_12_16_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i4_LC_12_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i4_LC_12_16_4  (
            .in0(_gnd_net_),
            .in1(N__9810),
            .in2(_gnd_net_),
            .in3(N__9060),
            .lcout(\transmit_module.video_signal_controller.VGA_X_4 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3183 ),
            .carryout(\transmit_module.video_signal_controller.n3184 ),
            .clk(N__24221),
            .ce(),
            .sr(N__11900));
    defparam \transmit_module.video_signal_controller.VGA_X_i5_LC_12_16_5 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i5_LC_12_16_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i5_LC_12_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i5_LC_12_16_5  (
            .in0(_gnd_net_),
            .in1(N__9756),
            .in2(_gnd_net_),
            .in3(N__9057),
            .lcout(\transmit_module.video_signal_controller.VGA_X_5 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3184 ),
            .carryout(\transmit_module.video_signal_controller.n3185 ),
            .clk(N__24221),
            .ce(),
            .sr(N__11900));
    defparam \transmit_module.video_signal_controller.VGA_X_i6_LC_12_16_6 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i6_LC_12_16_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i6_LC_12_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i6_LC_12_16_6  (
            .in0(_gnd_net_),
            .in1(N__9732),
            .in2(_gnd_net_),
            .in3(N__9054),
            .lcout(\transmit_module.video_signal_controller.VGA_X_6 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3185 ),
            .carryout(\transmit_module.video_signal_controller.n3186 ),
            .clk(N__24221),
            .ce(),
            .sr(N__11900));
    defparam \transmit_module.video_signal_controller.VGA_X_i7_LC_12_16_7 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i7_LC_12_16_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i7_LC_12_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i7_LC_12_16_7  (
            .in0(_gnd_net_),
            .in1(N__9709),
            .in2(_gnd_net_),
            .in3(N__9051),
            .lcout(\transmit_module.video_signal_controller.VGA_X_7 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3186 ),
            .carryout(\transmit_module.video_signal_controller.n3187 ),
            .clk(N__24221),
            .ce(),
            .sr(N__11900));
    defparam \transmit_module.video_signal_controller.VGA_X_i8_LC_12_17_0 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i8_LC_12_17_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i8_LC_12_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i8_LC_12_17_0  (
            .in0(_gnd_net_),
            .in1(N__11949),
            .in2(_gnd_net_),
            .in3(N__9189),
            .lcout(\transmit_module.video_signal_controller.VGA_X_8 ),
            .ltout(),
            .carryin(bfn_12_17_0_),
            .carryout(\transmit_module.video_signal_controller.n3188 ),
            .clk(N__24067),
            .ce(),
            .sr(N__11904));
    defparam \transmit_module.video_signal_controller.VGA_X_i9_LC_12_17_1 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i9_LC_12_17_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i9_LC_12_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i9_LC_12_17_1  (
            .in0(_gnd_net_),
            .in1(N__12150),
            .in2(_gnd_net_),
            .in3(N__9186),
            .lcout(\transmit_module.video_signal_controller.VGA_X_9 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3188 ),
            .carryout(\transmit_module.video_signal_controller.n3189 ),
            .clk(N__24067),
            .ce(),
            .sr(N__11904));
    defparam \transmit_module.video_signal_controller.VGA_X_i10_LC_12_17_2 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i10_LC_12_17_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i10_LC_12_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i10_LC_12_17_2  (
            .in0(_gnd_net_),
            .in1(N__12189),
            .in2(_gnd_net_),
            .in3(N__9183),
            .lcout(\transmit_module.video_signal_controller.VGA_X_10 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3189 ),
            .carryout(\transmit_module.video_signal_controller.n3190 ),
            .clk(N__24067),
            .ce(),
            .sr(N__11904));
    defparam \transmit_module.video_signal_controller.VGA_X_i11_LC_12_17_3 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.VGA_X_i11_LC_12_17_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i11_LC_12_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i11_LC_12_17_3  (
            .in0(_gnd_net_),
            .in1(N__12242),
            .in2(_gnd_net_),
            .in3(N__9180),
            .lcout(\transmit_module.video_signal_controller.VGA_X_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24067),
            .ce(),
            .sr(N__11904));
    defparam \transmit_module.Y_DELTA_PATTERN_i0_LC_12_18_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i0_LC_12_18_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i0_LC_12_18_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i0_LC_12_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9162),
            .lcout(\transmit_module.Y_DELTA_PATTERN_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23978),
            .ce(N__20526),
            .sr(N__23336));
    defparam \transmit_module.Y_DELTA_PATTERN_i2_LC_12_18_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i2_LC_12_18_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i2_LC_12_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i2_LC_12_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9177),
            .lcout(\transmit_module.Y_DELTA_PATTERN_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23978),
            .ce(N__20526),
            .sr(N__23336));
    defparam \transmit_module.Y_DELTA_PATTERN_i1_LC_12_18_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i1_LC_12_18_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i1_LC_12_18_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i1_LC_12_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9168),
            .lcout(\transmit_module.Y_DELTA_PATTERN_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23978),
            .ce(N__20526),
            .sr(N__23336));
    defparam \line_buffer.i2190_3_lut_LC_12_19_6 .C_ON=1'b0;
    defparam \line_buffer.i2190_3_lut_LC_12_19_6 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2190_3_lut_LC_12_19_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \line_buffer.i2190_3_lut_LC_12_19_6  (
            .in0(N__22808),
            .in1(N__9156),
            .in2(_gnd_net_),
            .in3(N__9144),
            .lcout(\line_buffer.n3527 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_LC_12_20_4 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_LC_12_20_4 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_LC_12_20_4 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \line_buffer.TX_ADDR_12__bdd_4_lut_LC_12_20_4  (
            .in0(N__21498),
            .in1(N__9123),
            .in2(N__21300),
            .in3(N__9432),
            .lcout(\line_buffer.n3617 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.VGA_R__i3_LC_12_22_6 .C_ON=1'b0;
    defparam \transmit_module.VGA_R__i3_LC_12_22_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.VGA_R__i3_LC_12_22_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.VGA_R__i3_LC_12_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9426),
            .lcout(n1816),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23951),
            .ce(),
            .sr(N__22424));
    defparam \line_buffer.i2193_3_lut_LC_12_25_0 .C_ON=1'b0;
    defparam \line_buffer.i2193_3_lut_LC_12_25_0 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2193_3_lut_LC_12_25_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \line_buffer.i2193_3_lut_LC_12_25_0  (
            .in0(N__9369),
            .in1(N__22830),
            .in2(_gnd_net_),
            .in3(N__9357),
            .lcout(\line_buffer.n3530 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.WIRE_OUT_i1_LC_13_4_6 .C_ON=1'b0;
    defparam \tvp_video_buffer.WIRE_OUT_i1_LC_13_4_6 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.WIRE_OUT_i1_LC_13_4_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.WIRE_OUT_i1_LC_13_4_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9345),
            .lcout(RX_DATA_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21929),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.WIRE_OUT_i5_LC_13_5_0 .C_ON=1'b0;
    defparam \tvp_video_buffer.WIRE_OUT_i5_LC_13_5_0 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.WIRE_OUT_i5_LC_13_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.WIRE_OUT_i5_LC_13_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9246),
            .lcout(RX_DATA_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21932),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.BUFFER_0__i14_LC_13_5_2 .C_ON=1'b0;
    defparam \tvp_video_buffer.BUFFER_0__i14_LC_13_5_2 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.BUFFER_0__i14_LC_13_5_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.BUFFER_0__i14_LC_13_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9204),
            .lcout(\tvp_video_buffer.BUFFER_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21932),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.BUFFER_0__i6_LC_13_5_6 .C_ON=1'b0;
    defparam \tvp_video_buffer.BUFFER_0__i6_LC_13_5_6 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.BUFFER_0__i6_LC_13_5_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \tvp_video_buffer.BUFFER_0__i6_LC_13_5_6  (
            .in0(N__9230),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\tvp_video_buffer.BUFFER_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21932),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.BUFFER_0__i11_LC_13_9_0 .C_ON=1'b0;
    defparam \tvp_video_buffer.BUFFER_0__i11_LC_13_9_0 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.BUFFER_0__i11_LC_13_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.BUFFER_0__i11_LC_13_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9198),
            .lcout(\tvp_video_buffer.BUFFER_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21951),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.Y_DELTA_PATTERN_i16_LC_13_10_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i16_LC_13_10_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i16_LC_13_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i16_LC_13_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9579),
            .lcout(\transmit_module.Y_DELTA_PATTERN_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24300),
            .ce(N__20503),
            .sr(N__23198));
    defparam \transmit_module.Y_DELTA_PATTERN_i17_LC_13_10_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i17_LC_13_10_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i17_LC_13_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i17_LC_13_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9549),
            .lcout(\transmit_module.Y_DELTA_PATTERN_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24300),
            .ce(N__20503),
            .sr(N__23198));
    defparam \transmit_module.Y_DELTA_PATTERN_i15_LC_13_10_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i15_LC_13_10_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i15_LC_13_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i15_LC_13_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9573),
            .lcout(\transmit_module.Y_DELTA_PATTERN_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24300),
            .ce(N__20503),
            .sr(N__23198));
    defparam \transmit_module.Y_DELTA_PATTERN_i13_LC_13_10_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i13_LC_13_10_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i13_LC_13_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i13_LC_13_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9555),
            .lcout(\transmit_module.Y_DELTA_PATTERN_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24300),
            .ce(N__20503),
            .sr(N__23198));
    defparam \transmit_module.Y_DELTA_PATTERN_i14_LC_13_10_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i14_LC_13_10_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i14_LC_13_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i14_LC_13_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9561),
            .lcout(\transmit_module.Y_DELTA_PATTERN_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24300),
            .ce(N__20503),
            .sr(N__23198));
    defparam \transmit_module.Y_DELTA_PATTERN_i18_LC_13_10_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i18_LC_13_10_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i18_LC_13_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i18_LC_13_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11451),
            .lcout(\transmit_module.Y_DELTA_PATTERN_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24300),
            .ce(N__20503),
            .sr(N__23198));
    defparam \tvp_video_buffer.WIRE_OUT_i2_LC_13_11_0 .C_ON=1'b0;
    defparam \tvp_video_buffer.WIRE_OUT_i2_LC_13_11_0 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.WIRE_OUT_i2_LC_13_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.WIRE_OUT_i2_LC_13_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9543),
            .lcout(RX_DATA_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21959),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.VGA_Y_i0_LC_13_12_0 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i0_LC_13_12_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i0_LC_13_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i0_LC_13_12_0  (
            .in0(_gnd_net_),
            .in1(N__11972),
            .in2(_gnd_net_),
            .in3(N__9441),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_0 ),
            .ltout(),
            .carryin(bfn_13_12_0_),
            .carryout(\transmit_module.video_signal_controller.n3191 ),
            .clk(N__24283),
            .ce(N__11899),
            .sr(N__9597));
    defparam \transmit_module.video_signal_controller.VGA_Y_i1_LC_13_12_1 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i1_LC_13_12_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i1_LC_13_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i1_LC_13_12_1  (
            .in0(_gnd_net_),
            .in1(N__11993),
            .in2(_gnd_net_),
            .in3(N__9438),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_1 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3191 ),
            .carryout(\transmit_module.video_signal_controller.n3192 ),
            .clk(N__24283),
            .ce(N__11899),
            .sr(N__9597));
    defparam \transmit_module.video_signal_controller.VGA_Y_i2_LC_13_12_2 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i2_LC_13_12_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i2_LC_13_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i2_LC_13_12_2  (
            .in0(_gnd_net_),
            .in1(N__12026),
            .in2(_gnd_net_),
            .in3(N__9435),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_2 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3192 ),
            .carryout(\transmit_module.video_signal_controller.n3193 ),
            .clk(N__24283),
            .ce(N__11899),
            .sr(N__9597));
    defparam \transmit_module.video_signal_controller.VGA_Y_i3_LC_13_12_3 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i3_LC_13_12_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i3_LC_13_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i3_LC_13_12_3  (
            .in0(_gnd_net_),
            .in1(N__11760),
            .in2(_gnd_net_),
            .in3(N__9624),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_3 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3193 ),
            .carryout(\transmit_module.video_signal_controller.n3194 ),
            .clk(N__24283),
            .ce(N__11899),
            .sr(N__9597));
    defparam \transmit_module.video_signal_controller.VGA_Y_i4_LC_13_12_4 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i4_LC_13_12_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i4_LC_13_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i4_LC_13_12_4  (
            .in0(_gnd_net_),
            .in1(N__11742),
            .in2(_gnd_net_),
            .in3(N__9621),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_4 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3194 ),
            .carryout(\transmit_module.video_signal_controller.n3195 ),
            .clk(N__24283),
            .ce(N__11899),
            .sr(N__9597));
    defparam \transmit_module.video_signal_controller.VGA_Y_i5_LC_13_12_5 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i5_LC_13_12_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i5_LC_13_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i5_LC_13_12_5  (
            .in0(_gnd_net_),
            .in1(N__11703),
            .in2(_gnd_net_),
            .in3(N__9618),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_5 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3195 ),
            .carryout(\transmit_module.video_signal_controller.n3196 ),
            .clk(N__24283),
            .ce(N__11899),
            .sr(N__9597));
    defparam \transmit_module.video_signal_controller.VGA_Y_i6_LC_13_12_6 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i6_LC_13_12_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i6_LC_13_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i6_LC_13_12_6  (
            .in0(_gnd_net_),
            .in1(N__11718),
            .in2(_gnd_net_),
            .in3(N__9615),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_6 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3196 ),
            .carryout(\transmit_module.video_signal_controller.n3197 ),
            .clk(N__24283),
            .ce(N__11899),
            .sr(N__9597));
    defparam \transmit_module.video_signal_controller.VGA_Y_i7_LC_13_12_7 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i7_LC_13_12_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i7_LC_13_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i7_LC_13_12_7  (
            .in0(_gnd_net_),
            .in1(N__11664),
            .in2(_gnd_net_),
            .in3(N__9612),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_7 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3197 ),
            .carryout(\transmit_module.video_signal_controller.n3198 ),
            .clk(N__24283),
            .ce(N__11899),
            .sr(N__9597));
    defparam \transmit_module.video_signal_controller.VGA_Y_i8_LC_13_13_0 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i8_LC_13_13_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i8_LC_13_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i8_LC_13_13_0  (
            .in0(_gnd_net_),
            .in1(N__11676),
            .in2(_gnd_net_),
            .in3(N__9609),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_8 ),
            .ltout(),
            .carryin(bfn_13_13_0_),
            .carryout(\transmit_module.video_signal_controller.n3199 ),
            .clk(N__24228),
            .ce(N__11898),
            .sr(N__9593));
    defparam \transmit_module.video_signal_controller.VGA_Y_i9_LC_13_13_1 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i9_LC_13_13_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i9_LC_13_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i9_LC_13_13_1  (
            .in0(_gnd_net_),
            .in1(N__13694),
            .in2(_gnd_net_),
            .in3(N__9606),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_9 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3199 ),
            .carryout(\transmit_module.video_signal_controller.n3200 ),
            .clk(N__24228),
            .ce(N__11898),
            .sr(N__9593));
    defparam \transmit_module.video_signal_controller.VGA_Y_i10_LC_13_13_2 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i10_LC_13_13_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i10_LC_13_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i10_LC_13_13_2  (
            .in0(_gnd_net_),
            .in1(N__13737),
            .in2(_gnd_net_),
            .in3(N__9603),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_10 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3200 ),
            .carryout(\transmit_module.video_signal_controller.n3201 ),
            .clk(N__24228),
            .ce(N__11898),
            .sr(N__9593));
    defparam \transmit_module.video_signal_controller.VGA_Y_i11_LC_13_13_3 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.VGA_Y_i11_LC_13_13_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i11_LC_13_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i11_LC_13_13_3  (
            .in0(_gnd_net_),
            .in1(N__13757),
            .in2(_gnd_net_),
            .in3(N__9600),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24228),
            .ce(N__11898),
            .sr(N__9593));
    defparam \transmit_module.video_signal_controller.VGA_HS_66_LC_13_14_0 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.VGA_HS_66_LC_13_14_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_HS_66_LC_13_14_0 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \transmit_module.video_signal_controller.VGA_HS_66_LC_13_14_0  (
            .in0(N__12159),
            .in1(N__11954),
            .in2(N__12256),
            .in3(N__9945),
            .lcout(ADV_HSYNC_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24270),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1712_2_lut_3_lut_LC_13_14_2 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1712_2_lut_3_lut_LC_13_14_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1712_2_lut_3_lut_LC_13_14_2 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \transmit_module.video_signal_controller.i1712_2_lut_3_lut_LC_13_14_2  (
            .in0(N__9686),
            .in1(N__9659),
            .in2(_gnd_net_),
            .in3(N__9938),
            .lcout(\transmit_module.video_signal_controller.n2955 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.old_VGA_HS_40_LC_13_14_3 .C_ON=1'b0;
    defparam \transmit_module.old_VGA_HS_40_LC_13_14_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.old_VGA_HS_40_LC_13_14_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \transmit_module.old_VGA_HS_40_LC_13_14_3  (
            .in0(N__11816),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.old_VGA_HS ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24270),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i124_2_lut_4_lut_rep_24_LC_13_14_4 .C_ON=1'b0;
    defparam \transmit_module.i124_2_lut_4_lut_rep_24_LC_13_14_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i124_2_lut_4_lut_rep_24_LC_13_14_4 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \transmit_module.i124_2_lut_4_lut_rep_24_LC_13_14_4  (
            .in0(N__11857),
            .in1(N__11787),
            .in2(N__23174),
            .in3(N__11815),
            .lcout(\transmit_module.n3680 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_2_lut_adj_33_LC_13_14_5 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_2_lut_adj_33_LC_13_14_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_2_lut_adj_33_LC_13_14_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \transmit_module.video_signal_controller.i1_2_lut_adj_33_LC_13_14_5  (
            .in0(_gnd_net_),
            .in1(N__9811),
            .in2(_gnd_net_),
            .in3(N__9781),
            .lcout(\transmit_module.video_signal_controller.n3363 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i2_3_lut_adj_34_LC_13_14_6 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i2_3_lut_adj_34_LC_13_14_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i2_3_lut_adj_34_LC_13_14_6 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \transmit_module.video_signal_controller.i2_3_lut_adj_34_LC_13_14_6  (
            .in0(N__9757),
            .in1(N__9733),
            .in2(_gnd_net_),
            .in3(N__9710),
            .lcout(\transmit_module.video_signal_controller.n2014 ),
            .ltout(\transmit_module.video_signal_controller.n2014_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1761_4_lut_LC_13_14_7 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1761_4_lut_LC_13_14_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1761_4_lut_LC_13_14_7 .LUT_INIT=16'b1010100010100000;
    LogicCell40 \transmit_module.video_signal_controller.i1761_4_lut_LC_13_14_7  (
            .in0(N__11953),
            .in1(N__9630),
            .in2(N__9690),
            .in3(N__11927),
            .lcout(\transmit_module.video_signal_controller.n3004 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1_3_lut_LC_13_15_0 .C_ON=1'b0;
    defparam \transmit_module.i1_3_lut_LC_13_15_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1_3_lut_LC_13_15_0 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \transmit_module.i1_3_lut_LC_13_15_0  (
            .in0(N__16240),
            .in1(N__23120),
            .in2(_gnd_net_),
            .in3(N__20633),
            .lcout(\transmit_module.n2310 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i506_2_lut_rep_20_LC_13_15_1 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i506_2_lut_rep_20_LC_13_15_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i506_2_lut_rep_20_LC_13_15_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \transmit_module.video_signal_controller.i506_2_lut_rep_20_LC_13_15_1  (
            .in0(_gnd_net_),
            .in1(N__9684),
            .in2(_gnd_net_),
            .in3(N__9654),
            .lcout(\transmit_module.video_signal_controller.n3676 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i7_LC_13_15_2 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i7_LC_13_15_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i7_LC_13_15_2 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \transmit_module.BRAM_ADDR__i7_LC_13_15_2  (
            .in0(N__16241),
            .in1(N__23121),
            .in2(N__13005),
            .in3(N__13020),
            .lcout(\transmit_module.TX_ADDR_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24115),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i1_LC_13_15_5 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i1_LC_13_15_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i1_LC_13_15_5 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \transmit_module.BRAM_ADDR__i1_LC_13_15_5  (
            .in0(N__16265),
            .in1(N__10683),
            .in2(N__23240),
            .in3(N__10182),
            .lcout(\transmit_module.TX_ADDR_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24115),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_14_i2_3_lut_LC_13_15_6 .C_ON=1'b0;
    defparam \transmit_module.mux_14_i2_3_lut_LC_13_15_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_14_i2_3_lut_LC_13_15_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \transmit_module.mux_14_i2_3_lut_LC_13_15_6  (
            .in0(N__12460),
            .in1(N__14024),
            .in2(_gnd_net_),
            .in3(N__12117),
            .lcout(\transmit_module.n146 ),
            .ltout(\transmit_module.n146_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1643_4_lut_LC_13_15_7 .C_ON=1'b0;
    defparam \transmit_module.i1643_4_lut_LC_13_15_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1643_4_lut_LC_13_15_7 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \transmit_module.i1643_4_lut_LC_13_15_7  (
            .in0(N__23119),
            .in1(N__16239),
            .in2(N__10176),
            .in3(N__10682),
            .lcout(n27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i10_3_lut_LC_13_16_0 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i10_3_lut_LC_13_16_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i10_3_lut_LC_13_16_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_12_i10_3_lut_LC_13_16_0  (
            .in0(N__20626),
            .in1(N__12477),
            .in2(_gnd_net_),
            .in3(N__12500),
            .lcout(\transmit_module.n107 ),
            .ltout(\transmit_module.n107_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i9_LC_13_16_1 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i9_LC_13_16_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i9_LC_13_16_1 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \transmit_module.BRAM_ADDR__i9_LC_13_16_1  (
            .in0(N__10428),
            .in1(N__23125),
            .in2(N__9951),
            .in3(N__16317),
            .lcout(\transmit_module.TX_ADDR_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24184),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_14_i3_3_lut_LC_13_16_2 .C_ON=1'b0;
    defparam \transmit_module.mux_14_i3_3_lut_LC_13_16_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_14_i3_3_lut_LC_13_16_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \transmit_module.mux_14_i3_3_lut_LC_13_16_2  (
            .in0(N__12106),
            .in1(N__14027),
            .in2(_gnd_net_),
            .in3(N__12084),
            .lcout(\transmit_module.n145 ),
            .ltout(\transmit_module.n145_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i2_LC_13_16_3 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i2_LC_13_16_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i2_LC_13_16_3 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \transmit_module.BRAM_ADDR__i2_LC_13_16_3  (
            .in0(N__23253),
            .in1(N__16314),
            .in2(N__9948),
            .in3(N__10956),
            .lcout(\transmit_module.TX_ADDR_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24184),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i3_LC_13_16_4 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i3_LC_13_16_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i3_LC_13_16_4 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \transmit_module.BRAM_ADDR__i3_LC_13_16_4  (
            .in0(N__16315),
            .in1(N__10704),
            .in2(N__23241),
            .in3(N__10941),
            .lcout(\transmit_module.TX_ADDR_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24184),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i5_LC_13_16_6 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i5_LC_13_16_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i5_LC_13_16_6 .LUT_INIT=16'b0000111000000100;
    LogicCell40 \transmit_module.BRAM_ADDR__i5_LC_13_16_6  (
            .in0(N__16316),
            .in1(N__10674),
            .in2(N__23242),
            .in3(N__10440),
            .lcout(\transmit_module.TX_ADDR_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24184),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i2_3_lut_LC_13_16_7 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i2_3_lut_LC_13_16_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i2_3_lut_LC_13_16_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \transmit_module.mux_12_i2_3_lut_LC_13_16_7  (
            .in0(N__12461),
            .in1(N__12435),
            .in2(_gnd_net_),
            .in3(N__20627),
            .lcout(\transmit_module.n115 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_14_i6_3_lut_LC_13_17_1 .C_ON=1'b0;
    defparam \transmit_module.mux_14_i6_3_lut_LC_13_17_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_14_i6_3_lut_LC_13_17_1 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \transmit_module.mux_14_i6_3_lut_LC_13_17_1  (
            .in0(_gnd_net_),
            .in1(N__14029),
            .in2(N__12327),
            .in3(N__12396),
            .lcout(\transmit_module.n142 ),
            .ltout(\transmit_module.n142_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1647_4_lut_LC_13_17_2 .C_ON=1'b0;
    defparam \transmit_module.i1647_4_lut_LC_13_17_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1647_4_lut_LC_13_17_2 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \transmit_module.i1647_4_lut_LC_13_17_2  (
            .in0(N__23212),
            .in1(N__16304),
            .in2(N__10668),
            .in3(N__10439),
            .lcout(n23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i8_LC_13_17_3 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i8_LC_13_17_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i8_LC_13_17_3 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \transmit_module.BRAM_ADDR__i8_LC_13_17_3  (
            .in0(N__16307),
            .in1(N__11439),
            .in2(N__23299),
            .in3(N__11445),
            .lcout(\transmit_module.TX_ADDR_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24208),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i6_3_lut_LC_13_17_4 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i6_3_lut_LC_13_17_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i6_3_lut_LC_13_17_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \transmit_module.mux_12_i6_3_lut_LC_13_17_4  (
            .in0(N__12397),
            .in1(N__20592),
            .in2(_gnd_net_),
            .in3(N__12375),
            .lcout(\transmit_module.n111 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_14_i10_3_lut_LC_13_17_5 .C_ON=1'b0;
    defparam \transmit_module.mux_14_i10_3_lut_LC_13_17_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_14_i10_3_lut_LC_13_17_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \transmit_module.mux_14_i10_3_lut_LC_13_17_5  (
            .in0(N__12499),
            .in1(N__14028),
            .in2(_gnd_net_),
            .in3(N__12294),
            .lcout(\transmit_module.n138 ),
            .ltout(\transmit_module.n138_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1651_4_lut_LC_13_17_6 .C_ON=1'b0;
    defparam \transmit_module.i1651_4_lut_LC_13_17_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1651_4_lut_LC_13_17_6 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \transmit_module.i1651_4_lut_LC_13_17_6  (
            .in0(N__23213),
            .in1(N__16305),
            .in2(N__10422),
            .in3(N__10419),
            .lcout(n19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i10_LC_13_17_7 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i10_LC_13_17_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i10_LC_13_17_7 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \transmit_module.BRAM_ADDR__i10_LC_13_17_7  (
            .in0(N__16306),
            .in1(N__12756),
            .in2(N__23298),
            .in3(N__12744),
            .lcout(\transmit_module.TX_ADDR_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24208),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i9_3_lut_LC_13_18_2 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i9_3_lut_LC_13_18_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i9_3_lut_LC_13_18_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \transmit_module.mux_12_i9_3_lut_LC_13_18_2  (
            .in0(N__12427),
            .in1(N__20580),
            .in2(_gnd_net_),
            .in3(N__12405),
            .lcout(\transmit_module.n108 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_14_i9_3_lut_LC_13_18_3 .C_ON=1'b0;
    defparam \transmit_module.mux_14_i9_3_lut_LC_13_18_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_14_i9_3_lut_LC_13_18_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_14_i9_3_lut_LC_13_18_3  (
            .in0(N__14041),
            .in1(N__12426),
            .in2(_gnd_net_),
            .in3(N__12306),
            .lcout(\transmit_module.n139 ),
            .ltout(\transmit_module.n139_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1650_4_lut_LC_13_18_4 .C_ON=1'b0;
    defparam \transmit_module.i1650_4_lut_LC_13_18_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1650_4_lut_LC_13_18_4 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \transmit_module.i1650_4_lut_LC_13_18_4  (
            .in0(N__11438),
            .in1(N__23234),
            .in2(N__11427),
            .in3(N__16308),
            .lcout(n20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i11_3_lut_LC_13_18_5 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i11_3_lut_LC_13_18_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i11_3_lut_LC_13_18_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_12_i11_3_lut_LC_13_18_5  (
            .in0(N__20579),
            .in1(N__11202),
            .in2(_gnd_net_),
            .in3(N__12362),
            .lcout(\transmit_module.n106 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1644_4_lut_LC_13_19_0 .C_ON=1'b0;
    defparam \transmit_module.i1644_4_lut_LC_13_19_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1644_4_lut_LC_13_19_0 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \transmit_module.i1644_4_lut_LC_13_19_0  (
            .in0(N__16322),
            .in1(N__10952),
            .in2(N__23302),
            .in3(N__11190),
            .lcout(n26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i3_3_lut_LC_13_19_1 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i3_3_lut_LC_13_19_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i3_3_lut_LC_13_19_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_12_i3_3_lut_LC_13_19_1  (
            .in0(N__20590),
            .in1(N__10689),
            .in2(_gnd_net_),
            .in3(N__12107),
            .lcout(\transmit_module.n114 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_14_i4_3_lut_LC_13_19_2 .C_ON=1'b0;
    defparam \transmit_module.mux_14_i4_3_lut_LC_13_19_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_14_i4_3_lut_LC_13_19_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \transmit_module.mux_14_i4_3_lut_LC_13_19_2  (
            .in0(N__12075),
            .in1(N__14042),
            .in2(_gnd_net_),
            .in3(N__12048),
            .lcout(\transmit_module.n144 ),
            .ltout(\transmit_module.n144_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1645_4_lut_LC_13_19_3 .C_ON=1'b0;
    defparam \transmit_module.i1645_4_lut_LC_13_19_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1645_4_lut_LC_13_19_3 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \transmit_module.i1645_4_lut_LC_13_19_3  (
            .in0(N__23286),
            .in1(N__16323),
            .in2(N__10932),
            .in3(N__10700),
            .lcout(n25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i4_3_lut_LC_13_19_4 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i4_3_lut_LC_13_19_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i4_3_lut_LC_13_19_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_12_i4_3_lut_LC_13_19_4  (
            .in0(N__20591),
            .in1(N__11586),
            .in2(_gnd_net_),
            .in3(N__12073),
            .lcout(\transmit_module.n113 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.ADDR_Y_COMPONENT__i2_LC_13_19_5 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i2_LC_13_19_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i2_LC_13_19_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i2_LC_13_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12108),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23852),
            .ce(N__15390),
            .sr(N__23238));
    defparam \transmit_module.ADDR_Y_COMPONENT__i3_LC_13_19_6 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i3_LC_13_19_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i3_LC_13_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i3_LC_13_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12074),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23852),
            .ce(N__15390),
            .sr(N__23238));
    defparam \line_buffer.i2194_3_lut_LC_13_21_5 .C_ON=1'b0;
    defparam \line_buffer.i2194_3_lut_LC_13_21_5 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2194_3_lut_LC_13_21_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \line_buffer.i2194_3_lut_LC_13_21_5  (
            .in0(N__11580),
            .in1(N__11565),
            .in2(_gnd_net_),
            .in3(N__22832),
            .lcout(),
            .ltout(\line_buffer.n3531_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i7_LC_13_21_6 .C_ON=1'b0;
    defparam \line_buffer.dout_i7_LC_13_21_6 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i7_LC_13_21_6 .LUT_INIT=16'b1111101001000100;
    LogicCell40 \line_buffer.dout_i7_LC_13_21_6  (
            .in0(N__21294),
            .in1(N__11547),
            .in2(N__11535),
            .in3(N__11532),
            .lcout(TX_DATA_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23798),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.VGA_R__i8_LC_13_22_2 .C_ON=1'b0;
    defparam \transmit_module.VGA_R__i8_LC_13_22_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.VGA_R__i8_LC_13_22_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.VGA_R__i8_LC_13_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11526),
            .lcout(ADV_B_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23835),
            .ce(),
            .sr(N__22414));
    defparam \transmit_module.X_DELTA_PATTERN_i6_LC_14_9_3 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i6_LC_14_9_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i6_LC_14_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i6_LC_14_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13866),
            .lcout(\transmit_module.X_DELTA_PATTERN_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24333),
            .ce(N__18663),
            .sr(N__20492));
    defparam \transmit_module.X_DELTA_PATTERN_i12_LC_14_9_7 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i12_LC_14_9_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.X_DELTA_PATTERN_i12_LC_14_9_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i12_LC_14_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11622),
            .lcout(\transmit_module.X_DELTA_PATTERN_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24333),
            .ce(N__18663),
            .sr(N__20492));
    defparam \transmit_module.Y_DELTA_PATTERN_i24_LC_14_10_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i24_LC_14_10_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i24_LC_14_10_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i24_LC_14_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11457),
            .lcout(\transmit_module.Y_DELTA_PATTERN_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24331),
            .ce(N__20487),
            .sr(N__23197));
    defparam \transmit_module.Y_DELTA_PATTERN_i25_LC_14_10_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i25_LC_14_10_2 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i25_LC_14_10_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i25_LC_14_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11469),
            .lcout(\transmit_module.Y_DELTA_PATTERN_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24331),
            .ce(N__20487),
            .sr(N__23197));
    defparam \transmit_module.Y_DELTA_PATTERN_i19_LC_14_10_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i19_LC_14_10_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i19_LC_14_10_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i19_LC_14_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11652),
            .lcout(\transmit_module.Y_DELTA_PATTERN_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24331),
            .ce(N__20487),
            .sr(N__23197));
    defparam \transmit_module.Y_DELTA_PATTERN_i20_LC_14_10_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i20_LC_14_10_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i20_LC_14_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i20_LC_14_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11646),
            .lcout(\transmit_module.Y_DELTA_PATTERN_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24331),
            .ce(N__20487),
            .sr(N__23197));
    defparam \transmit_module.Y_DELTA_PATTERN_i21_LC_14_10_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i21_LC_14_10_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i21_LC_14_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i21_LC_14_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11640),
            .lcout(\transmit_module.Y_DELTA_PATTERN_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24331),
            .ce(N__20487),
            .sr(N__23197));
    defparam \transmit_module.Y_DELTA_PATTERN_i22_LC_14_10_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i22_LC_14_10_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i22_LC_14_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i22_LC_14_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11628),
            .lcout(\transmit_module.Y_DELTA_PATTERN_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24331),
            .ce(N__20487),
            .sr(N__23197));
    defparam \transmit_module.Y_DELTA_PATTERN_i23_LC_14_10_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i23_LC_14_10_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i23_LC_14_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i23_LC_14_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11634),
            .lcout(\transmit_module.Y_DELTA_PATTERN_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24331),
            .ce(N__20487),
            .sr(N__23197));
    defparam \transmit_module.X_DELTA_PATTERN_i13_LC_14_11_0 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i13_LC_14_11_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i13_LC_14_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i13_LC_14_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11613),
            .lcout(\transmit_module.X_DELTA_PATTERN_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24273),
            .ce(N__18655),
            .sr(N__20486));
    defparam \transmit_module.X_DELTA_PATTERN_i14_LC_14_11_1 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i14_LC_14_11_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.X_DELTA_PATTERN_i14_LC_14_11_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i14_LC_14_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18675),
            .lcout(\transmit_module.X_DELTA_PATTERN_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24273),
            .ce(N__18655),
            .sr(N__20486));
    defparam \transmit_module.X_DELTA_PATTERN_i3_LC_14_11_2 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i3_LC_14_11_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.X_DELTA_PATTERN_i3_LC_14_11_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i3_LC_14_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11592),
            .lcout(\transmit_module.X_DELTA_PATTERN_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24273),
            .ce(N__18655),
            .sr(N__20486));
    defparam \transmit_module.X_DELTA_PATTERN_i5_LC_14_11_4 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i5_LC_14_11_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.X_DELTA_PATTERN_i5_LC_14_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i5_LC_14_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11607),
            .lcout(\transmit_module.X_DELTA_PATTERN_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24273),
            .ce(N__18655),
            .sr(N__20486));
    defparam \transmit_module.X_DELTA_PATTERN_i4_LC_14_11_7 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i4_LC_14_11_7 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i4_LC_14_11_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i4_LC_14_11_7  (
            .in0(N__11598),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.X_DELTA_PATTERN_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24273),
            .ce(N__18655),
            .sr(N__20486));
    defparam \transmit_module.video_signal_controller.i480_2_lut_LC_14_12_0 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i480_2_lut_LC_14_12_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i480_2_lut_LC_14_12_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \transmit_module.video_signal_controller.i480_2_lut_LC_14_12_0  (
            .in0(_gnd_net_),
            .in1(N__11992),
            .in2(_gnd_net_),
            .in3(N__12025),
            .lcout(),
            .ltout(\transmit_module.video_signal_controller.n6_adj_622_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_4_lut_adj_28_LC_14_12_1 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_4_lut_adj_28_LC_14_12_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_4_lut_adj_28_LC_14_12_1 .LUT_INIT=16'b1111111110101000;
    LogicCell40 \transmit_module.video_signal_controller.i1_4_lut_adj_28_LC_14_12_1  (
            .in0(N__11739),
            .in1(N__11758),
            .in2(N__11763),
            .in3(N__11684),
            .lcout(\transmit_module.video_signal_controller.VGA_VISIBLE_N_588 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i2180_3_lut_LC_14_12_3 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i2180_3_lut_LC_14_12_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i2180_3_lut_LC_14_12_3 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \transmit_module.video_signal_controller.i2180_3_lut_LC_14_12_3  (
            .in0(N__11740),
            .in1(N__11759),
            .in2(_gnd_net_),
            .in3(N__11685),
            .lcout(\transmit_module.video_signal_controller.n3517 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i2_3_lut_LC_14_12_4 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i2_3_lut_LC_14_12_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i2_3_lut_LC_14_12_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \transmit_module.video_signal_controller.i2_3_lut_LC_14_12_4  (
            .in0(N__11757),
            .in1(N__11991),
            .in2(_gnd_net_),
            .in3(N__12024),
            .lcout(),
            .ltout(\transmit_module.video_signal_controller.n3482_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i2_4_lut_LC_14_12_5 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i2_4_lut_LC_14_12_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i2_4_lut_LC_14_12_5 .LUT_INIT=16'b1010100000000000;
    LogicCell40 \transmit_module.video_signal_controller.i2_4_lut_LC_14_12_5  (
            .in0(N__11717),
            .in1(N__11741),
            .in2(N__11721),
            .in3(N__11702),
            .lcout(\transmit_module.video_signal_controller.n3461 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_2_lut_3_lut_LC_14_12_6 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_2_lut_3_lut_LC_14_12_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_2_lut_3_lut_LC_14_12_6 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \transmit_module.video_signal_controller.i1_2_lut_3_lut_LC_14_12_6  (
            .in0(N__13753),
            .in1(N__13729),
            .in2(_gnd_net_),
            .in3(N__11716),
            .lcout(),
            .ltout(\transmit_module.video_signal_controller.n6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i4_4_lut_LC_14_12_7 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i4_4_lut_LC_14_12_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i4_4_lut_LC_14_12_7 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \transmit_module.video_signal_controller.i4_4_lut_LC_14_12_7  (
            .in0(N__13690),
            .in1(N__11701),
            .in2(N__11688),
            .in3(N__13709),
            .lcout(\transmit_module.video_signal_controller.n2016 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.VGA_VISIBLE_Y_64_LC_14_13_0 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.VGA_VISIBLE_Y_64_LC_14_13_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_VISIBLE_Y_64_LC_14_13_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_VISIBLE_Y_64_LC_14_13_0  (
            .in0(_gnd_net_),
            .in1(N__12272),
            .in2(_gnd_net_),
            .in3(N__13673),
            .lcout(\transmit_module.VGA_VISIBLE_Y ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24272),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_2_lut_LC_14_13_1 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_2_lut_LC_14_13_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_2_lut_LC_14_13_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \transmit_module.video_signal_controller.i1_2_lut_LC_14_13_1  (
            .in0(_gnd_net_),
            .in1(N__11675),
            .in2(_gnd_net_),
            .in3(N__11663),
            .lcout(\transmit_module.video_signal_controller.n3375 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i124_2_lut_4_lut_LC_14_13_3 .C_ON=1'b0;
    defparam \transmit_module.i124_2_lut_4_lut_LC_14_13_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i124_2_lut_4_lut_LC_14_13_3 .LUT_INIT=16'b1100110011101100;
    LogicCell40 \transmit_module.i124_2_lut_4_lut_LC_14_13_3  (
            .in0(N__11786),
            .in1(N__23025),
            .in2(N__11859),
            .in3(N__11814),
            .lcout(\transmit_module.n2206 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.VGA_VS_67_LC_14_13_4 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.VGA_VS_67_LC_14_13_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_VS_67_LC_14_13_4 .LUT_INIT=16'b0001000100010000;
    LogicCell40 \transmit_module.video_signal_controller.VGA_VS_67_LC_14_13_4  (
            .in0(N__12033),
            .in1(N__12006),
            .in2(N__12000),
            .in3(N__11973),
            .lcout(ADV_VSYNC_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24272),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i124_2_lut_4_lut_rep_23_LC_14_13_5 .C_ON=1'b0;
    defparam \transmit_module.i124_2_lut_4_lut_rep_23_LC_14_13_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i124_2_lut_4_lut_rep_23_LC_14_13_5 .LUT_INIT=16'b1100110011101100;
    LogicCell40 \transmit_module.i124_2_lut_4_lut_rep_23_LC_14_13_5  (
            .in0(N__11785),
            .in1(N__23024),
            .in2(N__11858),
            .in3(N__11813),
            .lcout(\transmit_module.n3679 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1729_4_lut_LC_14_13_6 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1729_4_lut_LC_14_13_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1729_4_lut_LC_14_13_6 .LUT_INIT=16'b1100110010000000;
    LogicCell40 \transmit_module.video_signal_controller.i1729_4_lut_LC_14_13_6  (
            .in0(N__11961),
            .in1(N__11955),
            .in2(N__11928),
            .in3(N__11913),
            .lcout(),
            .ltout(\transmit_module.video_signal_controller.n2972_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1735_4_lut_LC_14_13_7 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1735_4_lut_LC_14_13_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1735_4_lut_LC_14_13_7 .LUT_INIT=16'b1110111011101010;
    LogicCell40 \transmit_module.video_signal_controller.i1735_4_lut_LC_14_13_7  (
            .in0(N__12255),
            .in1(N__12199),
            .in2(N__11907),
            .in3(N__12162),
            .lcout(\transmit_module.video_signal_controller.n2047 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i1_3_lut_LC_14_14_0 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i1_3_lut_LC_14_14_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i1_3_lut_LC_14_14_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_12_i1_3_lut_LC_14_14_0  (
            .in0(N__20628),
            .in1(N__12471),
            .in2(_gnd_net_),
            .in3(N__13909),
            .lcout(\transmit_module.n116 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i2_3_lut_rep_19_LC_14_14_1 .C_ON=1'b0;
    defparam \transmit_module.i2_3_lut_rep_19_LC_14_14_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i2_3_lut_rep_19_LC_14_14_1 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \transmit_module.i2_3_lut_rep_19_LC_14_14_1  (
            .in0(N__11850),
            .in1(N__11812),
            .in2(_gnd_net_),
            .in3(N__11784),
            .lcout(\transmit_module.n3675 ),
            .ltout(\transmit_module.n3675_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i2_3_lut_LC_14_14_2 .C_ON=1'b0;
    defparam \transmit_module.i2_3_lut_LC_14_14_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i2_3_lut_LC_14_14_2 .LUT_INIT=16'b1111111111111010;
    LogicCell40 \transmit_module.i2_3_lut_LC_14_14_2  (
            .in0(N__23091),
            .in1(_gnd_net_),
            .in2(N__11766),
            .in3(N__14026),
            .lcout(\transmit_module.n2084 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i2_2_lut_LC_14_14_3 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i2_2_lut_LC_14_14_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i2_2_lut_LC_14_14_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \transmit_module.video_signal_controller.i2_2_lut_LC_14_14_3  (
            .in0(_gnd_net_),
            .in1(N__12257),
            .in2(_gnd_net_),
            .in3(N__12160),
            .lcout(),
            .ltout(\transmit_module.video_signal_controller.n6_adj_623_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i2_4_lut_adj_35_LC_14_14_4 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i2_4_lut_adj_35_LC_14_14_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i2_4_lut_adj_35_LC_14_14_4 .LUT_INIT=16'b1111111000000000;
    LogicCell40 \transmit_module.video_signal_controller.i2_4_lut_adj_35_LC_14_14_4  (
            .in0(N__12201),
            .in1(N__12210),
            .in2(N__12276),
            .in3(N__12273),
            .lcout(),
            .ltout(\transmit_module.video_signal_controller.n7_adj_624_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.VGA_VISIBLE_65_LC_14_14_5 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.VGA_VISIBLE_65_LC_14_14_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_VISIBLE_65_LC_14_14_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \transmit_module.video_signal_controller.VGA_VISIBLE_65_LC_14_14_5  (
            .in0(N__12258),
            .in1(N__13674),
            .in2(N__12213),
            .in3(N__12123),
            .lcout(\transmit_module.VGA_VISIBLE ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24223),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1696_4_lut_LC_14_14_6 .C_ON=1'b0;
    defparam \transmit_module.i1696_4_lut_LC_14_14_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1696_4_lut_LC_14_14_6 .LUT_INIT=16'b1111011111110100;
    LogicCell40 \transmit_module.i1696_4_lut_LC_14_14_6  (
            .in0(N__20629),
            .in1(N__16264),
            .in2(N__23223),
            .in3(N__14025),
            .lcout(\transmit_module.n2070 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1771_3_lut_LC_14_14_7 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1771_3_lut_LC_14_14_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1771_3_lut_LC_14_14_7 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \transmit_module.video_signal_controller.i1771_3_lut_LC_14_14_7  (
            .in0(N__12209),
            .in1(N__12200),
            .in2(_gnd_net_),
            .in3(N__12161),
            .lcout(\transmit_module.video_signal_controller.n3014 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_2_lut_LC_14_15_0 .C_ON=1'b1;
    defparam \transmit_module.add_13_2_lut_LC_14_15_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_2_lut_LC_14_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_2_lut_LC_14_15_0  (
            .in0(_gnd_net_),
            .in1(N__18686),
            .in2(N__13913),
            .in3(_gnd_net_),
            .lcout(\transmit_module.n132 ),
            .ltout(),
            .carryin(bfn_14_15_0_),
            .carryout(\transmit_module.n3159 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_3_lut_LC_14_15_1 .C_ON=1'b1;
    defparam \transmit_module.add_13_3_lut_LC_14_15_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_3_lut_LC_14_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_3_lut_LC_14_15_1  (
            .in0(_gnd_net_),
            .in1(N__12453),
            .in2(_gnd_net_),
            .in3(N__12111),
            .lcout(\transmit_module.n131 ),
            .ltout(),
            .carryin(\transmit_module.n3159 ),
            .carryout(\transmit_module.n3160 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_4_lut_LC_14_15_2 .C_ON=1'b1;
    defparam \transmit_module.add_13_4_lut_LC_14_15_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_4_lut_LC_14_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_4_lut_LC_14_15_2  (
            .in0(_gnd_net_),
            .in1(N__12100),
            .in2(_gnd_net_),
            .in3(N__12078),
            .lcout(\transmit_module.n130 ),
            .ltout(),
            .carryin(\transmit_module.n3160 ),
            .carryout(\transmit_module.n3161 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_5_lut_LC_14_15_3 .C_ON=1'b1;
    defparam \transmit_module.add_13_5_lut_LC_14_15_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_5_lut_LC_14_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_5_lut_LC_14_15_3  (
            .in0(_gnd_net_),
            .in1(N__12064),
            .in2(_gnd_net_),
            .in3(N__12036),
            .lcout(\transmit_module.n129 ),
            .ltout(),
            .carryin(\transmit_module.n3161 ),
            .carryout(\transmit_module.n3162 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_6_lut_LC_14_15_4 .C_ON=1'b1;
    defparam \transmit_module.add_13_6_lut_LC_14_15_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_6_lut_LC_14_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_6_lut_LC_14_15_4  (
            .in0(_gnd_net_),
            .in1(N__15513),
            .in2(_gnd_net_),
            .in3(N__12330),
            .lcout(\transmit_module.n128 ),
            .ltout(),
            .carryin(\transmit_module.n3162 ),
            .carryout(\transmit_module.n3163 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_7_lut_LC_14_15_5 .C_ON=1'b1;
    defparam \transmit_module.add_13_7_lut_LC_14_15_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_7_lut_LC_14_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_7_lut_LC_14_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12399),
            .in3(N__12315),
            .lcout(\transmit_module.n127 ),
            .ltout(),
            .carryin(\transmit_module.n3163 ),
            .carryout(\transmit_module.n3164 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_8_lut_LC_14_15_6 .C_ON=1'b1;
    defparam \transmit_module.add_13_8_lut_LC_14_15_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_8_lut_LC_14_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_8_lut_LC_14_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15439),
            .in3(N__12312),
            .lcout(\transmit_module.n126 ),
            .ltout(),
            .carryin(\transmit_module.n3164 ),
            .carryout(\transmit_module.n3165 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_9_lut_LC_14_15_7 .C_ON=1'b1;
    defparam \transmit_module.add_13_9_lut_LC_14_15_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_9_lut_LC_14_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_9_lut_LC_14_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15477),
            .in3(N__12309),
            .lcout(\transmit_module.n125 ),
            .ltout(),
            .carryin(\transmit_module.n3165 ),
            .carryout(\transmit_module.n3166 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_10_lut_LC_14_16_0 .C_ON=1'b1;
    defparam \transmit_module.add_13_10_lut_LC_14_16_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_10_lut_LC_14_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_10_lut_LC_14_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12429),
            .in3(N__12297),
            .lcout(\transmit_module.n124 ),
            .ltout(),
            .carryin(bfn_14_16_0_),
            .carryout(\transmit_module.n3167 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_11_lut_LC_14_16_1 .C_ON=1'b1;
    defparam \transmit_module.add_13_11_lut_LC_14_16_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_11_lut_LC_14_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_11_lut_LC_14_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12501),
            .in3(N__12288),
            .lcout(\transmit_module.n123 ),
            .ltout(),
            .carryin(\transmit_module.n3167 ),
            .carryout(\transmit_module.n3168 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_12_lut_LC_14_16_2 .C_ON=1'b1;
    defparam \transmit_module.add_13_12_lut_LC_14_16_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_12_lut_LC_14_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_12_lut_LC_14_16_2  (
            .in0(_gnd_net_),
            .in1(N__12360),
            .in2(_gnd_net_),
            .in3(N__12285),
            .lcout(\transmit_module.n122 ),
            .ltout(),
            .carryin(\transmit_module.n3168 ),
            .carryout(\transmit_module.n3169 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_13_lut_LC_14_16_3 .C_ON=1'b1;
    defparam \transmit_module.add_13_13_lut_LC_14_16_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_13_lut_LC_14_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_13_lut_LC_14_16_3  (
            .in0(_gnd_net_),
            .in1(N__22763),
            .in2(_gnd_net_),
            .in3(N__12282),
            .lcout(\transmit_module.n121 ),
            .ltout(),
            .carryin(\transmit_module.n3169 ),
            .carryout(\transmit_module.n3170 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_14_lut_LC_14_16_4 .C_ON=1'b1;
    defparam \transmit_module.add_13_14_lut_LC_14_16_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_14_lut_LC_14_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_14_lut_LC_14_16_4  (
            .in0(_gnd_net_),
            .in1(N__21439),
            .in2(_gnd_net_),
            .in3(N__12279),
            .lcout(\transmit_module.n120 ),
            .ltout(),
            .carryin(\transmit_module.n3170 ),
            .carryout(\transmit_module.n3171 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_15_lut_LC_14_16_5 .C_ON=1'b0;
    defparam \transmit_module.add_13_15_lut_LC_14_16_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_15_lut_LC_14_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_15_lut_LC_14_16_5  (
            .in0(_gnd_net_),
            .in1(N__21228),
            .in2(_gnd_net_),
            .in3(N__12504),
            .lcout(\transmit_module.n119 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.ADDR_Y_COMPONENT__i9_LC_14_16_6 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i9_LC_14_16_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i9_LC_14_16_6 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i9_LC_14_16_6  (
            .in0(_gnd_net_),
            .in1(N__12498),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24146),
            .ce(N__15397),
            .sr(N__23140));
    defparam \transmit_module.ADDR_Y_COMPONENT__i0_LC_14_17_0 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i0_LC_14_17_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i0_LC_14_17_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i0_LC_14_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13914),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24066),
            .ce(N__15389),
            .sr(N__23239));
    defparam \transmit_module.ADDR_Y_COMPONENT__i1_LC_14_17_1 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i1_LC_14_17_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i1_LC_14_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i1_LC_14_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12462),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24066),
            .ce(N__15389),
            .sr(N__23239));
    defparam \transmit_module.ADDR_Y_COMPONENT__i8_LC_14_17_2 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i8_LC_14_17_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i8_LC_14_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i8_LC_14_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12428),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24066),
            .ce(N__15389),
            .sr(N__23239));
    defparam \transmit_module.ADDR_Y_COMPONENT__i12_LC_14_17_4 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i12_LC_14_17_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i12_LC_14_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i12_LC_14_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21484),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24066),
            .ce(N__15389),
            .sr(N__23239));
    defparam \transmit_module.ADDR_Y_COMPONENT__i13_LC_14_17_5 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i13_LC_14_17_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i13_LC_14_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i13_LC_14_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21270),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24066),
            .ce(N__15389),
            .sr(N__23239));
    defparam \transmit_module.ADDR_Y_COMPONENT__i5_LC_14_17_7 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i5_LC_14_17_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i5_LC_14_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i5_LC_14_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12398),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24066),
            .ce(N__15389),
            .sr(N__23239));
    defparam \transmit_module.mux_14_i11_3_lut_LC_14_18_1 .C_ON=1'b0;
    defparam \transmit_module.mux_14_i11_3_lut_LC_14_18_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_14_i11_3_lut_LC_14_18_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_14_i11_3_lut_LC_14_18_1  (
            .in0(N__14039),
            .in1(N__12361),
            .in2(_gnd_net_),
            .in3(N__12339),
            .lcout(\transmit_module.n137 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i7_3_lut_LC_14_18_5 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i7_3_lut_LC_14_18_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i7_3_lut_LC_14_18_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_12_i7_3_lut_LC_14_18_5  (
            .in0(N__20604),
            .in1(N__15408),
            .in2(_gnd_net_),
            .in3(N__15444),
            .lcout(\transmit_module.n110 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i8_3_lut_LC_14_18_6 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i8_3_lut_LC_14_18_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i8_3_lut_LC_14_18_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_12_i8_3_lut_LC_14_18_6  (
            .in0(N__20605),
            .in1(N__15450),
            .in2(_gnd_net_),
            .in3(N__15488),
            .lcout(\transmit_module.n109 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1648_4_lut_LC_14_19_0 .C_ON=1'b0;
    defparam \transmit_module.i1648_4_lut_LC_14_19_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1648_4_lut_LC_14_19_0 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \transmit_module.i1648_4_lut_LC_14_19_0  (
            .in0(N__16299),
            .in1(N__13778),
            .in2(N__23297),
            .in3(N__13797),
            .lcout(n22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i5_3_lut_LC_14_19_1 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i5_3_lut_LC_14_19_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i5_3_lut_LC_14_19_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_12_i5_3_lut_LC_14_19_1  (
            .in0(N__20625),
            .in1(N__15495),
            .in2(_gnd_net_),
            .in3(N__15525),
            .lcout(\transmit_module.n112 ),
            .ltout(\transmit_module.n112_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1646_4_lut_LC_14_19_2 .C_ON=1'b0;
    defparam \transmit_module.i1646_4_lut_LC_14_19_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1646_4_lut_LC_14_19_2 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \transmit_module.i1646_4_lut_LC_14_19_2  (
            .in0(N__16298),
            .in1(N__23233),
            .in2(N__13242),
            .in3(N__13956),
            .lcout(n24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_14_i8_3_lut_LC_14_19_5 .C_ON=1'b0;
    defparam \transmit_module.mux_14_i8_3_lut_LC_14_19_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_14_i8_3_lut_LC_14_19_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_14_i8_3_lut_LC_14_19_5  (
            .in0(N__14040),
            .in1(N__15487),
            .in2(_gnd_net_),
            .in3(N__13029),
            .lcout(\transmit_module.n140 ),
            .ltout(\transmit_module.n140_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1649_4_lut_LC_14_19_6 .C_ON=1'b0;
    defparam \transmit_module.i1649_4_lut_LC_14_19_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1649_4_lut_LC_14_19_6 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \transmit_module.i1649_4_lut_LC_14_19_6  (
            .in0(N__16300),
            .in1(N__23229),
            .in2(N__13008),
            .in3(N__12995),
            .lcout(n21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1652_4_lut_LC_14_19_7 .C_ON=1'b0;
    defparam \transmit_module.i1652_4_lut_LC_14_19_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1652_4_lut_LC_14_19_7 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \transmit_module.i1652_4_lut_LC_14_19_7  (
            .in0(N__16321),
            .in1(N__12755),
            .in2(N__23301),
            .in3(N__12743),
            .lcout(n18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1141_1_lut_LC_14_20_1 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1141_1_lut_LC_14_20_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1141_1_lut_LC_14_20_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \transmit_module.video_signal_controller.i1141_1_lut_LC_14_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14043),
            .lcout(\transmit_module.n2385 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.BUFFER_0__i4_LC_15_1_3 .C_ON=1'b0;
    defparam \tvp_video_buffer.BUFFER_0__i4_LC_15_1_3 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.BUFFER_0__i4_LC_15_1_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \tvp_video_buffer.BUFFER_0__i4_LC_15_1_3  (
            .in0(N__13635),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\tvp_video_buffer.BUFFER_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21926),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_vs_buffer.BUFFER_0__i1_LC_15_7_2 .C_ON=1'b0;
    defparam \tvp_vs_buffer.BUFFER_0__i1_LC_15_7_2 .SEQ_MODE=4'b1000;
    defparam \tvp_vs_buffer.BUFFER_0__i1_LC_15_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_vs_buffer.BUFFER_0__i1_LC_15_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13610),
            .lcout(\tvp_vs_buffer.BUFFER_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21933),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_vs_buffer.BUFFER_0__i2_LC_15_7_5 .C_ON=1'b0;
    defparam \tvp_vs_buffer.BUFFER_0__i2_LC_15_7_5 .SEQ_MODE=4'b1000;
    defparam \tvp_vs_buffer.BUFFER_0__i2_LC_15_7_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_vs_buffer.BUFFER_0__i2_LC_15_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13593),
            .lcout(\tvp_vs_buffer.BUFFER_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21933),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_vs_buffer.BUFFER_0__i3_LC_15_8_5 .C_ON=1'b0;
    defparam \tvp_vs_buffer.BUFFER_0__i3_LC_15_8_5 .SEQ_MODE=4'b1000;
    defparam \tvp_vs_buffer.BUFFER_0__i3_LC_15_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_vs_buffer.BUFFER_0__i3_LC_15_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13587),
            .lcout(\tvp_vs_buffer.BUFFER_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21936),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.sync_wd.i2_2_lut_LC_15_9_1 .C_ON=1'b0;
    defparam \receive_module.sync_wd.i2_2_lut_LC_15_9_1 .SEQ_MODE=4'b0000;
    defparam \receive_module.sync_wd.i2_2_lut_LC_15_9_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \receive_module.sync_wd.i2_2_lut_LC_15_9_1  (
            .in0(_gnd_net_),
            .in1(N__19873),
            .in2(_gnd_net_),
            .in3(N__21007),
            .lcout(),
            .ltout(\receive_module.sync_wd.n6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.sync_wd.i1_4_lut_LC_15_9_2 .C_ON=1'b0;
    defparam \receive_module.sync_wd.i1_4_lut_LC_15_9_2 .SEQ_MODE=4'b0000;
    defparam \receive_module.sync_wd.i1_4_lut_LC_15_9_2 .LUT_INIT=16'b1111111100000001;
    LogicCell40 \receive_module.sync_wd.i1_4_lut_LC_15_9_2  (
            .in0(N__21692),
            .in1(N__13549),
            .in2(N__13476),
            .in3(N__19668),
            .lcout(),
            .ltout(\receive_module.sync_wd.n4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.sync_wd.SYNC_BAD_16_LC_15_9_3 .C_ON=1'b0;
    defparam \receive_module.sync_wd.SYNC_BAD_16_LC_15_9_3 .SEQ_MODE=4'b1000;
    defparam \receive_module.sync_wd.SYNC_BAD_16_LC_15_9_3 .LUT_INIT=16'b1100111000000000;
    LogicCell40 \receive_module.sync_wd.SYNC_BAD_16_LC_15_9_3  (
            .in0(N__13470),
            .in1(N__18163),
            .in2(N__13473),
            .in3(N__20096),
            .lcout(DEBUG_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21941),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.sync_wd.old_visible_17_LC_15_9_4 .C_ON=1'b0;
    defparam \receive_module.sync_wd.old_visible_17_LC_15_9_4 .SEQ_MODE=4'b1000;
    defparam \receive_module.sync_wd.old_visible_17_LC_15_9_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \receive_module.sync_wd.old_visible_17_LC_15_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19669),
            .lcout(\receive_module.sync_wd.old_visible ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21941),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.X_243__i0_LC_15_10_0 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_243__i0_LC_15_10_0 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_243__i0_LC_15_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_243__i0_LC_15_10_0  (
            .in0(_gnd_net_),
            .in1(N__15705),
            .in2(_gnd_net_),
            .in3(N__13464),
            .lcout(\receive_module.rx_counter.X_0 ),
            .ltout(),
            .carryin(bfn_15_10_0_),
            .carryout(\receive_module.rx_counter.n3207 ),
            .clk(N__21947),
            .ce(),
            .sr(N__15746));
    defparam \receive_module.rx_counter.X_243__i1_LC_15_10_1 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_243__i1_LC_15_10_1 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_243__i1_LC_15_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_243__i1_LC_15_10_1  (
            .in0(_gnd_net_),
            .in1(N__15729),
            .in2(_gnd_net_),
            .in3(N__13662),
            .lcout(\receive_module.rx_counter.X_1 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3207 ),
            .carryout(\receive_module.rx_counter.n3208 ),
            .clk(N__21947),
            .ce(),
            .sr(N__15746));
    defparam \receive_module.rx_counter.X_243__i2_LC_15_10_2 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_243__i2_LC_15_10_2 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_243__i2_LC_15_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_243__i2_LC_15_10_2  (
            .in0(_gnd_net_),
            .in1(N__15717),
            .in2(_gnd_net_),
            .in3(N__13659),
            .lcout(\receive_module.rx_counter.X_2 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3208 ),
            .carryout(\receive_module.rx_counter.n3209 ),
            .clk(N__21947),
            .ce(),
            .sr(N__15746));
    defparam \receive_module.rx_counter.X_243__i3_LC_15_10_3 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_243__i3_LC_15_10_3 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_243__i3_LC_15_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_243__i3_LC_15_10_3  (
            .in0(_gnd_net_),
            .in1(N__16003),
            .in2(_gnd_net_),
            .in3(N__13656),
            .lcout(\receive_module.rx_counter.X_3 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3209 ),
            .carryout(\receive_module.rx_counter.n3210 ),
            .clk(N__21947),
            .ce(),
            .sr(N__15746));
    defparam \receive_module.rx_counter.X_243__i4_LC_15_10_4 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_243__i4_LC_15_10_4 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_243__i4_LC_15_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_243__i4_LC_15_10_4  (
            .in0(_gnd_net_),
            .in1(N__15946),
            .in2(_gnd_net_),
            .in3(N__13653),
            .lcout(\receive_module.rx_counter.X_4 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3210 ),
            .carryout(\receive_module.rx_counter.n3211 ),
            .clk(N__21947),
            .ce(),
            .sr(N__15746));
    defparam \receive_module.rx_counter.X_243__i5_LC_15_10_5 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_243__i5_LC_15_10_5 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_243__i5_LC_15_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_243__i5_LC_15_10_5  (
            .in0(_gnd_net_),
            .in1(N__15976),
            .in2(_gnd_net_),
            .in3(N__13650),
            .lcout(\receive_module.rx_counter.X_5 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3211 ),
            .carryout(\receive_module.rx_counter.n3212 ),
            .clk(N__21947),
            .ce(),
            .sr(N__15746));
    defparam \receive_module.rx_counter.X_243__i6_LC_15_10_6 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_243__i6_LC_15_10_6 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_243__i6_LC_15_10_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_243__i6_LC_15_10_6  (
            .in0(_gnd_net_),
            .in1(N__15871),
            .in2(_gnd_net_),
            .in3(N__13647),
            .lcout(\receive_module.rx_counter.X_6 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3212 ),
            .carryout(\receive_module.rx_counter.n3213 ),
            .clk(N__21947),
            .ce(),
            .sr(N__15746));
    defparam \receive_module.rx_counter.X_243__i7_LC_15_10_7 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_243__i7_LC_15_10_7 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_243__i7_LC_15_10_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_243__i7_LC_15_10_7  (
            .in0(_gnd_net_),
            .in1(N__15901),
            .in2(_gnd_net_),
            .in3(N__13644),
            .lcout(\receive_module.rx_counter.X_7 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3213 ),
            .carryout(\receive_module.rx_counter.n3214 ),
            .clk(N__21947),
            .ce(),
            .sr(N__15746));
    defparam \receive_module.rx_counter.X_243__i8_LC_15_11_0 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_243__i8_LC_15_11_0 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_243__i8_LC_15_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_243__i8_LC_15_11_0  (
            .in0(_gnd_net_),
            .in1(N__15842),
            .in2(_gnd_net_),
            .in3(N__13641),
            .lcout(\receive_module.rx_counter.X_8 ),
            .ltout(),
            .carryin(bfn_15_11_0_),
            .carryout(\receive_module.rx_counter.n3215 ),
            .clk(N__21952),
            .ce(),
            .sr(N__15750));
    defparam \receive_module.rx_counter.X_243__i9_LC_15_11_1 .C_ON=1'b0;
    defparam \receive_module.rx_counter.X_243__i9_LC_15_11_1 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_243__i9_LC_15_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_243__i9_LC_15_11_1  (
            .in0(_gnd_net_),
            .in1(N__15824),
            .in2(_gnd_net_),
            .in3(N__13638),
            .lcout(\receive_module.rx_counter.X_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21952),
            .ce(),
            .sr(N__15750));
    defparam \receive_module.rx_counter.old_VS_52_LC_15_12_2 .C_ON=1'b0;
    defparam \receive_module.rx_counter.old_VS_52_LC_15_12_2 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.old_VS_52_LC_15_12_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \receive_module.rx_counter.old_VS_52_LC_15_12_2  (
            .in0(N__20067),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\receive_module.rx_counter.old_VS ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21955),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i2_2_lut_adj_25_LC_15_12_4 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i2_2_lut_adj_25_LC_15_12_4 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i2_2_lut_adj_25_LC_15_12_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \receive_module.rx_counter.i2_2_lut_adj_25_LC_15_12_4  (
            .in0(_gnd_net_),
            .in1(N__16004),
            .in2(_gnd_net_),
            .in3(N__15977),
            .lcout(\receive_module.rx_counter.n7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i131_2_lut_rep_16_2_lut_LC_15_12_5 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i131_2_lut_rep_16_2_lut_LC_15_12_5 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i131_2_lut_rep_16_2_lut_LC_15_12_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \receive_module.rx_counter.i131_2_lut_rep_16_2_lut_LC_15_12_5  (
            .in0(_gnd_net_),
            .in1(N__18998),
            .in2(_gnd_net_),
            .in3(N__20066),
            .lcout(\receive_module.rx_counter.n3672 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_vs_buffer.WIRE_OUT_0__9_LC_15_12_6 .C_ON=1'b0;
    defparam \tvp_vs_buffer.WIRE_OUT_0__9_LC_15_12_6 .SEQ_MODE=4'b1000;
    defparam \tvp_vs_buffer.WIRE_OUT_0__9_LC_15_12_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_vs_buffer.WIRE_OUT_0__9_LC_15_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13767),
            .lcout(TVP_VSYNC_buff),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21955),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i1_2_lut_adj_24_LC_15_12_7 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i1_2_lut_adj_24_LC_15_12_7 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i1_2_lut_adj_24_LC_15_12_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \receive_module.rx_counter.i1_2_lut_adj_24_LC_15_12_7  (
            .in0(_gnd_net_),
            .in1(N__15950),
            .in2(_gnd_net_),
            .in3(N__15872),
            .lcout(\receive_module.rx_counter.n6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.O_VS_I_0_1_lut_rep_18_LC_15_13_2 .C_ON=1'b0;
    defparam \receive_module.rx_counter.O_VS_I_0_1_lut_rep_18_LC_15_13_2 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.O_VS_I_0_1_lut_rep_18_LC_15_13_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \receive_module.rx_counter.O_VS_I_0_1_lut_rep_18_LC_15_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20056),
            .lcout(\receive_module.n3674 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_17_LC_15_13_3 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_17_LC_15_13_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_17_LC_15_13_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \transmit_module.video_signal_controller.i1_2_lut_rep_17_LC_15_13_3  (
            .in0(_gnd_net_),
            .in1(N__13758),
            .in2(_gnd_net_),
            .in3(N__13736),
            .lcout(),
            .ltout(\transmit_module.video_signal_controller.n3673_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_4_lut_LC_15_13_4 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_4_lut_LC_15_13_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_4_lut_LC_15_13_4 .LUT_INIT=16'b1111111011110000;
    LogicCell40 \transmit_module.video_signal_controller.i1_4_lut_LC_15_13_4  (
            .in0(N__13716),
            .in1(N__13710),
            .in2(N__13698),
            .in3(N__13695),
            .lcout(\transmit_module.video_signal_controller.n3379 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.X_DELTA_PATTERN_i0_LC_15_14_0 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i0_LC_15_14_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i0_LC_15_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i0_LC_15_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13809),
            .lcout(\transmit_module.X_DELTA_PATTERN_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24250),
            .ce(N__18645),
            .sr(N__20419));
    defparam \transmit_module.X_DELTA_PATTERN_i8_LC_15_14_1 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i8_LC_15_14_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.X_DELTA_PATTERN_i8_LC_15_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i8_LC_15_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13845),
            .lcout(\transmit_module.X_DELTA_PATTERN_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24250),
            .ce(N__18645),
            .sr(N__20419));
    defparam \transmit_module.X_DELTA_PATTERN_i7_LC_15_14_2 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i7_LC_15_14_2 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i7_LC_15_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i7_LC_15_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13872),
            .lcout(\transmit_module.X_DELTA_PATTERN_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24250),
            .ce(N__18645),
            .sr(N__20419));
    defparam \transmit_module.X_DELTA_PATTERN_i2_LC_15_14_3 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i2_LC_15_14_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i2_LC_15_14_3 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i2_LC_15_14_3  (
            .in0(_gnd_net_),
            .in1(N__13854),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.X_DELTA_PATTERN_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24250),
            .ce(N__18645),
            .sr(N__20419));
    defparam \transmit_module.X_DELTA_PATTERN_i9_LC_15_14_4 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i9_LC_15_14_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i9_LC_15_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i9_LC_15_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13839),
            .lcout(\transmit_module.X_DELTA_PATTERN_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24250),
            .ce(N__18645),
            .sr(N__20419));
    defparam \transmit_module.X_DELTA_PATTERN_i10_LC_15_14_5 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i10_LC_15_14_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.X_DELTA_PATTERN_i10_LC_15_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i10_LC_15_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13821),
            .lcout(\transmit_module.X_DELTA_PATTERN_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24250),
            .ce(N__18645),
            .sr(N__20419));
    defparam \transmit_module.X_DELTA_PATTERN_i11_LC_15_14_6 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i11_LC_15_14_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i11_LC_15_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i11_LC_15_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13833),
            .lcout(\transmit_module.X_DELTA_PATTERN_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24250),
            .ce(N__18645),
            .sr(N__20419));
    defparam \transmit_module.X_DELTA_PATTERN_i1_LC_15_14_7 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i1_LC_15_14_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.X_DELTA_PATTERN_i1_LC_15_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i1_LC_15_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13815),
            .lcout(\transmit_module.X_DELTA_PATTERN_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24250),
            .ce(N__18645),
            .sr(N__20419));
    defparam \transmit_module.mux_14_i7_3_lut_LC_15_15_0 .C_ON=1'b0;
    defparam \transmit_module.mux_14_i7_3_lut_LC_15_15_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_14_i7_3_lut_LC_15_15_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_14_i7_3_lut_LC_15_15_0  (
            .in0(N__14001),
            .in1(N__15432),
            .in2(_gnd_net_),
            .in3(N__13803),
            .lcout(\transmit_module.n141 ),
            .ltout(\transmit_module.n141_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i6_LC_15_15_1 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i6_LC_15_15_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i6_LC_15_15_1 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \transmit_module.BRAM_ADDR__i6_LC_15_15_1  (
            .in0(N__23143),
            .in1(N__16238),
            .in2(N__13785),
            .in3(N__13782),
            .lcout(\transmit_module.TX_ADDR_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24092),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_14_i1_3_lut_LC_15_15_2 .C_ON=1'b0;
    defparam \transmit_module.mux_14_i1_3_lut_LC_15_15_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_14_i1_3_lut_LC_15_15_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \transmit_module.mux_14_i1_3_lut_LC_15_15_2  (
            .in0(N__14002),
            .in1(N__14274),
            .in2(_gnd_net_),
            .in3(N__13908),
            .lcout(\transmit_module.n147 ),
            .ltout(\transmit_module.n147_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1637_4_lut_LC_15_15_3 .C_ON=1'b0;
    defparam \transmit_module.i1637_4_lut_LC_15_15_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1637_4_lut_LC_15_15_3 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \transmit_module.i1637_4_lut_LC_15_15_3  (
            .in0(N__23141),
            .in1(N__16233),
            .in2(N__14268),
            .in3(N__13928),
            .lcout(n28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_14_i5_3_lut_LC_15_15_4 .C_ON=1'b0;
    defparam \transmit_module.mux_14_i5_3_lut_LC_15_15_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_14_i5_3_lut_LC_15_15_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_14_i5_3_lut_LC_15_15_4  (
            .in0(N__14000),
            .in1(N__15514),
            .in2(_gnd_net_),
            .in3(N__13962),
            .lcout(\transmit_module.n143 ),
            .ltout(\transmit_module.n143_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i4_LC_15_15_5 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i4_LC_15_15_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i4_LC_15_15_5 .LUT_INIT=16'b0100010001010000;
    LogicCell40 \transmit_module.BRAM_ADDR__i4_LC_15_15_5  (
            .in0(N__23142),
            .in1(N__13944),
            .in2(N__13932),
            .in3(N__16237),
            .lcout(\transmit_module.TX_ADDR_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24092),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i0_LC_15_15_6 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i0_LC_15_15_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i0_LC_15_15_6 .LUT_INIT=16'b0010001100100000;
    LogicCell40 \transmit_module.BRAM_ADDR__i0_LC_15_15_6  (
            .in0(N__13929),
            .in1(N__23144),
            .in2(N__16266),
            .in3(N__13920),
            .lcout(\transmit_module.TX_ADDR_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24092),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_2_lut_LC_15_16_0 .C_ON=1'b1;
    defparam \receive_module.add_12_2_lut_LC_15_16_0 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_2_lut_LC_15_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_2_lut_LC_15_16_0  (
            .in0(_gnd_net_),
            .in1(N__14637),
            .in2(_gnd_net_),
            .in3(N__13884),
            .lcout(\receive_module.n137 ),
            .ltout(),
            .carryin(bfn_15_16_0_),
            .carryout(\receive_module.n3146 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_3_lut_LC_15_16_1 .C_ON=1'b1;
    defparam \receive_module.add_12_3_lut_LC_15_16_1 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_3_lut_LC_15_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_3_lut_LC_15_16_1  (
            .in0(_gnd_net_),
            .in1(N__15123),
            .in2(_gnd_net_),
            .in3(N__13881),
            .lcout(\receive_module.n136 ),
            .ltout(),
            .carryin(\receive_module.n3146 ),
            .carryout(\receive_module.n3147 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_4_lut_LC_15_16_2 .C_ON=1'b1;
    defparam \receive_module.add_12_4_lut_LC_15_16_2 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_4_lut_LC_15_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_4_lut_LC_15_16_2  (
            .in0(_gnd_net_),
            .in1(N__14356),
            .in2(_gnd_net_),
            .in3(N__13878),
            .lcout(\receive_module.n135 ),
            .ltout(),
            .carryin(\receive_module.n3147 ),
            .carryout(\receive_module.n3148 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_5_lut_LC_15_16_3 .C_ON=1'b1;
    defparam \receive_module.add_12_5_lut_LC_15_16_3 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_5_lut_LC_15_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_5_lut_LC_15_16_3  (
            .in0(_gnd_net_),
            .in1(N__17617),
            .in2(_gnd_net_),
            .in3(N__13875),
            .lcout(\receive_module.n134 ),
            .ltout(),
            .carryin(\receive_module.n3148 ),
            .carryout(\receive_module.n3149 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_6_lut_LC_15_16_4 .C_ON=1'b1;
    defparam \receive_module.add_12_6_lut_LC_15_16_4 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_6_lut_LC_15_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_6_lut_LC_15_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17362),
            .in3(N__14301),
            .lcout(\receive_module.n133 ),
            .ltout(),
            .carryin(\receive_module.n3149 ),
            .carryout(\receive_module.n3150 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_7_lut_LC_15_16_5 .C_ON=1'b1;
    defparam \receive_module.add_12_7_lut_LC_15_16_5 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_7_lut_LC_15_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_7_lut_LC_15_16_5  (
            .in0(_gnd_net_),
            .in1(N__19348),
            .in2(_gnd_net_),
            .in3(N__14298),
            .lcout(\receive_module.n132 ),
            .ltout(),
            .carryin(\receive_module.n3150 ),
            .carryout(\receive_module.n3151 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_8_lut_LC_15_16_6 .C_ON=1'b1;
    defparam \receive_module.add_12_8_lut_LC_15_16_6 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_8_lut_LC_15_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_8_lut_LC_15_16_6  (
            .in0(_gnd_net_),
            .in1(N__16864),
            .in2(_gnd_net_),
            .in3(N__14295),
            .lcout(\receive_module.n131 ),
            .ltout(),
            .carryin(\receive_module.n3151 ),
            .carryout(\receive_module.n3152 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_9_lut_LC_15_16_7 .C_ON=1'b1;
    defparam \receive_module.add_12_9_lut_LC_15_16_7 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_9_lut_LC_15_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_9_lut_LC_15_16_7  (
            .in0(_gnd_net_),
            .in1(N__16618),
            .in2(_gnd_net_),
            .in3(N__14292),
            .lcout(\receive_module.n130 ),
            .ltout(),
            .carryin(\receive_module.n3152 ),
            .carryout(\receive_module.n3153 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_10_lut_LC_15_17_0 .C_ON=1'b1;
    defparam \receive_module.add_12_10_lut_LC_15_17_0 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_10_lut_LC_15_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_10_lut_LC_15_17_0  (
            .in0(_gnd_net_),
            .in1(N__17116),
            .in2(_gnd_net_),
            .in3(N__14289),
            .lcout(\receive_module.n129 ),
            .ltout(),
            .carryin(bfn_15_17_0_),
            .carryout(\receive_module.n3154 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_11_lut_LC_15_17_1 .C_ON=1'b1;
    defparam \receive_module.add_12_11_lut_LC_15_17_1 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_11_lut_LC_15_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_11_lut_LC_15_17_1  (
            .in0(_gnd_net_),
            .in1(N__17853),
            .in2(_gnd_net_),
            .in3(N__14286),
            .lcout(\receive_module.n128 ),
            .ltout(),
            .carryin(\receive_module.n3154 ),
            .carryout(\receive_module.n3155 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_12_12_lut_LC_15_17_2 .C_ON=1'b1;
    defparam \receive_module.add_12_12_lut_LC_15_17_2 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_12_12_lut_LC_15_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_12_12_lut_LC_15_17_2  (
            .in0(_gnd_net_),
            .in1(N__14880),
            .in2(_gnd_net_),
            .in3(N__14283),
            .lcout(\receive_module.n127 ),
            .ltout(),
            .carryin(\receive_module.n3155 ),
            .carryout(\receive_module.n3156 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.BRAM_ADDR__i11_LC_15_17_3 .C_ON=1'b1;
    defparam \receive_module.BRAM_ADDR__i11_LC_15_17_3 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i11_LC_15_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.BRAM_ADDR__i11_LC_15_17_3  (
            .in0(_gnd_net_),
            .in1(N__18762),
            .in2(_gnd_net_),
            .in3(N__14280),
            .lcout(RX_ADDR_11),
            .ltout(),
            .carryin(\receive_module.n3156 ),
            .carryout(\receive_module.n3157 ),
            .clk(N__21966),
            .ce(N__16164),
            .sr(N__19272));
    defparam \receive_module.BRAM_ADDR__i12_LC_15_17_4 .C_ON=1'b1;
    defparam \receive_module.BRAM_ADDR__i12_LC_15_17_4 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i12_LC_15_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.BRAM_ADDR__i12_LC_15_17_4  (
            .in0(_gnd_net_),
            .in1(N__18919),
            .in2(_gnd_net_),
            .in3(N__14277),
            .lcout(RX_ADDR_12),
            .ltout(),
            .carryin(\receive_module.n3157 ),
            .carryout(\receive_module.n3158 ),
            .clk(N__21966),
            .ce(N__16164),
            .sr(N__19272));
    defparam \receive_module.BRAM_ADDR__i13_LC_15_17_5 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i13_LC_15_17_5 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i13_LC_15_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.BRAM_ADDR__i13_LC_15_17_5  (
            .in0(_gnd_net_),
            .in1(N__18834),
            .in2(_gnd_net_),
            .in3(N__15528),
            .lcout(RX_ADDR_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21966),
            .ce(N__16164),
            .sr(N__19272));
    defparam \transmit_module.ADDR_Y_COMPONENT__i4_LC_15_18_3 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i4_LC_15_18_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i4_LC_15_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i4_LC_15_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15524),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23977),
            .ce(N__15402),
            .sr(N__23252));
    defparam \transmit_module.ADDR_Y_COMPONENT__i7_LC_15_18_4 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i7_LC_15_18_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i7_LC_15_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i7_LC_15_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15489),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23977),
            .ce(N__15402),
            .sr(N__23252));
    defparam \transmit_module.ADDR_Y_COMPONENT__i6_LC_15_18_5 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i6_LC_15_18_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i6_LC_15_18_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i6_LC_15_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15443),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23977),
            .ce(N__15402),
            .sr(N__23252));
    defparam \receive_module.BRAM_ADDR__i1_LC_15_19_1 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i1_LC_15_19_1 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i1_LC_15_19_1 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \receive_module.BRAM_ADDR__i1_LC_15_19_1  (
            .in0(N__20132),
            .in1(N__15327),
            .in2(N__15124),
            .in3(N__19672),
            .lcout(RX_ADDR_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21971),
            .ce(),
            .sr(N__19291));
    defparam \receive_module.BRAM_ADDR__i10_LC_15_19_2 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i10_LC_15_19_2 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i10_LC_15_19_2 .LUT_INIT=16'b1111101101000000;
    LogicCell40 \receive_module.BRAM_ADDR__i10_LC_15_19_2  (
            .in0(N__19671),
            .in1(N__20131),
            .in2(N__14881),
            .in3(N__15090),
            .lcout(RX_ADDR_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21971),
            .ce(),
            .sr(N__19291));
    defparam \receive_module.BRAM_ADDR__i0_LC_15_19_3 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i0_LC_15_19_3 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i0_LC_15_19_3 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \receive_module.BRAM_ADDR__i0_LC_15_19_3  (
            .in0(N__20130),
            .in1(N__14844),
            .in2(N__14638),
            .in3(N__19670),
            .lcout(RX_ADDR_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21971),
            .ce(),
            .sr(N__19291));
    defparam \transmit_module.VGA_R__i1_LC_15_20_5 .C_ON=1'b0;
    defparam \transmit_module.VGA_R__i1_LC_15_20_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.VGA_R__i1_LC_15_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.VGA_R__i1_LC_15_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20919),
            .lcout(n1818),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23845),
            .ce(),
            .sr(N__22397));
    defparam \receive_module.BRAM_ADDR__i2_LC_15_31_2 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i2_LC_15_31_2 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i2_LC_15_31_2 .LUT_INIT=16'b1100111011000100;
    LogicCell40 \receive_module.BRAM_ADDR__i2_LC_15_31_2  (
            .in0(N__20139),
            .in1(N__14553),
            .in2(N__19697),
            .in3(N__14328),
            .lcout(RX_ADDR_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21987),
            .ce(),
            .sr(N__19302));
    defparam \tvp_video_buffer.BUFFER_0__i12_LC_16_3_5 .C_ON=1'b0;
    defparam \tvp_video_buffer.BUFFER_0__i12_LC_16_3_5 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.BUFFER_0__i12_LC_16_3_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.BUFFER_0__i12_LC_16_3_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15681),
            .lcout(\tvp_video_buffer.BUFFER_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21927),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i2_4_lut_LC_16_9_0 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i2_4_lut_LC_16_9_0 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i2_4_lut_LC_16_9_0 .LUT_INIT=16'b1111111111101100;
    LogicCell40 \receive_module.rx_counter.i2_4_lut_LC_16_9_0  (
            .in0(N__18621),
            .in1(N__18544),
            .in2(N__18600),
            .in3(N__18570),
            .lcout(),
            .ltout(\receive_module.rx_counter.n3452_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i1_4_lut_adj_22_LC_16_9_1 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i1_4_lut_adj_22_LC_16_9_1 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i1_4_lut_adj_22_LC_16_9_1 .LUT_INIT=16'b1100110010000000;
    LogicCell40 \receive_module.rx_counter.i1_4_lut_adj_22_LC_16_9_1  (
            .in0(N__18521),
            .in1(N__18461),
            .in2(N__15672),
            .in3(N__15761),
            .lcout(\receive_module.rx_counter.n4_adj_612 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i2_2_lut_LC_16_9_3 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i2_2_lut_LC_16_9_3 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i2_2_lut_LC_16_9_3 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \receive_module.rx_counter.i2_2_lut_LC_16_9_3  (
            .in0(N__18520),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18460),
            .lcout(\receive_module.rx_counter.n10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.WIRE_OUT_i3_LC_16_9_5 .C_ON=1'b0;
    defparam \tvp_video_buffer.WIRE_OUT_i3_LC_16_9_5 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.WIRE_OUT_i3_LC_16_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.WIRE_OUT_i3_LC_16_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15669),
            .lcout(RX_DATA_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21937),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i1_2_lut_adj_27_LC_16_9_6 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i1_2_lut_adj_27_LC_16_9_6 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i1_2_lut_adj_27_LC_16_9_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \receive_module.rx_counter.i1_2_lut_adj_27_LC_16_9_6  (
            .in0(_gnd_net_),
            .in1(N__18519),
            .in2(_gnd_net_),
            .in3(N__18543),
            .lcout(\receive_module.rx_counter.n4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i2_3_lut_LC_16_10_0 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i2_3_lut_LC_16_10_0 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i2_3_lut_LC_16_10_0 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \receive_module.rx_counter.i2_3_lut_LC_16_10_0  (
            .in0(N__18594),
            .in1(N__18622),
            .in2(_gnd_net_),
            .in3(N__18571),
            .lcout(\receive_module.rx_counter.n3450 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i6_4_lut_LC_16_10_1 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i6_4_lut_LC_16_10_1 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i6_4_lut_LC_16_10_1 .LUT_INIT=16'b1111111111011111;
    LogicCell40 \receive_module.rx_counter.i6_4_lut_LC_16_10_1  (
            .in0(N__18572),
            .in1(N__18595),
            .in2(N__18549),
            .in3(N__19179),
            .lcout(),
            .ltout(\receive_module.rx_counter.n14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.SYNC_46_LC_16_10_2 .C_ON=1'b0;
    defparam \receive_module.rx_counter.SYNC_46_LC_16_10_2 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.SYNC_46_LC_16_10_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \receive_module.rx_counter.SYNC_46_LC_16_10_2  (
            .in0(N__15552),
            .in1(N__18623),
            .in2(N__15543),
            .in3(N__15762),
            .lcout(RX_TX_SYNC),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21942),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i1_2_lut_3_lut_LC_16_10_3 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i1_2_lut_3_lut_LC_16_10_3 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i1_2_lut_3_lut_LC_16_10_3 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \receive_module.rx_counter.i1_2_lut_3_lut_LC_16_10_3  (
            .in0(N__18500),
            .in1(N__18459),
            .in2(_gnd_net_),
            .in3(N__18482),
            .lcout(),
            .ltout(\receive_module.rx_counter.n5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i3_4_lut_adj_21_LC_16_10_4 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i3_4_lut_adj_21_LC_16_10_4 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i3_4_lut_adj_21_LC_16_10_4 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \receive_module.rx_counter.i3_4_lut_adj_21_LC_16_10_4  (
            .in0(N__19180),
            .in1(N__15780),
            .in2(N__15771),
            .in3(N__15768),
            .lcout(\receive_module.rx_counter.n3478 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i606_2_lut_rep_21_LC_16_10_6 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i606_2_lut_rep_21_LC_16_10_6 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i606_2_lut_rep_21_LC_16_10_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \receive_module.rx_counter.i606_2_lut_rep_21_LC_16_10_6  (
            .in0(_gnd_net_),
            .in1(N__18481),
            .in2(_gnd_net_),
            .in3(N__18499),
            .lcout(\receive_module.rx_counter.n3677 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i5_1_lut_LC_16_10_7 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i5_1_lut_LC_16_10_7 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i5_1_lut_LC_16_10_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \receive_module.rx_counter.i5_1_lut_LC_16_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20001),
            .lcout(\receive_module.rx_counter.n3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i2_3_lut_adj_23_LC_16_11_5 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i2_3_lut_adj_23_LC_16_11_5 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i2_3_lut_adj_23_LC_16_11_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \receive_module.rx_counter.i2_3_lut_adj_23_LC_16_11_5  (
            .in0(N__15728),
            .in1(N__15716),
            .in2(_gnd_net_),
            .in3(N__15704),
            .lcout(\receive_module.rx_counter.n3222 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.FRAME_COUNTER_244__i0_LC_16_12_0 .C_ON=1'b1;
    defparam \receive_module.rx_counter.FRAME_COUNTER_244__i0_LC_16_12_0 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.FRAME_COUNTER_244__i0_LC_16_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.FRAME_COUNTER_244__i0_LC_16_12_0  (
            .in0(_gnd_net_),
            .in1(N__19032),
            .in2(_gnd_net_),
            .in3(N__15693),
            .lcout(\receive_module.rx_counter.FRAME_COUNTER_0 ),
            .ltout(),
            .carryin(bfn_16_12_0_),
            .carryout(\receive_module.rx_counter.n3202 ),
            .clk(N__21953),
            .ce(N__18947),
            .sr(N__18981));
    defparam \receive_module.rx_counter.FRAME_COUNTER_244__i1_LC_16_12_1 .C_ON=1'b1;
    defparam \receive_module.rx_counter.FRAME_COUNTER_244__i1_LC_16_12_1 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.FRAME_COUNTER_244__i1_LC_16_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.FRAME_COUNTER_244__i1_LC_16_12_1  (
            .in0(_gnd_net_),
            .in1(N__16020),
            .in2(_gnd_net_),
            .in3(N__15690),
            .lcout(\receive_module.rx_counter.FRAME_COUNTER_1 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3202 ),
            .carryout(\receive_module.rx_counter.n3203 ),
            .clk(N__21953),
            .ce(N__18947),
            .sr(N__18981));
    defparam \receive_module.rx_counter.FRAME_COUNTER_244__i2_LC_16_12_2 .C_ON=1'b1;
    defparam \receive_module.rx_counter.FRAME_COUNTER_244__i2_LC_16_12_2 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.FRAME_COUNTER_244__i2_LC_16_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.FRAME_COUNTER_244__i2_LC_16_12_2  (
            .in0(_gnd_net_),
            .in1(N__19044),
            .in2(_gnd_net_),
            .in3(N__15687),
            .lcout(\receive_module.rx_counter.FRAME_COUNTER_2 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3203 ),
            .carryout(\receive_module.rx_counter.n3204 ),
            .clk(N__21953),
            .ce(N__18947),
            .sr(N__18981));
    defparam \receive_module.rx_counter.FRAME_COUNTER_244__i3_LC_16_12_3 .C_ON=1'b1;
    defparam \receive_module.rx_counter.FRAME_COUNTER_244__i3_LC_16_12_3 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.FRAME_COUNTER_244__i3_LC_16_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.FRAME_COUNTER_244__i3_LC_16_12_3  (
            .in0(_gnd_net_),
            .in1(N__19020),
            .in2(_gnd_net_),
            .in3(N__15684),
            .lcout(\receive_module.rx_counter.FRAME_COUNTER_3 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3204 ),
            .carryout(\receive_module.rx_counter.n3205 ),
            .clk(N__21953),
            .ce(N__18947),
            .sr(N__18981));
    defparam \receive_module.rx_counter.FRAME_COUNTER_244__i4_LC_16_12_4 .C_ON=1'b1;
    defparam \receive_module.rx_counter.FRAME_COUNTER_244__i4_LC_16_12_4 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.FRAME_COUNTER_244__i4_LC_16_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.FRAME_COUNTER_244__i4_LC_16_12_4  (
            .in0(_gnd_net_),
            .in1(N__19056),
            .in2(_gnd_net_),
            .in3(N__16050),
            .lcout(\receive_module.rx_counter.FRAME_COUNTER_4 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3205 ),
            .carryout(\receive_module.rx_counter.n3206 ),
            .clk(N__21953),
            .ce(N__18947),
            .sr(N__18981));
    defparam \receive_module.rx_counter.FRAME_COUNTER_244__i5_LC_16_12_5 .C_ON=1'b0;
    defparam \receive_module.rx_counter.FRAME_COUNTER_244__i5_LC_16_12_5 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.FRAME_COUNTER_244__i5_LC_16_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.FRAME_COUNTER_244__i5_LC_16_12_5  (
            .in0(_gnd_net_),
            .in1(N__16032),
            .in2(_gnd_net_),
            .in3(N__16047),
            .lcout(\receive_module.rx_counter.FRAME_COUNTER_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21953),
            .ce(N__18947),
            .sr(N__18981));
    defparam \receive_module.rx_counter.i2089_4_lut_LC_16_13_3 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i2089_4_lut_LC_16_13_3 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i2089_4_lut_LC_16_13_3 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \receive_module.rx_counter.i2089_4_lut_LC_16_13_3  (
            .in0(N__16044),
            .in1(N__16038),
            .in2(N__15909),
            .in3(N__15924),
            .lcout(\receive_module.rx_counter.n3426 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i2182_2_lut_LC_16_13_5 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i2182_2_lut_LC_16_13_5 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i2182_2_lut_LC_16_13_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \receive_module.rx_counter.i2182_2_lut_LC_16_13_5  (
            .in0(_gnd_net_),
            .in1(N__16031),
            .in2(_gnd_net_),
            .in3(N__16019),
            .lcout(\receive_module.rx_counter.n3519 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i3_4_lut_LC_16_14_2 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i3_4_lut_LC_16_14_2 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i3_4_lut_LC_16_14_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \receive_module.rx_counter.i3_4_lut_LC_16_14_2  (
            .in0(N__16008),
            .in1(N__15981),
            .in2(N__15954),
            .in3(N__15923),
            .lcout(),
            .ltout(\receive_module.rx_counter.n3455_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i1_4_lut_LC_16_14_3 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i1_4_lut_LC_16_14_3 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i1_4_lut_LC_16_14_3 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \receive_module.rx_counter.i1_4_lut_LC_16_14_3  (
            .in0(N__15908),
            .in1(N__15848),
            .in2(N__15879),
            .in3(N__15876),
            .lcout(),
            .ltout(\receive_module.rx_counter.n39_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i58_4_lut_LC_16_14_4 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i58_4_lut_LC_16_14_4 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i58_4_lut_LC_16_14_4 .LUT_INIT=16'b1100000011010001;
    LogicCell40 \receive_module.rx_counter.i58_4_lut_LC_16_14_4  (
            .in0(N__15849),
            .in1(N__15828),
            .in2(N__15810),
            .in3(N__15807),
            .lcout(),
            .ltout(\receive_module.rx_counter.n54_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.O_VISIBLE_53_LC_16_14_5 .C_ON=1'b0;
    defparam \receive_module.rx_counter.O_VISIBLE_53_LC_16_14_5 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.O_VISIBLE_53_LC_16_14_5 .LUT_INIT=16'b0000010000001100;
    LogicCell40 \receive_module.rx_counter.O_VISIBLE_53_LC_16_14_5  (
            .in0(N__19191),
            .in1(N__15801),
            .in2(N__15792),
            .in3(N__15789),
            .lcout(DEBUG_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21960),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_17_LC_16_15_3 .C_ON=1'b0;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_17_LC_16_15_3 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_17_LC_16_15_3 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \line_buffer.i1_2_lut_3_lut_4_lut_adj_17_LC_16_15_3  (
            .in0(N__18920),
            .in1(N__19592),
            .in2(N__18866),
            .in3(N__18779),
            .lcout(\line_buffer.n473 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_19_LC_16_15_5 .C_ON=1'b0;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_19_LC_16_15_5 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_19_LC_16_15_5 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \line_buffer.i1_2_lut_3_lut_4_lut_adj_19_LC_16_15_5  (
            .in0(N__18921),
            .in1(N__19591),
            .in2(N__18867),
            .in3(N__18780),
            .lcout(\line_buffer.n570 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_20_LC_16_15_6 .C_ON=1'b0;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_20_LC_16_15_6 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_20_LC_16_15_6 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \line_buffer.i1_2_lut_3_lut_4_lut_adj_20_LC_16_15_6  (
            .in0(N__18781),
            .in1(N__18922),
            .in2(N__18871),
            .in3(N__19593),
            .lcout(\line_buffer.n571 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__rep_1_i0_LC_16_16_1 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__rep_1_i0_LC_16_16_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__rep_1_i0_LC_16_16_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \transmit_module.BRAM_ADDR__rep_1_i0_LC_16_16_1  (
            .in0(N__16377),
            .in1(N__16320),
            .in2(_gnd_net_),
            .in3(N__16365),
            .lcout(TX_ADDR_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24102),
            .ce(N__16179),
            .sr(N__23243));
    defparam \transmit_module.BRAM_ADDR__i13_LC_16_16_4 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i13_LC_16_16_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i13_LC_16_16_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \transmit_module.BRAM_ADDR__i13_LC_16_16_4  (
            .in0(N__16319),
            .in1(N__16356),
            .in2(_gnd_net_),
            .in3(N__16344),
            .lcout(TX_ADDR_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24102),
            .ce(N__16179),
            .sr(N__23243));
    defparam \transmit_module.BRAM_ADDR__i12_LC_16_16_5 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i12_LC_16_16_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i12_LC_16_16_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \transmit_module.BRAM_ADDR__i12_LC_16_16_5  (
            .in0(N__16335),
            .in1(N__16318),
            .in2(_gnd_net_),
            .in3(N__16188),
            .lcout(TX_ADDR_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24102),
            .ce(N__16179),
            .sr(N__23243));
    defparam \receive_module.rx_counter.i246_2_lut_rep_15_2_lut_LC_16_17_0 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i246_2_lut_rep_15_2_lut_LC_16_17_0 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i246_2_lut_rep_15_2_lut_LC_16_17_0 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \receive_module.rx_counter.i246_2_lut_rep_15_2_lut_LC_16_17_0  (
            .in0(_gnd_net_),
            .in1(N__19645),
            .in2(_gnd_net_),
            .in3(N__20104),
            .lcout(\receive_module.n3671 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_16_LC_16_17_1 .C_ON=1'b0;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_16_LC_16_17_1 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_16_LC_16_17_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \line_buffer.i1_2_lut_3_lut_4_lut_adj_16_LC_16_17_1  (
            .in0(N__18777),
            .in1(N__18833),
            .in2(N__19676),
            .in3(N__18918),
            .lcout(\line_buffer.n603 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_LC_16_17_4 .C_ON=1'b0;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_LC_16_17_4 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_LC_16_17_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \line_buffer.i1_2_lut_3_lut_4_lut_LC_16_17_4  (
            .in0(N__18917),
            .in1(N__19641),
            .in2(N__18850),
            .in3(N__18776),
            .lcout(\line_buffer.n539 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_18_LC_16_18_7 .C_ON=1'b0;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_18_LC_16_18_7 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_18_LC_16_18_7 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \line_buffer.i1_2_lut_3_lut_4_lut_adj_18_LC_16_18_7  (
            .in0(N__18916),
            .in1(N__19649),
            .in2(N__18849),
            .in3(N__18778),
            .lcout(\line_buffer.n474 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.BRAM_ADDR__i9_LC_16_19_0 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i9_LC_16_19_0 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i9_LC_16_19_0 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \receive_module.BRAM_ADDR__i9_LC_16_19_0  (
            .in0(N__20135),
            .in1(N__19667),
            .in2(N__17854),
            .in3(N__18069),
            .lcout(RX_ADDR_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21968),
            .ce(),
            .sr(N__19300));
    defparam \receive_module.BRAM_ADDR__i3_LC_16_19_3 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i3_LC_16_19_3 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i3_LC_16_19_3 .LUT_INIT=16'b1010111010100010;
    LogicCell40 \receive_module.BRAM_ADDR__i3_LC_16_19_3  (
            .in0(N__17817),
            .in1(N__20133),
            .in2(N__19684),
            .in3(N__17598),
            .lcout(RX_ADDR_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21968),
            .ce(),
            .sr(N__19300));
    defparam \receive_module.BRAM_ADDR__i4_LC_16_19_4 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i4_LC_16_19_4 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i4_LC_16_19_4 .LUT_INIT=16'b1010101011100010;
    LogicCell40 \receive_module.BRAM_ADDR__i4_LC_16_19_4  (
            .in0(N__17571),
            .in1(N__20136),
            .in2(N__17361),
            .in3(N__19659),
            .lcout(RX_ADDR_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21968),
            .ce(),
            .sr(N__19300));
    defparam \receive_module.BRAM_ADDR__i8_LC_16_19_5 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i8_LC_16_19_5 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i8_LC_16_19_5 .LUT_INIT=16'b1111110100001000;
    LogicCell40 \receive_module.BRAM_ADDR__i8_LC_16_19_5  (
            .in0(N__20138),
            .in1(N__17100),
            .in2(N__19686),
            .in3(N__17319),
            .lcout(RX_ADDR_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21968),
            .ce(),
            .sr(N__19300));
    defparam \receive_module.BRAM_ADDR__i6_LC_16_19_6 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i6_LC_16_19_6 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i6_LC_16_19_6 .LUT_INIT=16'b1111110100100000;
    LogicCell40 \receive_module.BRAM_ADDR__i6_LC_16_19_6  (
            .in0(N__20134),
            .in1(N__19660),
            .in2(N__16857),
            .in3(N__17073),
            .lcout(RX_ADDR_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21968),
            .ce(),
            .sr(N__19300));
    defparam \receive_module.BRAM_ADDR__i7_LC_16_19_7 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i7_LC_16_19_7 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i7_LC_16_19_7 .LUT_INIT=16'b1111110100001000;
    LogicCell40 \receive_module.BRAM_ADDR__i7_LC_16_19_7  (
            .in0(N__20137),
            .in1(N__16599),
            .in2(N__19685),
            .in3(N__16818),
            .lcout(RX_ADDR_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21968),
            .ce(),
            .sr(N__19300));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2257_LC_16_20_3 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2257_LC_16_20_3 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2257_LC_16_20_3 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_2257_LC_16_20_3  (
            .in0(N__22754),
            .in1(N__16572),
            .in2(N__21497),
            .in3(N__16551),
            .lcout(\line_buffer.n3587 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n3623_bdd_4_lut_LC_16_20_7 .C_ON=1'b0;
    defparam \line_buffer.n3623_bdd_4_lut_LC_16_20_7 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3623_bdd_4_lut_LC_16_20_7 .LUT_INIT=16'b1110111001010000;
    LogicCell40 \line_buffer.n3623_bdd_4_lut_LC_16_20_7  (
            .in0(N__21458),
            .in1(N__18438),
            .in2(N__18414),
            .in3(N__19200),
            .lcout(\line_buffer.n3626 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n3587_bdd_4_lut_LC_16_21_5 .C_ON=1'b0;
    defparam \line_buffer.n3587_bdd_4_lut_LC_16_21_5 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3587_bdd_4_lut_LC_16_21_5 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \line_buffer.n3587_bdd_4_lut_LC_16_21_5  (
            .in0(N__18393),
            .in1(N__21459),
            .in2(N__18381),
            .in3(N__18360),
            .lcout(),
            .ltout(\line_buffer.n3590_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i3_LC_16_21_6 .C_ON=1'b0;
    defparam \line_buffer.dout_i3_LC_16_21_6 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i3_LC_16_21_6 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \line_buffer.dout_i3_LC_16_21_6  (
            .in0(_gnd_net_),
            .in1(N__21293),
            .in2(N__18354),
            .in3(N__18351),
            .lcout(TX_DATA_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23771),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.VGA_R__i4_LC_16_22_7 .C_ON=1'b0;
    defparam \transmit_module.VGA_R__i4_LC_16_22_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.VGA_R__i4_LC_16_22_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.VGA_R__i4_LC_16_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18345),
            .lcout(n1815),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23653),
            .ce(),
            .sr(N__22426));
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_15_LC_16_23_6 .C_ON=1'b0;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_15_LC_16_23_6 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_15_LC_16_23_6 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \line_buffer.i1_2_lut_3_lut_4_lut_adj_15_LC_16_23_6  (
            .in0(N__18930),
            .in1(N__19680),
            .in2(N__18872),
            .in3(N__18789),
            .lcout(\line_buffer.n602 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam GB_BUFFER_DEBUG_c_3_c_THRU_LUT4_0_LC_16_26_4.C_ON=1'b0;
    defparam GB_BUFFER_DEBUG_c_3_c_THRU_LUT4_0_LC_16_26_4.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_DEBUG_c_3_c_THRU_LUT4_0_LC_16_26_4.LUT_INIT=16'b1010101010101010;
    LogicCell40 GB_BUFFER_DEBUG_c_3_c_THRU_LUT4_0_LC_16_26_4 (
            .in0(N__21999),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(GB_BUFFER_DEBUG_c_3_c_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam PULSE_1HZ_I_0_2_lut_LC_17_5_5.C_ON=1'b0;
    defparam PULSE_1HZ_I_0_2_lut_LC_17_5_5.SEQ_MODE=4'b0000;
    defparam PULSE_1HZ_I_0_2_lut_LC_17_5_5.LUT_INIT=16'b1111111111001100;
    LogicCell40 PULSE_1HZ_I_0_2_lut_LC_17_5_5 (
            .in0(_gnd_net_),
            .in1(N__18176),
            .in2(_gnd_net_),
            .in3(N__18966),
            .lcout(LED_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.BUFFER_0__i1_LC_17_8_4 .C_ON=1'b0;
    defparam \tvp_video_buffer.BUFFER_0__i1_LC_17_8_4 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.BUFFER_0__i1_LC_17_8_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \tvp_video_buffer.BUFFER_0__i1_LC_17_8_4  (
            .in0(N__18132),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\tvp_video_buffer.BUFFER_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21928),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.BUFFER_0__i9_LC_17_8_5 .C_ON=1'b0;
    defparam \tvp_video_buffer.BUFFER_0__i9_LC_17_8_5 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.BUFFER_0__i9_LC_17_8_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.BUFFER_0__i9_LC_17_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18114),
            .lcout(\tvp_video_buffer.BUFFER_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21928),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.Y__i0_LC_17_9_0 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i0_LC_17_9_0 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i0_LC_17_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i0_LC_17_9_0  (
            .in0(_gnd_net_),
            .in1(N__18624),
            .in2(_gnd_net_),
            .in3(N__18603),
            .lcout(\receive_module.rx_counter.Y_0 ),
            .ltout(),
            .carryin(bfn_17_9_0_),
            .carryout(\receive_module.rx_counter.n3172 ),
            .clk(N__21930),
            .ce(N__20022),
            .sr(N__19299));
    defparam \receive_module.rx_counter.Y__i1_LC_17_9_1 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i1_LC_17_9_1 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i1_LC_17_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i1_LC_17_9_1  (
            .in0(_gnd_net_),
            .in1(N__18599),
            .in2(_gnd_net_),
            .in3(N__18576),
            .lcout(\receive_module.rx_counter.Y_1 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3172 ),
            .carryout(\receive_module.rx_counter.n3173 ),
            .clk(N__21930),
            .ce(N__20022),
            .sr(N__19299));
    defparam \receive_module.rx_counter.Y__i2_LC_17_9_2 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i2_LC_17_9_2 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i2_LC_17_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i2_LC_17_9_2  (
            .in0(_gnd_net_),
            .in1(N__18573),
            .in2(_gnd_net_),
            .in3(N__18552),
            .lcout(\receive_module.rx_counter.Y_2 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3173 ),
            .carryout(\receive_module.rx_counter.n3174 ),
            .clk(N__21930),
            .ce(N__20022),
            .sr(N__19299));
    defparam \receive_module.rx_counter.Y__i3_LC_17_9_3 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i3_LC_17_9_3 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i3_LC_17_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i3_LC_17_9_3  (
            .in0(_gnd_net_),
            .in1(N__18545),
            .in2(_gnd_net_),
            .in3(N__18525),
            .lcout(\receive_module.rx_counter.Y_3 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3174 ),
            .carryout(\receive_module.rx_counter.n3175 ),
            .clk(N__21930),
            .ce(N__20022),
            .sr(N__19299));
    defparam \receive_module.rx_counter.Y__i4_LC_17_9_4 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i4_LC_17_9_4 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i4_LC_17_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i4_LC_17_9_4  (
            .in0(_gnd_net_),
            .in1(N__18522),
            .in2(_gnd_net_),
            .in3(N__18504),
            .lcout(\receive_module.rx_counter.Y_4 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3175 ),
            .carryout(\receive_module.rx_counter.n3176 ),
            .clk(N__21930),
            .ce(N__20022),
            .sr(N__19299));
    defparam \receive_module.rx_counter.Y__i5_LC_17_9_5 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i5_LC_17_9_5 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i5_LC_17_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i5_LC_17_9_5  (
            .in0(_gnd_net_),
            .in1(N__18501),
            .in2(_gnd_net_),
            .in3(N__18486),
            .lcout(\receive_module.rx_counter.Y_5 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3176 ),
            .carryout(\receive_module.rx_counter.n3177 ),
            .clk(N__21930),
            .ce(N__20022),
            .sr(N__19299));
    defparam \receive_module.rx_counter.Y__i6_LC_17_9_6 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i6_LC_17_9_6 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i6_LC_17_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i6_LC_17_9_6  (
            .in0(_gnd_net_),
            .in1(N__18483),
            .in2(_gnd_net_),
            .in3(N__18465),
            .lcout(\receive_module.rx_counter.Y_6 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3177 ),
            .carryout(\receive_module.rx_counter.n3178 ),
            .clk(N__21930),
            .ce(N__20022),
            .sr(N__19299));
    defparam \receive_module.rx_counter.Y__i7_LC_17_9_7 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i7_LC_17_9_7 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i7_LC_17_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i7_LC_17_9_7  (
            .in0(_gnd_net_),
            .in1(N__18462),
            .in2(_gnd_net_),
            .in3(N__18441),
            .lcout(\receive_module.rx_counter.Y_7 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3178 ),
            .carryout(\receive_module.rx_counter.n3179 ),
            .clk(N__21930),
            .ce(N__20022),
            .sr(N__19299));
    defparam \receive_module.rx_counter.Y__i8_LC_17_10_0 .C_ON=1'b0;
    defparam \receive_module.rx_counter.Y__i8_LC_17_10_0 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i8_LC_17_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i8_LC_17_10_0  (
            .in0(_gnd_net_),
            .in1(N__19190),
            .in2(_gnd_net_),
            .in3(N__19194),
            .lcout(\receive_module.rx_counter.Y_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21935),
            .ce(N__20018),
            .sr(N__19298));
    defparam \tvp_video_buffer.WIRE_OUT_i0_LC_17_11_4 .C_ON=1'b0;
    defparam \tvp_video_buffer.WIRE_OUT_i0_LC_17_11_4 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.WIRE_OUT_i0_LC_17_11_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.WIRE_OUT_i0_LC_17_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19164),
            .lcout(RX_DATA_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21940),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i1_2_lut_adj_26_LC_17_12_1 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i1_2_lut_adj_26_LC_17_12_1 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i1_2_lut_adj_26_LC_17_12_1 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \receive_module.rx_counter.i1_2_lut_adj_26_LC_17_12_1  (
            .in0(_gnd_net_),
            .in1(N__19055),
            .in2(_gnd_net_),
            .in3(N__19043),
            .lcout(),
            .ltout(\receive_module.rx_counter.n7_adj_619_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i5_4_lut_LC_17_12_2 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i5_4_lut_LC_17_12_2 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i5_4_lut_LC_17_12_2 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \receive_module.rx_counter.i5_4_lut_LC_17_12_2  (
            .in0(N__19031),
            .in1(N__19019),
            .in2(N__19008),
            .in3(N__19005),
            .lcout(\receive_module.rx_counter.n11 ),
            .ltout(\receive_module.rx_counter.n11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i1304_2_lut_3_lut_3_lut_LC_17_12_3 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i1304_2_lut_3_lut_3_lut_LC_17_12_3 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i1304_2_lut_3_lut_3_lut_LC_17_12_3 .LUT_INIT=16'b0000000000001010;
    LogicCell40 \receive_module.rx_counter.i1304_2_lut_3_lut_3_lut_LC_17_12_3  (
            .in0(N__18999),
            .in1(_gnd_net_),
            .in2(N__18984),
            .in3(N__20079),
            .lcout(\receive_module.rx_counter.n2547 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.PULSE_1HZ_49_LC_17_12_7 .C_ON=1'b0;
    defparam \receive_module.rx_counter.PULSE_1HZ_49_LC_17_12_7 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.PULSE_1HZ_49_LC_17_12_7 .LUT_INIT=16'b1001100110011001;
    LogicCell40 \receive_module.rx_counter.PULSE_1HZ_49_LC_17_12_7  (
            .in0(N__18972),
            .in1(N__18959),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(PULSE_1HZ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21946),
            .ce(N__18948),
            .sr(_gnd_net_));
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_14_LC_17_13_0 .C_ON=1'b0;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_14_LC_17_13_0 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_14_LC_17_13_0 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \line_buffer.i1_2_lut_3_lut_4_lut_adj_14_LC_17_13_0  (
            .in0(N__18929),
            .in1(N__19594),
            .in2(N__18873),
            .in3(N__18788),
            .lcout(\line_buffer.n538 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.X_DELTA_PATTERN_i15_LC_17_14_7 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i15_LC_17_14_7 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i15_LC_17_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i15_LC_17_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18690),
            .lcout(\transmit_module.X_DELTA_PATTERN_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24251),
            .ce(N__18662),
            .sr(N__20515));
    defparam \tvp_video_buffer.BUFFER_0__i7_LC_17_15_0 .C_ON=1'b0;
    defparam \tvp_video_buffer.BUFFER_0__i7_LC_17_15_0 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.BUFFER_0__i7_LC_17_15_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \tvp_video_buffer.BUFFER_0__i7_LC_17_15_0  (
            .in0(N__19955),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\tvp_video_buffer.BUFFER_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21957),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.WIRE_OUT_i6_LC_17_15_4 .C_ON=1'b0;
    defparam \tvp_video_buffer.WIRE_OUT_i6_LC_17_15_4 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.WIRE_OUT_i6_LC_17_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.WIRE_OUT_i6_LC_17_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19812),
            .lcout(RX_DATA_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21957),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.BUFFER_0__i15_LC_17_15_6 .C_ON=1'b0;
    defparam \tvp_video_buffer.BUFFER_0__i15_LC_17_15_6 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.BUFFER_0__i15_LC_17_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.BUFFER_0__i15_LC_17_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19818),
            .lcout(\tvp_video_buffer.BUFFER_1_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21957),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2281_LC_17_16_2 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2281_LC_17_16_2 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2281_LC_17_16_2 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_2281_LC_17_16_2  (
            .in0(N__22707),
            .in1(N__19806),
            .in2(N__21464),
            .in3(N__19791),
            .lcout(),
            .ltout(\line_buffer.n3593_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n3593_bdd_4_lut_LC_17_16_3 .C_ON=1'b0;
    defparam \line_buffer.n3593_bdd_4_lut_LC_17_16_3 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3593_bdd_4_lut_LC_17_16_3 .LUT_INIT=16'b1111000011001010;
    LogicCell40 \line_buffer.n3593_bdd_4_lut_LC_17_16_3  (
            .in0(N__19779),
            .in1(N__19764),
            .in2(N__19743),
            .in3(N__21414),
            .lcout(\line_buffer.n3596 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2291_LC_17_17_3 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2291_LC_17_17_3 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2291_LC_17_17_3 .LUT_INIT=16'b1110101001001010;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_2291_LC_17_17_3  (
            .in0(N__22633),
            .in1(N__19740),
            .in2(N__21463),
            .in3(N__19731),
            .lcout(\line_buffer.n3629 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.BRAM_ADDR__i5_LC_17_19_3 .C_ON=1'b0;
    defparam \receive_module.BRAM_ADDR__i5_LC_17_19_3 .SEQ_MODE=4'b1000;
    defparam \receive_module.BRAM_ADDR__i5_LC_17_19_3 .LUT_INIT=16'b1100111011000100;
    LogicCell40 \receive_module.BRAM_ADDR__i5_LC_17_19_3  (
            .in0(N__20129),
            .in1(N__19713),
            .in2(N__19690),
            .in3(N__19329),
            .lcout(RX_ADDR_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21965),
            .ce(),
            .sr(N__19301));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2286_LC_17_20_6 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2286_LC_17_20_6 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2286_LC_17_20_6 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_2286_LC_17_20_6  (
            .in0(N__22753),
            .in1(N__19227),
            .in2(N__21499),
            .in3(N__19212),
            .lcout(\line_buffer.n3623 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_hs_buffer.BUFFER_0__i2_LC_18_9_0 .C_ON=1'b0;
    defparam \tvp_hs_buffer.BUFFER_0__i2_LC_18_9_0 .SEQ_MODE=4'b1000;
    defparam \tvp_hs_buffer.BUFFER_0__i2_LC_18_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_hs_buffer.BUFFER_0__i2_LC_18_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20151),
            .lcout(\tvp_hs_buffer.BUFFER_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21938),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_hs_buffer.BUFFER_0__i1_LC_18_9_5 .C_ON=1'b0;
    defparam \tvp_hs_buffer.BUFFER_0__i1_LC_18_9_5 .SEQ_MODE=4'b1000;
    defparam \tvp_hs_buffer.BUFFER_0__i1_LC_18_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_hs_buffer.BUFFER_0__i1_LC_18_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20168),
            .lcout(\tvp_hs_buffer.BUFFER_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21938),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_hs_buffer.WIRE_OUT_0__9_LC_18_10_5 .C_ON=1'b0;
    defparam \tvp_hs_buffer.WIRE_OUT_0__9_LC_18_10_5 .SEQ_MODE=4'b1000;
    defparam \tvp_hs_buffer.WIRE_OUT_0__9_LC_18_10_5 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \tvp_hs_buffer.WIRE_OUT_0__9_LC_18_10_5  (
            .in0(_gnd_net_),
            .in1(N__20145),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(TVP_HSYNC_buff),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21943),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i249_3_lut_LC_18_10_6 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i249_3_lut_LC_18_10_6 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i249_3_lut_LC_18_10_6 .LUT_INIT=16'b0010001011111111;
    LogicCell40 \receive_module.rx_counter.i249_3_lut_LC_18_10_6  (
            .in0(N__19983),
            .in1(N__19999),
            .in2(_gnd_net_),
            .in3(N__20100),
            .lcout(\receive_module.rx_counter.n2078 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.old_HS_51_LC_18_10_7 .C_ON=1'b0;
    defparam \receive_module.rx_counter.old_HS_51_LC_18_10_7 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.old_HS_51_LC_18_10_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \receive_module.rx_counter.old_HS_51_LC_18_10_7  (
            .in0(N__20000),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\receive_module.rx_counter.old_HS ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21943),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.Y_DELTA_PATTERN_i92_LC_18_12_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i92_LC_18_12_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i92_LC_18_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i92_LC_18_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21141),
            .lcout(\transmit_module.Y_DELTA_PATTERN_92 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24314),
            .ce(N__23395),
            .sr(N__23283));
    defparam \transmit_module.Y_DELTA_PATTERN_i97_LC_18_13_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i97_LC_18_13_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i97_LC_18_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i97_LC_18_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19977),
            .lcout(\transmit_module.Y_DELTA_PATTERN_97 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24220),
            .ce(N__23387),
            .sr(N__23285));
    defparam \transmit_module.Y_DELTA_PATTERN_i98_LC_18_13_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i98_LC_18_13_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i98_LC_18_13_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i98_LC_18_13_3  (
            .in0(N__20532),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.Y_DELTA_PATTERN_98 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24220),
            .ce(N__23387),
            .sr(N__23285));
    defparam \transmit_module.Y_DELTA_PATTERN_i89_LC_18_13_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i89_LC_18_13_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i89_LC_18_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i89_LC_18_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20640),
            .lcout(\transmit_module.Y_DELTA_PATTERN_89 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24220),
            .ce(N__23387),
            .sr(N__23285));
    defparam \transmit_module.Y_DELTA_PATTERN_i88_LC_18_13_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i88_LC_18_13_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i88_LC_18_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i88_LC_18_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19971),
            .lcout(\transmit_module.Y_DELTA_PATTERN_88 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24220),
            .ce(N__23387),
            .sr(N__23285));
    defparam \transmit_module.Y_DELTA_PATTERN_i91_LC_18_13_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i91_LC_18_13_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i91_LC_18_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i91_LC_18_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20652),
            .lcout(\transmit_module.Y_DELTA_PATTERN_91 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24220),
            .ce(N__23387),
            .sr(N__23285));
    defparam \transmit_module.Y_DELTA_PATTERN_i90_LC_18_13_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i90_LC_18_13_7 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i90_LC_18_13_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i90_LC_18_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20646),
            .lcout(\transmit_module.Y_DELTA_PATTERN_90 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24220),
            .ce(N__23387),
            .sr(N__23285));
    defparam \transmit_module.Y_DELTA_PATTERN_i99_LC_18_14_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i99_LC_18_14_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i99_LC_18_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i99_LC_18_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20634),
            .lcout(\transmit_module.Y_DELTA_PATTERN_99 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24227),
            .ce(N__20516),
            .sr(N__23282));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_LC_18_15_5 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_LC_18_15_5 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_LC_18_15_5 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_LC_18_15_5  (
            .in0(N__22755),
            .in1(N__20370),
            .in2(N__21505),
            .in3(N__20352),
            .lcout(\line_buffer.n3653 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n3629_bdd_4_lut_LC_18_17_0 .C_ON=1'b0;
    defparam \line_buffer.n3629_bdd_4_lut_LC_18_17_0 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3629_bdd_4_lut_LC_18_17_0 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \line_buffer.n3629_bdd_4_lut_LC_18_17_0  (
            .in0(N__20337),
            .in1(N__21478),
            .in2(N__20319),
            .in3(N__20301),
            .lcout(\line_buffer.n3632 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2296_LC_18_17_3 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2296_LC_18_17_3 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2296_LC_18_17_3 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_2296_LC_18_17_3  (
            .in0(N__22723),
            .in1(N__20295),
            .in2(N__21502),
            .in3(N__20277),
            .lcout(),
            .ltout(\line_buffer.n3635_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n3635_bdd_4_lut_LC_18_17_4 .C_ON=1'b0;
    defparam \line_buffer.n3635_bdd_4_lut_LC_18_17_4 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3635_bdd_4_lut_LC_18_17_4 .LUT_INIT=16'b1111000011001010;
    LogicCell40 \line_buffer.n3635_bdd_4_lut_LC_18_17_4  (
            .in0(N__20262),
            .in1(N__20241),
            .in2(N__20223),
            .in3(N__21479),
            .lcout(\line_buffer.n3638 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n3653_bdd_4_lut_LC_18_17_6 .C_ON=1'b0;
    defparam \line_buffer.n3653_bdd_4_lut_LC_18_17_6 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3653_bdd_4_lut_LC_18_17_6 .LUT_INIT=16'b1111101000001100;
    LogicCell40 \line_buffer.n3653_bdd_4_lut_LC_18_17_6  (
            .in0(N__20220),
            .in1(N__20205),
            .in2(N__21503),
            .in3(N__20190),
            .lcout(),
            .ltout(\line_buffer.n3656_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i5_LC_18_17_7 .C_ON=1'b0;
    defparam \line_buffer.dout_i5_LC_18_17_7 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i5_LC_18_17_7 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \line_buffer.dout_i5_LC_18_17_7  (
            .in0(_gnd_net_),
            .in1(N__21267),
            .in2(N__20934),
            .in3(N__20931),
            .lcout(TX_DATA_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24074),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i0_LC_18_18_2 .C_ON=1'b0;
    defparam \line_buffer.dout_i0_LC_18_18_2 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i0_LC_18_18_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \line_buffer.dout_i0_LC_18_18_2  (
            .in0(N__21268),
            .in1(N__20781),
            .in2(_gnd_net_),
            .in3(N__20925),
            .lcout(TX_DATA_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24112),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n3647_bdd_4_lut_LC_18_18_4 .C_ON=1'b0;
    defparam \line_buffer.n3647_bdd_4_lut_LC_18_18_4 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3647_bdd_4_lut_LC_18_18_4 .LUT_INIT=16'b1100110010111000;
    LogicCell40 \line_buffer.n3647_bdd_4_lut_LC_18_18_4  (
            .in0(N__20907),
            .in1(N__20829),
            .in2(N__20886),
            .in3(N__21483),
            .lcout(),
            .ltout(\line_buffer.n3650_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i1_LC_18_18_5 .C_ON=1'b0;
    defparam \line_buffer.dout_i1_LC_18_18_5 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i1_LC_18_18_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \line_buffer.dout_i1_LC_18_18_5  (
            .in0(_gnd_net_),
            .in1(N__20865),
            .in2(N__20859),
            .in3(N__21269),
            .lcout(TX_DATA_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24112),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2306_LC_18_19_1 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2306_LC_18_19_1 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2306_LC_18_19_1 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_2306_LC_18_19_1  (
            .in0(N__22759),
            .in1(N__20856),
            .in2(N__21501),
            .in3(N__20844),
            .lcout(\line_buffer.n3647 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n3641_bdd_4_lut_LC_18_19_3 .C_ON=1'b0;
    defparam \line_buffer.n3641_bdd_4_lut_LC_18_19_3 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n3641_bdd_4_lut_LC_18_19_3 .LUT_INIT=16'b1111101001000100;
    LogicCell40 \line_buffer.n3641_bdd_4_lut_LC_18_19_3  (
            .in0(N__21474),
            .in1(N__20823),
            .in2(N__20805),
            .in3(N__21090),
            .lcout(\line_buffer.n3644 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.VGA_R__i6_LC_18_21_6 .C_ON=1'b0;
    defparam \transmit_module.VGA_R__i6_LC_18_21_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.VGA_R__i6_LC_18_21_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.VGA_R__i6_LC_18_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20775),
            .lcout(n1813),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23772),
            .ce(),
            .sr(N__22425));
    defparam \transmit_module.VGA_R__i2_LC_18_22_7 .C_ON=1'b0;
    defparam \transmit_module.VGA_R__i2_LC_18_22_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.VGA_R__i2_LC_18_22_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.VGA_R__i2_LC_18_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20709),
            .lcout(n1817),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23815),
            .ce(),
            .sr(N__22427));
    defparam \transmit_module.Y_DELTA_PATTERN_i96_LC_19_13_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i96_LC_19_13_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i96_LC_19_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i96_LC_19_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20658),
            .lcout(\transmit_module.Y_DELTA_PATTERN_96 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24213),
            .ce(N__23391),
            .sr(N__23280));
    defparam \transmit_module.Y_DELTA_PATTERN_i94_LC_19_13_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i94_LC_19_13_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i94_LC_19_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i94_LC_19_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21153),
            .lcout(\transmit_module.Y_DELTA_PATTERN_94 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24213),
            .ce(N__23391),
            .sr(N__23280));
    defparam \transmit_module.Y_DELTA_PATTERN_i95_LC_19_13_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i95_LC_19_13_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i95_LC_19_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i95_LC_19_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21159),
            .lcout(\transmit_module.Y_DELTA_PATTERN_95 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24213),
            .ce(N__23391),
            .sr(N__23280));
    defparam \transmit_module.Y_DELTA_PATTERN_i93_LC_19_13_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i93_LC_19_13_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i93_LC_19_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i93_LC_19_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21147),
            .lcout(\transmit_module.Y_DELTA_PATTERN_93 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24213),
            .ce(N__23391),
            .sr(N__23280));
    defparam \transmit_module.Y_DELTA_PATTERN_i83_LC_19_13_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i83_LC_19_13_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i83_LC_19_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i83_LC_19_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21774),
            .lcout(\transmit_module.Y_DELTA_PATTERN_83 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24213),
            .ce(N__23391),
            .sr(N__23280));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2301_LC_19_19_4 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2301_LC_19_19_4 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2301_LC_19_19_4 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_2301_LC_19_19_4  (
            .in0(N__22769),
            .in1(N__21126),
            .in2(N__21504),
            .in3(N__21111),
            .lcout(\line_buffer.n3641 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2196_3_lut_LC_20_7_7 .C_ON=1'b0;
    defparam \line_buffer.i2196_3_lut_LC_20_7_7 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2196_3_lut_LC_20_7_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \line_buffer.i2196_3_lut_LC_20_7_7  (
            .in0(N__22833),
            .in1(N__21084),
            .in2(_gnd_net_),
            .in3(N__21072),
            .lcout(\line_buffer.n3533 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.WIRE_OUT_i7_LC_20_9_0 .C_ON=1'b0;
    defparam \tvp_video_buffer.WIRE_OUT_i7_LC_20_9_0 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.WIRE_OUT_i7_LC_20_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.WIRE_OUT_i7_LC_20_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22005),
            .lcout(RX_DATA_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21948),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2212_3_lut_LC_20_12_6 .C_ON=1'b0;
    defparam \line_buffer.i2212_3_lut_LC_20_12_6 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2212_3_lut_LC_20_12_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \line_buffer.i2212_3_lut_LC_20_12_6  (
            .in0(N__20961),
            .in1(N__20949),
            .in2(_gnd_net_),
            .in3(N__22825),
            .lcout(\line_buffer.n3549 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_2276_LC_20_15_5 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_2276_LC_20_15_5 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_2276_LC_20_15_5 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \line_buffer.TX_ADDR_12__bdd_4_lut_2276_LC_20_15_5  (
            .in0(N__21506),
            .in1(N__22839),
            .in2(N__21299),
            .in3(N__21762),
            .lcout(),
            .ltout(\line_buffer.n3611_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i4_LC_20_15_6 .C_ON=1'b0;
    defparam \line_buffer.dout_i4_LC_20_15_6 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i4_LC_20_15_6 .LUT_INIT=16'b1110010111100000;
    LogicCell40 \line_buffer.dout_i4_LC_20_15_6  (
            .in0(N__21283),
            .in1(N__21750),
            .in2(N__21741),
            .in3(N__21549),
            .lcout(TX_DATA_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24209),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.WIRE_OUT_i4_LC_20_17_1 .C_ON=1'b0;
    defparam \tvp_video_buffer.WIRE_OUT_i4_LC_20_17_1 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.WIRE_OUT_i4_LC_20_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.WIRE_OUT_i4_LC_20_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21633),
            .lcout(RX_DATA_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21969),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.BUFFER_0__i13_LC_20_17_2 .C_ON=1'b0;
    defparam \tvp_video_buffer.BUFFER_0__i13_LC_20_17_2 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.BUFFER_0__i13_LC_20_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.BUFFER_0__i13_LC_20_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21585),
            .lcout(\tvp_video_buffer.BUFFER_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21969),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.BUFFER_0__i5_LC_20_17_5 .C_ON=1'b0;
    defparam \tvp_video_buffer.BUFFER_0__i5_LC_20_17_5 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.BUFFER_0__i5_LC_20_17_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \tvp_video_buffer.BUFFER_0__i5_LC_20_17_5  (
            .in0(N__21623),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\tvp_video_buffer.BUFFER_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21969),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2211_3_lut_LC_20_18_0 .C_ON=1'b0;
    defparam \line_buffer.i2211_3_lut_LC_20_18_0 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2211_3_lut_LC_20_18_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \line_buffer.i2211_3_lut_LC_20_18_0  (
            .in0(N__21579),
            .in1(N__21564),
            .in2(_gnd_net_),
            .in3(N__22771),
            .lcout(\line_buffer.n3548 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2236_3_lut_LC_20_20_2 .C_ON=1'b0;
    defparam \line_buffer.i2236_3_lut_LC_20_20_2 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2236_3_lut_LC_20_20_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \line_buffer.i2236_3_lut_LC_20_20_2  (
            .in0(N__21540),
            .in1(N__21528),
            .in2(_gnd_net_),
            .in3(N__22770),
            .lcout(\line_buffer.n3573 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_2271_LC_20_20_7 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_2271_LC_20_20_7 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_2271_LC_20_20_7 .LUT_INIT=16'b1101101010001010;
    LogicCell40 \line_buffer.TX_ADDR_12__bdd_4_lut_2271_LC_20_20_7  (
            .in0(N__21500),
            .in1(N__21324),
            .in2(N__21295),
            .in3(N__22566),
            .lcout(\line_buffer.n3605 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i6_LC_20_21_4 .C_ON=1'b0;
    defparam \line_buffer.dout_i6_LC_20_21_4 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i6_LC_20_21_4 .LUT_INIT=16'b1111110000001010;
    LogicCell40 \line_buffer.dout_i6_LC_20_21_4  (
            .in0(N__22335),
            .in1(N__21312),
            .in2(N__21305),
            .in3(N__21165),
            .lcout(TX_DATA_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23910),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.VGA_R__i5_LC_20_22_1 .C_ON=1'b0;
    defparam \transmit_module.VGA_R__i5_LC_20_22_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.VGA_R__i5_LC_20_22_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.VGA_R__i5_LC_20_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22560),
            .lcout(n1814),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23957),
            .ce(),
            .sr(N__22431));
    defparam \transmit_module.VGA_R__i7_LC_20_22_3 .C_ON=1'b0;
    defparam \transmit_module.VGA_R__i7_LC_20_22_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.VGA_R__i7_LC_20_22_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.VGA_R__i7_LC_20_22_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22494),
            .lcout(n1812),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__23957),
            .ce(),
            .sr(N__22431));
    defparam \line_buffer.i2235_3_lut_LC_20_24_4 .C_ON=1'b0;
    defparam \line_buffer.i2235_3_lut_LC_20_24_4 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2235_3_lut_LC_20_24_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \line_buffer.i2235_3_lut_LC_20_24_4  (
            .in0(N__22362),
            .in1(N__22347),
            .in2(_gnd_net_),
            .in3(N__22807),
            .lcout(\line_buffer.n3572 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_20_30_4.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_20_30_4.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_20_30_4.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_20_30_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.BUFFER_0__i8_LC_21_7_0 .C_ON=1'b0;
    defparam \tvp_video_buffer.BUFFER_0__i8_LC_21_7_0 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.BUFFER_0__i8_LC_21_7_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \tvp_video_buffer.BUFFER_0__i8_LC_21_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22026),
            .lcout(\tvp_video_buffer.BUFFER_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21944),
            .ce(),
            .sr(_gnd_net_));
    defparam \tvp_video_buffer.BUFFER_0__i16_LC_21_8_7 .C_ON=1'b0;
    defparam \tvp_video_buffer.BUFFER_0__i16_LC_21_8_7 .SEQ_MODE=4'b1000;
    defparam \tvp_video_buffer.BUFFER_0__i16_LC_21_8_7 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \tvp_video_buffer.BUFFER_0__i16_LC_21_8_7  (
            .in0(_gnd_net_),
            .in1(N__22011),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\tvp_video_buffer.BUFFER_1_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21949),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.Y_DELTA_PATTERN_i87_LC_21_13_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i87_LC_21_13_2 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i87_LC_21_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i87_LC_21_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21783),
            .lcout(\transmit_module.Y_DELTA_PATTERN_87 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24295),
            .ce(N__23396),
            .sr(N__23281));
    defparam \transmit_module.Y_DELTA_PATTERN_i84_LC_21_14_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i84_LC_21_14_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i84_LC_21_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i84_LC_21_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24381),
            .lcout(\transmit_module.Y_DELTA_PATTERN_84 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24315),
            .ce(N__23397),
            .sr(N__23325));
    defparam \transmit_module.Y_DELTA_PATTERN_i85_LC_21_14_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i85_LC_21_14_2 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i85_LC_21_14_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i85_LC_21_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24369),
            .lcout(\transmit_module.Y_DELTA_PATTERN_85 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24315),
            .ce(N__23397),
            .sr(N__23325));
    defparam \transmit_module.Y_DELTA_PATTERN_i86_LC_21_14_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i86_LC_21_14_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i86_LC_21_14_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i86_LC_21_14_5  (
            .in0(N__24375),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.Y_DELTA_PATTERN_86 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__24315),
            .ce(N__23397),
            .sr(N__23325));
    defparam \line_buffer.i2197_3_lut_LC_21_16_7 .C_ON=1'b0;
    defparam \line_buffer.i2197_3_lut_LC_21_16_7 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2197_3_lut_LC_21_16_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \line_buffer.i2197_3_lut_LC_21_16_7  (
            .in0(N__22768),
            .in1(N__22869),
            .in2(_gnd_net_),
            .in3(N__22854),
            .lcout(\line_buffer.n3534 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2202_3_lut_LC_21_20_3 .C_ON=1'b0;
    defparam \line_buffer.i2202_3_lut_LC_21_20_3 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2202_3_lut_LC_21_20_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \line_buffer.i2202_3_lut_LC_21_20_3  (
            .in0(N__22798),
            .in1(N__22602),
            .in2(_gnd_net_),
            .in3(N__22587),
            .lcout(\line_buffer.n3539 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // main
