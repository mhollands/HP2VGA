// ******************************************************************************

// iCEcube Netlister

// Version:            2017.08.27940

// Build Date:         Sep 11 2017 17:30:03

// File Generated:     Sep 23 2018 23:07:24

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "main" view "INTERFACE"

module main (
    TVP_VIDEO,
    ADV_B,
    ADV_G,
    ADV_R,
    DEBUG,
    TVP_CLK,
    ADV_CLK,
    TVP_HSYNC,
    ADV_HSYNC,
    TVP_VSYNC,
    ADV_VSYNC,
    ADV_BLANK_N,
    LED,
    ADV_SYNC_N);

    input [9:0] TVP_VIDEO;
    output [7:0] ADV_B;
    output [7:0] ADV_G;
    output [7:0] ADV_R;
    inout [7:0] DEBUG;
    input TVP_CLK;
    output ADV_CLK;
    input TVP_HSYNC;
    output ADV_HSYNC;
    input TVP_VSYNC;
    output ADV_VSYNC;
    output ADV_BLANK_N;
    output LED;
    output ADV_SYNC_N;

    wire N__24376;
    wire N__24375;
    wire N__24374;
    wire N__24365;
    wire N__24364;
    wire N__24363;
    wire N__24356;
    wire N__24355;
    wire N__24354;
    wire N__24347;
    wire N__24346;
    wire N__24345;
    wire N__24338;
    wire N__24337;
    wire N__24336;
    wire N__24329;
    wire N__24328;
    wire N__24327;
    wire N__24320;
    wire N__24319;
    wire N__24318;
    wire N__24311;
    wire N__24310;
    wire N__24309;
    wire N__24302;
    wire N__24301;
    wire N__24300;
    wire N__24293;
    wire N__24292;
    wire N__24291;
    wire N__24284;
    wire N__24283;
    wire N__24282;
    wire N__24275;
    wire N__24274;
    wire N__24273;
    wire N__24266;
    wire N__24265;
    wire N__24264;
    wire N__24257;
    wire N__24256;
    wire N__24255;
    wire N__24248;
    wire N__24247;
    wire N__24246;
    wire N__24239;
    wire N__24238;
    wire N__24237;
    wire N__24230;
    wire N__24229;
    wire N__24228;
    wire N__24221;
    wire N__24220;
    wire N__24219;
    wire N__24212;
    wire N__24211;
    wire N__24210;
    wire N__24203;
    wire N__24202;
    wire N__24201;
    wire N__24194;
    wire N__24193;
    wire N__24192;
    wire N__24185;
    wire N__24184;
    wire N__24183;
    wire N__24176;
    wire N__24175;
    wire N__24174;
    wire N__24167;
    wire N__24166;
    wire N__24165;
    wire N__24158;
    wire N__24157;
    wire N__24156;
    wire N__24149;
    wire N__24148;
    wire N__24147;
    wire N__24140;
    wire N__24139;
    wire N__24138;
    wire N__24131;
    wire N__24130;
    wire N__24129;
    wire N__24122;
    wire N__24121;
    wire N__24120;
    wire N__24113;
    wire N__24112;
    wire N__24111;
    wire N__24104;
    wire N__24103;
    wire N__24102;
    wire N__24095;
    wire N__24094;
    wire N__24093;
    wire N__24086;
    wire N__24085;
    wire N__24084;
    wire N__24077;
    wire N__24076;
    wire N__24075;
    wire N__24068;
    wire N__24067;
    wire N__24066;
    wire N__24059;
    wire N__24058;
    wire N__24057;
    wire N__24050;
    wire N__24049;
    wire N__24048;
    wire N__24041;
    wire N__24040;
    wire N__24039;
    wire N__24032;
    wire N__24031;
    wire N__24030;
    wire N__24023;
    wire N__24022;
    wire N__24021;
    wire N__24014;
    wire N__24013;
    wire N__24012;
    wire N__24005;
    wire N__24004;
    wire N__24003;
    wire N__23996;
    wire N__23995;
    wire N__23994;
    wire N__23987;
    wire N__23986;
    wire N__23985;
    wire N__23978;
    wire N__23977;
    wire N__23976;
    wire N__23969;
    wire N__23968;
    wire N__23967;
    wire N__23960;
    wire N__23959;
    wire N__23958;
    wire N__23951;
    wire N__23950;
    wire N__23949;
    wire N__23942;
    wire N__23941;
    wire N__23940;
    wire N__23923;
    wire N__23920;
    wire N__23917;
    wire N__23914;
    wire N__23911;
    wire N__23908;
    wire N__23905;
    wire N__23902;
    wire N__23899;
    wire N__23896;
    wire N__23893;
    wire N__23890;
    wire N__23887;
    wire N__23884;
    wire N__23881;
    wire N__23878;
    wire N__23875;
    wire N__23872;
    wire N__23869;
    wire N__23866;
    wire N__23863;
    wire N__23860;
    wire N__23859;
    wire N__23856;
    wire N__23855;
    wire N__23852;
    wire N__23851;
    wire N__23850;
    wire N__23849;
    wire N__23848;
    wire N__23847;
    wire N__23846;
    wire N__23845;
    wire N__23844;
    wire N__23843;
    wire N__23842;
    wire N__23841;
    wire N__23840;
    wire N__23839;
    wire N__23838;
    wire N__23837;
    wire N__23836;
    wire N__23833;
    wire N__23830;
    wire N__23829;
    wire N__23828;
    wire N__23825;
    wire N__23822;
    wire N__23819;
    wire N__23818;
    wire N__23813;
    wire N__23808;
    wire N__23807;
    wire N__23806;
    wire N__23803;
    wire N__23800;
    wire N__23795;
    wire N__23790;
    wire N__23783;
    wire N__23780;
    wire N__23775;
    wire N__23772;
    wire N__23769;
    wire N__23762;
    wire N__23759;
    wire N__23756;
    wire N__23753;
    wire N__23750;
    wire N__23747;
    wire N__23742;
    wire N__23741;
    wire N__23736;
    wire N__23731;
    wire N__23720;
    wire N__23715;
    wire N__23712;
    wire N__23709;
    wire N__23706;
    wire N__23703;
    wire N__23700;
    wire N__23697;
    wire N__23694;
    wire N__23685;
    wire N__23674;
    wire N__23671;
    wire N__23668;
    wire N__23665;
    wire N__23662;
    wire N__23659;
    wire N__23656;
    wire N__23653;
    wire N__23650;
    wire N__23647;
    wire N__23644;
    wire N__23641;
    wire N__23638;
    wire N__23635;
    wire N__23632;
    wire N__23629;
    wire N__23626;
    wire N__23623;
    wire N__23620;
    wire N__23617;
    wire N__23614;
    wire N__23613;
    wire N__23612;
    wire N__23611;
    wire N__23608;
    wire N__23605;
    wire N__23604;
    wire N__23603;
    wire N__23602;
    wire N__23601;
    wire N__23600;
    wire N__23599;
    wire N__23598;
    wire N__23595;
    wire N__23592;
    wire N__23591;
    wire N__23590;
    wire N__23587;
    wire N__23586;
    wire N__23583;
    wire N__23578;
    wire N__23577;
    wire N__23576;
    wire N__23573;
    wire N__23570;
    wire N__23563;
    wire N__23560;
    wire N__23557;
    wire N__23554;
    wire N__23553;
    wire N__23550;
    wire N__23547;
    wire N__23544;
    wire N__23543;
    wire N__23540;
    wire N__23537;
    wire N__23536;
    wire N__23535;
    wire N__23532;
    wire N__23529;
    wire N__23522;
    wire N__23519;
    wire N__23518;
    wire N__23513;
    wire N__23510;
    wire N__23503;
    wire N__23500;
    wire N__23497;
    wire N__23494;
    wire N__23493;
    wire N__23492;
    wire N__23489;
    wire N__23486;
    wire N__23485;
    wire N__23482;
    wire N__23479;
    wire N__23474;
    wire N__23471;
    wire N__23468;
    wire N__23465;
    wire N__23462;
    wire N__23459;
    wire N__23454;
    wire N__23449;
    wire N__23444;
    wire N__23441;
    wire N__23438;
    wire N__23431;
    wire N__23422;
    wire N__23419;
    wire N__23414;
    wire N__23401;
    wire N__23398;
    wire N__23395;
    wire N__23394;
    wire N__23391;
    wire N__23388;
    wire N__23387;
    wire N__23386;
    wire N__23385;
    wire N__23380;
    wire N__23377;
    wire N__23374;
    wire N__23373;
    wire N__23372;
    wire N__23371;
    wire N__23370;
    wire N__23367;
    wire N__23360;
    wire N__23357;
    wire N__23354;
    wire N__23353;
    wire N__23352;
    wire N__23349;
    wire N__23346;
    wire N__23345;
    wire N__23344;
    wire N__23343;
    wire N__23340;
    wire N__23333;
    wire N__23330;
    wire N__23327;
    wire N__23326;
    wire N__23325;
    wire N__23324;
    wire N__23323;
    wire N__23318;
    wire N__23315;
    wire N__23312;
    wire N__23311;
    wire N__23310;
    wire N__23309;
    wire N__23308;
    wire N__23307;
    wire N__23306;
    wire N__23305;
    wire N__23304;
    wire N__23303;
    wire N__23300;
    wire N__23299;
    wire N__23296;
    wire N__23289;
    wire N__23286;
    wire N__23283;
    wire N__23282;
    wire N__23281;
    wire N__23278;
    wire N__23275;
    wire N__23268;
    wire N__23265;
    wire N__23262;
    wire N__23261;
    wire N__23260;
    wire N__23257;
    wire N__23256;
    wire N__23253;
    wire N__23252;
    wire N__23249;
    wire N__23246;
    wire N__23245;
    wire N__23242;
    wire N__23239;
    wire N__23238;
    wire N__23235;
    wire N__23232;
    wire N__23229;
    wire N__23228;
    wire N__23227;
    wire N__23224;
    wire N__23217;
    wire N__23214;
    wire N__23211;
    wire N__23206;
    wire N__23199;
    wire N__23196;
    wire N__23193;
    wire N__23192;
    wire N__23191;
    wire N__23190;
    wire N__23189;
    wire N__23178;
    wire N__23175;
    wire N__23164;
    wire N__23161;
    wire N__23158;
    wire N__23155;
    wire N__23152;
    wire N__23143;
    wire N__23140;
    wire N__23139;
    wire N__23138;
    wire N__23131;
    wire N__23128;
    wire N__23125;
    wire N__23124;
    wire N__23121;
    wire N__23118;
    wire N__23117;
    wire N__23112;
    wire N__23109;
    wire N__23098;
    wire N__23095;
    wire N__23092;
    wire N__23089;
    wire N__23082;
    wire N__23079;
    wire N__23074;
    wire N__23071;
    wire N__23068;
    wire N__23065;
    wire N__23062;
    wire N__23055;
    wire N__23046;
    wire N__23043;
    wire N__23040;
    wire N__23037;
    wire N__23032;
    wire N__23029;
    wire N__23026;
    wire N__23023;
    wire N__23020;
    wire N__23011;
    wire N__23008;
    wire N__23005;
    wire N__23002;
    wire N__22999;
    wire N__22996;
    wire N__22993;
    wire N__22990;
    wire N__22987;
    wire N__22984;
    wire N__22981;
    wire N__22978;
    wire N__22975;
    wire N__22972;
    wire N__22969;
    wire N__22966;
    wire N__22963;
    wire N__22960;
    wire N__22957;
    wire N__22954;
    wire N__22951;
    wire N__22948;
    wire N__22945;
    wire N__22942;
    wire N__22939;
    wire N__22936;
    wire N__22933;
    wire N__22930;
    wire N__22927;
    wire N__22924;
    wire N__22921;
    wire N__22918;
    wire N__22915;
    wire N__22912;
    wire N__22909;
    wire N__22906;
    wire N__22903;
    wire N__22900;
    wire N__22897;
    wire N__22894;
    wire N__22891;
    wire N__22888;
    wire N__22885;
    wire N__22882;
    wire N__22879;
    wire N__22876;
    wire N__22873;
    wire N__22870;
    wire N__22869;
    wire N__22866;
    wire N__22865;
    wire N__22862;
    wire N__22859;
    wire N__22858;
    wire N__22857;
    wire N__22856;
    wire N__22853;
    wire N__22850;
    wire N__22847;
    wire N__22846;
    wire N__22843;
    wire N__22842;
    wire N__22839;
    wire N__22836;
    wire N__22835;
    wire N__22830;
    wire N__22829;
    wire N__22826;
    wire N__22823;
    wire N__22820;
    wire N__22819;
    wire N__22818;
    wire N__22815;
    wire N__22812;
    wire N__22809;
    wire N__22806;
    wire N__22803;
    wire N__22802;
    wire N__22799;
    wire N__22794;
    wire N__22793;
    wire N__22790;
    wire N__22787;
    wire N__22784;
    wire N__22779;
    wire N__22776;
    wire N__22771;
    wire N__22768;
    wire N__22765;
    wire N__22764;
    wire N__22761;
    wire N__22758;
    wire N__22755;
    wire N__22748;
    wire N__22741;
    wire N__22738;
    wire N__22735;
    wire N__22726;
    wire N__22723;
    wire N__22714;
    wire N__22711;
    wire N__22708;
    wire N__22705;
    wire N__22702;
    wire N__22699;
    wire N__22696;
    wire N__22693;
    wire N__22690;
    wire N__22689;
    wire N__22688;
    wire N__22685;
    wire N__22684;
    wire N__22681;
    wire N__22678;
    wire N__22677;
    wire N__22676;
    wire N__22675;
    wire N__22672;
    wire N__22669;
    wire N__22668;
    wire N__22665;
    wire N__22662;
    wire N__22659;
    wire N__22656;
    wire N__22655;
    wire N__22654;
    wire N__22651;
    wire N__22650;
    wire N__22649;
    wire N__22644;
    wire N__22641;
    wire N__22640;
    wire N__22633;
    wire N__22630;
    wire N__22627;
    wire N__22624;
    wire N__22623;
    wire N__22622;
    wire N__22621;
    wire N__22620;
    wire N__22619;
    wire N__22616;
    wire N__22613;
    wire N__22610;
    wire N__22609;
    wire N__22604;
    wire N__22601;
    wire N__22600;
    wire N__22593;
    wire N__22590;
    wire N__22587;
    wire N__22584;
    wire N__22583;
    wire N__22582;
    wire N__22581;
    wire N__22580;
    wire N__22579;
    wire N__22578;
    wire N__22575;
    wire N__22574;
    wire N__22573;
    wire N__22572;
    wire N__22569;
    wire N__22566;
    wire N__22565;
    wire N__22564;
    wire N__22563;
    wire N__22562;
    wire N__22561;
    wire N__22560;
    wire N__22555;
    wire N__22552;
    wire N__22549;
    wire N__22548;
    wire N__22547;
    wire N__22542;
    wire N__22539;
    wire N__22538;
    wire N__22537;
    wire N__22536;
    wire N__22535;
    wire N__22534;
    wire N__22533;
    wire N__22526;
    wire N__22523;
    wire N__22520;
    wire N__22517;
    wire N__22516;
    wire N__22515;
    wire N__22514;
    wire N__22513;
    wire N__22512;
    wire N__22509;
    wire N__22506;
    wire N__22503;
    wire N__22500;
    wire N__22499;
    wire N__22498;
    wire N__22495;
    wire N__22492;
    wire N__22489;
    wire N__22488;
    wire N__22487;
    wire N__22486;
    wire N__22483;
    wire N__22478;
    wire N__22475;
    wire N__22474;
    wire N__22471;
    wire N__22470;
    wire N__22467;
    wire N__22466;
    wire N__22465;
    wire N__22462;
    wire N__22459;
    wire N__22456;
    wire N__22449;
    wire N__22446;
    wire N__22445;
    wire N__22444;
    wire N__22441;
    wire N__22440;
    wire N__22439;
    wire N__22438;
    wire N__22437;
    wire N__22436;
    wire N__22435;
    wire N__22434;
    wire N__22429;
    wire N__22426;
    wire N__22423;
    wire N__22422;
    wire N__22421;
    wire N__22420;
    wire N__22419;
    wire N__22416;
    wire N__22413;
    wire N__22410;
    wire N__22409;
    wire N__22408;
    wire N__22407;
    wire N__22404;
    wire N__22397;
    wire N__22394;
    wire N__22391;
    wire N__22388;
    wire N__22387;
    wire N__22386;
    wire N__22383;
    wire N__22380;
    wire N__22377;
    wire N__22374;
    wire N__22371;
    wire N__22366;
    wire N__22363;
    wire N__22360;
    wire N__22353;
    wire N__22352;
    wire N__22349;
    wire N__22348;
    wire N__22347;
    wire N__22344;
    wire N__22341;
    wire N__22340;
    wire N__22337;
    wire N__22332;
    wire N__22329;
    wire N__22326;
    wire N__22323;
    wire N__22322;
    wire N__22319;
    wire N__22316;
    wire N__22315;
    wire N__22314;
    wire N__22311;
    wire N__22308;
    wire N__22303;
    wire N__22298;
    wire N__22295;
    wire N__22292;
    wire N__22289;
    wire N__22286;
    wire N__22283;
    wire N__22282;
    wire N__22279;
    wire N__22276;
    wire N__22273;
    wire N__22270;
    wire N__22267;
    wire N__22266;
    wire N__22263;
    wire N__22258;
    wire N__22255;
    wire N__22252;
    wire N__22249;
    wire N__22248;
    wire N__22247;
    wire N__22244;
    wire N__22243;
    wire N__22240;
    wire N__22239;
    wire N__22234;
    wire N__22231;
    wire N__22230;
    wire N__22229;
    wire N__22226;
    wire N__22225;
    wire N__22222;
    wire N__22219;
    wire N__22212;
    wire N__22209;
    wire N__22206;
    wire N__22205;
    wire N__22202;
    wire N__22199;
    wire N__22196;
    wire N__22193;
    wire N__22180;
    wire N__22177;
    wire N__22174;
    wire N__22171;
    wire N__22168;
    wire N__22165;
    wire N__22162;
    wire N__22159;
    wire N__22154;
    wire N__22151;
    wire N__22146;
    wire N__22143;
    wire N__22140;
    wire N__22137;
    wire N__22134;
    wire N__22131;
    wire N__22128;
    wire N__22117;
    wire N__22112;
    wire N__22109;
    wire N__22106;
    wire N__22101;
    wire N__22096;
    wire N__22093;
    wire N__22090;
    wire N__22083;
    wire N__22080;
    wire N__22077;
    wire N__22074;
    wire N__22071;
    wire N__22070;
    wire N__22069;
    wire N__22066;
    wire N__22063;
    wire N__22062;
    wire N__22061;
    wire N__22058;
    wire N__22055;
    wire N__22050;
    wire N__22047;
    wire N__22044;
    wire N__22041;
    wire N__22038;
    wire N__22037;
    wire N__22034;
    wire N__22031;
    wire N__22024;
    wire N__22021;
    wire N__22020;
    wire N__22017;
    wire N__22006;
    wire N__21999;
    wire N__21992;
    wire N__21985;
    wire N__21982;
    wire N__21977;
    wire N__21972;
    wire N__21965;
    wire N__21960;
    wire N__21959;
    wire N__21958;
    wire N__21949;
    wire N__21938;
    wire N__21935;
    wire N__21932;
    wire N__21927;
    wire N__21924;
    wire N__21921;
    wire N__21918;
    wire N__21915;
    wire N__21908;
    wire N__21903;
    wire N__21900;
    wire N__21897;
    wire N__21894;
    wire N__21891;
    wire N__21888;
    wire N__21885;
    wire N__21882;
    wire N__21875;
    wire N__21870;
    wire N__21865;
    wire N__21860;
    wire N__21857;
    wire N__21854;
    wire N__21845;
    wire N__21838;
    wire N__21833;
    wire N__21830;
    wire N__21825;
    wire N__21820;
    wire N__21815;
    wire N__21812;
    wire N__21809;
    wire N__21806;
    wire N__21801;
    wire N__21798;
    wire N__21793;
    wire N__21788;
    wire N__21785;
    wire N__21780;
    wire N__21773;
    wire N__21768;
    wire N__21765;
    wire N__21762;
    wire N__21757;
    wire N__21752;
    wire N__21739;
    wire N__21736;
    wire N__21733;
    wire N__21730;
    wire N__21727;
    wire N__21724;
    wire N__21721;
    wire N__21718;
    wire N__21715;
    wire N__21712;
    wire N__21709;
    wire N__21706;
    wire N__21703;
    wire N__21700;
    wire N__21697;
    wire N__21694;
    wire N__21691;
    wire N__21688;
    wire N__21685;
    wire N__21682;
    wire N__21679;
    wire N__21676;
    wire N__21673;
    wire N__21670;
    wire N__21667;
    wire N__21664;
    wire N__21661;
    wire N__21658;
    wire N__21655;
    wire N__21652;
    wire N__21649;
    wire N__21646;
    wire N__21643;
    wire N__21640;
    wire N__21637;
    wire N__21634;
    wire N__21631;
    wire N__21628;
    wire N__21625;
    wire N__21622;
    wire N__21619;
    wire N__21616;
    wire N__21613;
    wire N__21610;
    wire N__21607;
    wire N__21604;
    wire N__21601;
    wire N__21598;
    wire N__21595;
    wire N__21592;
    wire N__21589;
    wire N__21586;
    wire N__21583;
    wire N__21580;
    wire N__21577;
    wire N__21574;
    wire N__21571;
    wire N__21568;
    wire N__21565;
    wire N__21562;
    wire N__21559;
    wire N__21556;
    wire N__21553;
    wire N__21550;
    wire N__21547;
    wire N__21544;
    wire N__21541;
    wire N__21538;
    wire N__21535;
    wire N__21532;
    wire N__21529;
    wire N__21526;
    wire N__21523;
    wire N__21520;
    wire N__21517;
    wire N__21514;
    wire N__21511;
    wire N__21508;
    wire N__21505;
    wire N__21502;
    wire N__21499;
    wire N__21496;
    wire N__21493;
    wire N__21490;
    wire N__21489;
    wire N__21488;
    wire N__21487;
    wire N__21484;
    wire N__21481;
    wire N__21480;
    wire N__21477;
    wire N__21474;
    wire N__21473;
    wire N__21468;
    wire N__21465;
    wire N__21464;
    wire N__21463;
    wire N__21460;
    wire N__21459;
    wire N__21458;
    wire N__21457;
    wire N__21456;
    wire N__21453;
    wire N__21450;
    wire N__21447;
    wire N__21444;
    wire N__21441;
    wire N__21438;
    wire N__21437;
    wire N__21436;
    wire N__21433;
    wire N__21430;
    wire N__21427;
    wire N__21424;
    wire N__21421;
    wire N__21416;
    wire N__21409;
    wire N__21406;
    wire N__21403;
    wire N__21400;
    wire N__21395;
    wire N__21392;
    wire N__21389;
    wire N__21386;
    wire N__21379;
    wire N__21374;
    wire N__21371;
    wire N__21368;
    wire N__21365;
    wire N__21360;
    wire N__21357;
    wire N__21346;
    wire N__21345;
    wire N__21344;
    wire N__21343;
    wire N__21342;
    wire N__21341;
    wire N__21340;
    wire N__21339;
    wire N__21338;
    wire N__21337;
    wire N__21336;
    wire N__21335;
    wire N__21332;
    wire N__21329;
    wire N__21326;
    wire N__21325;
    wire N__21324;
    wire N__21323;
    wire N__21322;
    wire N__21321;
    wire N__21318;
    wire N__21317;
    wire N__21314;
    wire N__21311;
    wire N__21308;
    wire N__21307;
    wire N__21306;
    wire N__21303;
    wire N__21300;
    wire N__21297;
    wire N__21296;
    wire N__21295;
    wire N__21294;
    wire N__21293;
    wire N__21292;
    wire N__21289;
    wire N__21288;
    wire N__21285;
    wire N__21282;
    wire N__21281;
    wire N__21280;
    wire N__21279;
    wire N__21278;
    wire N__21273;
    wire N__21270;
    wire N__21269;
    wire N__21268;
    wire N__21267;
    wire N__21266;
    wire N__21263;
    wire N__21262;
    wire N__21261;
    wire N__21260;
    wire N__21259;
    wire N__21256;
    wire N__21253;
    wire N__21252;
    wire N__21251;
    wire N__21248;
    wire N__21245;
    wire N__21242;
    wire N__21237;
    wire N__21234;
    wire N__21231;
    wire N__21228;
    wire N__21225;
    wire N__21220;
    wire N__21219;
    wire N__21218;
    wire N__21217;
    wire N__21214;
    wire N__21211;
    wire N__21210;
    wire N__21209;
    wire N__21206;
    wire N__21203;
    wire N__21200;
    wire N__21199;
    wire N__21198;
    wire N__21197;
    wire N__21196;
    wire N__21195;
    wire N__21194;
    wire N__21191;
    wire N__21188;
    wire N__21185;
    wire N__21182;
    wire N__21181;
    wire N__21180;
    wire N__21179;
    wire N__21176;
    wire N__21173;
    wire N__21172;
    wire N__21171;
    wire N__21168;
    wire N__21167;
    wire N__21166;
    wire N__21163;
    wire N__21158;
    wire N__21155;
    wire N__21152;
    wire N__21151;
    wire N__21148;
    wire N__21147;
    wire N__21144;
    wire N__21141;
    wire N__21138;
    wire N__21135;
    wire N__21132;
    wire N__21129;
    wire N__21124;
    wire N__21121;
    wire N__21118;
    wire N__21115;
    wire N__21108;
    wire N__21097;
    wire N__21094;
    wire N__21093;
    wire N__21092;
    wire N__21087;
    wire N__21084;
    wire N__21081;
    wire N__21078;
    wire N__21063;
    wire N__21060;
    wire N__21057;
    wire N__21056;
    wire N__21055;
    wire N__21052;
    wire N__21049;
    wire N__21046;
    wire N__21041;
    wire N__21038;
    wire N__21037;
    wire N__21036;
    wire N__21035;
    wire N__21034;
    wire N__21033;
    wire N__21030;
    wire N__21027;
    wire N__21024;
    wire N__21019;
    wire N__21016;
    wire N__21013;
    wire N__21010;
    wire N__21007;
    wire N__21000;
    wire N__20997;
    wire N__20994;
    wire N__20991;
    wire N__20988;
    wire N__20985;
    wire N__20976;
    wire N__20973;
    wire N__20970;
    wire N__20959;
    wire N__20956;
    wire N__20955;
    wire N__20952;
    wire N__20949;
    wire N__20946;
    wire N__20937;
    wire N__20932;
    wire N__20929;
    wire N__20926;
    wire N__20923;
    wire N__20920;
    wire N__20915;
    wire N__20912;
    wire N__20909;
    wire N__20906;
    wire N__20903;
    wire N__20896;
    wire N__20889;
    wire N__20886;
    wire N__20881;
    wire N__20874;
    wire N__20871;
    wire N__20862;
    wire N__20853;
    wire N__20850;
    wire N__20845;
    wire N__20838;
    wire N__20835;
    wire N__20832;
    wire N__20829;
    wire N__20824;
    wire N__20811;
    wire N__20808;
    wire N__20805;
    wire N__20802;
    wire N__20797;
    wire N__20794;
    wire N__20787;
    wire N__20776;
    wire N__20761;
    wire N__20758;
    wire N__20755;
    wire N__20752;
    wire N__20749;
    wire N__20746;
    wire N__20743;
    wire N__20740;
    wire N__20737;
    wire N__20734;
    wire N__20731;
    wire N__20728;
    wire N__20725;
    wire N__20722;
    wire N__20719;
    wire N__20716;
    wire N__20713;
    wire N__20710;
    wire N__20707;
    wire N__20704;
    wire N__20701;
    wire N__20698;
    wire N__20695;
    wire N__20692;
    wire N__20689;
    wire N__20686;
    wire N__20683;
    wire N__20680;
    wire N__20677;
    wire N__20674;
    wire N__20671;
    wire N__20668;
    wire N__20665;
    wire N__20662;
    wire N__20659;
    wire N__20656;
    wire N__20653;
    wire N__20650;
    wire N__20647;
    wire N__20644;
    wire N__20641;
    wire N__20638;
    wire N__20635;
    wire N__20632;
    wire N__20629;
    wire N__20626;
    wire N__20623;
    wire N__20622;
    wire N__20619;
    wire N__20618;
    wire N__20615;
    wire N__20614;
    wire N__20611;
    wire N__20608;
    wire N__20607;
    wire N__20606;
    wire N__20603;
    wire N__20600;
    wire N__20599;
    wire N__20598;
    wire N__20597;
    wire N__20596;
    wire N__20591;
    wire N__20588;
    wire N__20587;
    wire N__20584;
    wire N__20583;
    wire N__20578;
    wire N__20575;
    wire N__20572;
    wire N__20569;
    wire N__20566;
    wire N__20565;
    wire N__20560;
    wire N__20557;
    wire N__20554;
    wire N__20551;
    wire N__20550;
    wire N__20547;
    wire N__20542;
    wire N__20539;
    wire N__20536;
    wire N__20533;
    wire N__20530;
    wire N__20527;
    wire N__20522;
    wire N__20519;
    wire N__20514;
    wire N__20511;
    wire N__20508;
    wire N__20505;
    wire N__20496;
    wire N__20485;
    wire N__20482;
    wire N__20479;
    wire N__20476;
    wire N__20473;
    wire N__20470;
    wire N__20467;
    wire N__20464;
    wire N__20461;
    wire N__20458;
    wire N__20455;
    wire N__20452;
    wire N__20449;
    wire N__20446;
    wire N__20443;
    wire N__20440;
    wire N__20437;
    wire N__20434;
    wire N__20431;
    wire N__20428;
    wire N__20425;
    wire N__20422;
    wire N__20419;
    wire N__20416;
    wire N__20413;
    wire N__20410;
    wire N__20407;
    wire N__20404;
    wire N__20401;
    wire N__20398;
    wire N__20395;
    wire N__20392;
    wire N__20389;
    wire N__20386;
    wire N__20383;
    wire N__20380;
    wire N__20377;
    wire N__20374;
    wire N__20371;
    wire N__20368;
    wire N__20365;
    wire N__20362;
    wire N__20359;
    wire N__20356;
    wire N__20353;
    wire N__20350;
    wire N__20347;
    wire N__20344;
    wire N__20341;
    wire N__20338;
    wire N__20335;
    wire N__20332;
    wire N__20329;
    wire N__20326;
    wire N__20323;
    wire N__20320;
    wire N__20317;
    wire N__20314;
    wire N__20311;
    wire N__20308;
    wire N__20305;
    wire N__20302;
    wire N__20299;
    wire N__20296;
    wire N__20293;
    wire N__20290;
    wire N__20287;
    wire N__20284;
    wire N__20281;
    wire N__20278;
    wire N__20275;
    wire N__20274;
    wire N__20271;
    wire N__20268;
    wire N__20265;
    wire N__20260;
    wire N__20259;
    wire N__20256;
    wire N__20253;
    wire N__20250;
    wire N__20245;
    wire N__20242;
    wire N__20241;
    wire N__20240;
    wire N__20239;
    wire N__20236;
    wire N__20233;
    wire N__20230;
    wire N__20229;
    wire N__20228;
    wire N__20225;
    wire N__20220;
    wire N__20217;
    wire N__20216;
    wire N__20215;
    wire N__20210;
    wire N__20209;
    wire N__20202;
    wire N__20199;
    wire N__20198;
    wire N__20197;
    wire N__20196;
    wire N__20195;
    wire N__20194;
    wire N__20193;
    wire N__20192;
    wire N__20191;
    wire N__20188;
    wire N__20185;
    wire N__20182;
    wire N__20179;
    wire N__20176;
    wire N__20171;
    wire N__20170;
    wire N__20169;
    wire N__20168;
    wire N__20167;
    wire N__20166;
    wire N__20153;
    wire N__20150;
    wire N__20139;
    wire N__20132;
    wire N__20127;
    wire N__20116;
    wire N__20115;
    wire N__20112;
    wire N__20109;
    wire N__20106;
    wire N__20103;
    wire N__20100;
    wire N__20097;
    wire N__20094;
    wire N__20091;
    wire N__20088;
    wire N__20085;
    wire N__20082;
    wire N__20079;
    wire N__20076;
    wire N__20073;
    wire N__20070;
    wire N__20067;
    wire N__20064;
    wire N__20061;
    wire N__20058;
    wire N__20055;
    wire N__20052;
    wire N__20049;
    wire N__20046;
    wire N__20043;
    wire N__20040;
    wire N__20037;
    wire N__20034;
    wire N__20031;
    wire N__20028;
    wire N__20025;
    wire N__20022;
    wire N__20019;
    wire N__20016;
    wire N__20013;
    wire N__20010;
    wire N__20007;
    wire N__20004;
    wire N__20001;
    wire N__19998;
    wire N__19995;
    wire N__19992;
    wire N__19989;
    wire N__19986;
    wire N__19983;
    wire N__19980;
    wire N__19977;
    wire N__19974;
    wire N__19971;
    wire N__19968;
    wire N__19965;
    wire N__19962;
    wire N__19959;
    wire N__19956;
    wire N__19953;
    wire N__19950;
    wire N__19947;
    wire N__19944;
    wire N__19941;
    wire N__19938;
    wire N__19935;
    wire N__19932;
    wire N__19929;
    wire N__19926;
    wire N__19923;
    wire N__19920;
    wire N__19917;
    wire N__19912;
    wire N__19909;
    wire N__19906;
    wire N__19903;
    wire N__19900;
    wire N__19897;
    wire N__19894;
    wire N__19891;
    wire N__19888;
    wire N__19885;
    wire N__19882;
    wire N__19881;
    wire N__19878;
    wire N__19877;
    wire N__19876;
    wire N__19875;
    wire N__19874;
    wire N__19871;
    wire N__19870;
    wire N__19869;
    wire N__19866;
    wire N__19863;
    wire N__19860;
    wire N__19857;
    wire N__19854;
    wire N__19853;
    wire N__19850;
    wire N__19847;
    wire N__19844;
    wire N__19841;
    wire N__19836;
    wire N__19831;
    wire N__19828;
    wire N__19825;
    wire N__19822;
    wire N__19819;
    wire N__19814;
    wire N__19809;
    wire N__19804;
    wire N__19799;
    wire N__19796;
    wire N__19789;
    wire N__19786;
    wire N__19783;
    wire N__19780;
    wire N__19777;
    wire N__19774;
    wire N__19771;
    wire N__19768;
    wire N__19765;
    wire N__19762;
    wire N__19759;
    wire N__19756;
    wire N__19753;
    wire N__19750;
    wire N__19747;
    wire N__19744;
    wire N__19741;
    wire N__19738;
    wire N__19735;
    wire N__19732;
    wire N__19729;
    wire N__19726;
    wire N__19723;
    wire N__19720;
    wire N__19717;
    wire N__19716;
    wire N__19715;
    wire N__19714;
    wire N__19713;
    wire N__19710;
    wire N__19707;
    wire N__19702;
    wire N__19701;
    wire N__19698;
    wire N__19697;
    wire N__19694;
    wire N__19693;
    wire N__19692;
    wire N__19691;
    wire N__19686;
    wire N__19683;
    wire N__19680;
    wire N__19677;
    wire N__19674;
    wire N__19671;
    wire N__19670;
    wire N__19667;
    wire N__19664;
    wire N__19663;
    wire N__19662;
    wire N__19661;
    wire N__19658;
    wire N__19651;
    wire N__19646;
    wire N__19643;
    wire N__19638;
    wire N__19635;
    wire N__19632;
    wire N__19629;
    wire N__19626;
    wire N__19623;
    wire N__19612;
    wire N__19603;
    wire N__19600;
    wire N__19597;
    wire N__19594;
    wire N__19591;
    wire N__19588;
    wire N__19587;
    wire N__19584;
    wire N__19583;
    wire N__19582;
    wire N__19579;
    wire N__19576;
    wire N__19573;
    wire N__19572;
    wire N__19569;
    wire N__19566;
    wire N__19563;
    wire N__19560;
    wire N__19557;
    wire N__19552;
    wire N__19543;
    wire N__19540;
    wire N__19537;
    wire N__19534;
    wire N__19533;
    wire N__19532;
    wire N__19529;
    wire N__19526;
    wire N__19525;
    wire N__19522;
    wire N__19521;
    wire N__19520;
    wire N__19517;
    wire N__19514;
    wire N__19513;
    wire N__19512;
    wire N__19511;
    wire N__19508;
    wire N__19505;
    wire N__19502;
    wire N__19501;
    wire N__19500;
    wire N__19497;
    wire N__19496;
    wire N__19495;
    wire N__19494;
    wire N__19493;
    wire N__19492;
    wire N__19487;
    wire N__19480;
    wire N__19477;
    wire N__19472;
    wire N__19471;
    wire N__19470;
    wire N__19469;
    wire N__19468;
    wire N__19467;
    wire N__19462;
    wire N__19459;
    wire N__19448;
    wire N__19443;
    wire N__19438;
    wire N__19433;
    wire N__19426;
    wire N__19411;
    wire N__19410;
    wire N__19407;
    wire N__19404;
    wire N__19401;
    wire N__19398;
    wire N__19397;
    wire N__19394;
    wire N__19391;
    wire N__19388;
    wire N__19381;
    wire N__19378;
    wire N__19375;
    wire N__19372;
    wire N__19369;
    wire N__19368;
    wire N__19367;
    wire N__19366;
    wire N__19365;
    wire N__19364;
    wire N__19363;
    wire N__19362;
    wire N__19361;
    wire N__19360;
    wire N__19359;
    wire N__19356;
    wire N__19355;
    wire N__19354;
    wire N__19353;
    wire N__19352;
    wire N__19351;
    wire N__19350;
    wire N__19349;
    wire N__19348;
    wire N__19347;
    wire N__19346;
    wire N__19345;
    wire N__19344;
    wire N__19343;
    wire N__19342;
    wire N__19341;
    wire N__19340;
    wire N__19339;
    wire N__19338;
    wire N__19337;
    wire N__19336;
    wire N__19335;
    wire N__19334;
    wire N__19333;
    wire N__19332;
    wire N__19331;
    wire N__19330;
    wire N__19329;
    wire N__19328;
    wire N__19327;
    wire N__19326;
    wire N__19325;
    wire N__19324;
    wire N__19323;
    wire N__19322;
    wire N__19321;
    wire N__19228;
    wire N__19225;
    wire N__19222;
    wire N__19219;
    wire N__19216;
    wire N__19215;
    wire N__19212;
    wire N__19209;
    wire N__19206;
    wire N__19203;
    wire N__19200;
    wire N__19197;
    wire N__19192;
    wire N__19189;
    wire N__19186;
    wire N__19183;
    wire N__19180;
    wire N__19177;
    wire N__19174;
    wire N__19171;
    wire N__19168;
    wire N__19165;
    wire N__19162;
    wire N__19159;
    wire N__19156;
    wire N__19153;
    wire N__19150;
    wire N__19147;
    wire N__19144;
    wire N__19141;
    wire N__19138;
    wire N__19135;
    wire N__19132;
    wire N__19129;
    wire N__19128;
    wire N__19127;
    wire N__19126;
    wire N__19123;
    wire N__19122;
    wire N__19121;
    wire N__19120;
    wire N__19117;
    wire N__19114;
    wire N__19111;
    wire N__19108;
    wire N__19105;
    wire N__19104;
    wire N__19103;
    wire N__19102;
    wire N__19101;
    wire N__19100;
    wire N__19099;
    wire N__19096;
    wire N__19095;
    wire N__19092;
    wire N__19089;
    wire N__19084;
    wire N__19079;
    wire N__19076;
    wire N__19071;
    wire N__19068;
    wire N__19065;
    wire N__19058;
    wire N__19053;
    wire N__19042;
    wire N__19037;
    wire N__19030;
    wire N__19027;
    wire N__19026;
    wire N__19023;
    wire N__19022;
    wire N__19021;
    wire N__19018;
    wire N__19013;
    wire N__19010;
    wire N__19003;
    wire N__19000;
    wire N__18997;
    wire N__18994;
    wire N__18991;
    wire N__18988;
    wire N__18987;
    wire N__18984;
    wire N__18983;
    wire N__18982;
    wire N__18979;
    wire N__18976;
    wire N__18971;
    wire N__18968;
    wire N__18961;
    wire N__18960;
    wire N__18957;
    wire N__18954;
    wire N__18949;
    wire N__18946;
    wire N__18943;
    wire N__18942;
    wire N__18939;
    wire N__18936;
    wire N__18933;
    wire N__18930;
    wire N__18927;
    wire N__18924;
    wire N__18921;
    wire N__18918;
    wire N__18915;
    wire N__18912;
    wire N__18909;
    wire N__18906;
    wire N__18903;
    wire N__18900;
    wire N__18897;
    wire N__18894;
    wire N__18891;
    wire N__18888;
    wire N__18885;
    wire N__18882;
    wire N__18879;
    wire N__18876;
    wire N__18873;
    wire N__18870;
    wire N__18867;
    wire N__18864;
    wire N__18861;
    wire N__18858;
    wire N__18855;
    wire N__18852;
    wire N__18849;
    wire N__18846;
    wire N__18843;
    wire N__18840;
    wire N__18837;
    wire N__18834;
    wire N__18831;
    wire N__18828;
    wire N__18825;
    wire N__18822;
    wire N__18819;
    wire N__18816;
    wire N__18813;
    wire N__18810;
    wire N__18807;
    wire N__18804;
    wire N__18801;
    wire N__18798;
    wire N__18795;
    wire N__18792;
    wire N__18789;
    wire N__18786;
    wire N__18783;
    wire N__18780;
    wire N__18777;
    wire N__18774;
    wire N__18771;
    wire N__18768;
    wire N__18765;
    wire N__18762;
    wire N__18759;
    wire N__18756;
    wire N__18753;
    wire N__18750;
    wire N__18747;
    wire N__18744;
    wire N__18739;
    wire N__18736;
    wire N__18733;
    wire N__18732;
    wire N__18729;
    wire N__18726;
    wire N__18723;
    wire N__18718;
    wire N__18715;
    wire N__18712;
    wire N__18711;
    wire N__18708;
    wire N__18705;
    wire N__18702;
    wire N__18699;
    wire N__18696;
    wire N__18693;
    wire N__18690;
    wire N__18687;
    wire N__18684;
    wire N__18681;
    wire N__18678;
    wire N__18675;
    wire N__18672;
    wire N__18669;
    wire N__18666;
    wire N__18663;
    wire N__18660;
    wire N__18657;
    wire N__18654;
    wire N__18651;
    wire N__18648;
    wire N__18645;
    wire N__18642;
    wire N__18639;
    wire N__18636;
    wire N__18633;
    wire N__18630;
    wire N__18627;
    wire N__18624;
    wire N__18621;
    wire N__18618;
    wire N__18615;
    wire N__18612;
    wire N__18609;
    wire N__18606;
    wire N__18603;
    wire N__18600;
    wire N__18597;
    wire N__18594;
    wire N__18591;
    wire N__18588;
    wire N__18585;
    wire N__18582;
    wire N__18579;
    wire N__18576;
    wire N__18573;
    wire N__18570;
    wire N__18567;
    wire N__18564;
    wire N__18561;
    wire N__18558;
    wire N__18555;
    wire N__18552;
    wire N__18549;
    wire N__18546;
    wire N__18543;
    wire N__18540;
    wire N__18537;
    wire N__18534;
    wire N__18531;
    wire N__18528;
    wire N__18525;
    wire N__18522;
    wire N__18519;
    wire N__18516;
    wire N__18513;
    wire N__18510;
    wire N__18507;
    wire N__18504;
    wire N__18499;
    wire N__18496;
    wire N__18493;
    wire N__18490;
    wire N__18487;
    wire N__18484;
    wire N__18481;
    wire N__18478;
    wire N__18475;
    wire N__18472;
    wire N__18469;
    wire N__18466;
    wire N__18465;
    wire N__18464;
    wire N__18461;
    wire N__18458;
    wire N__18457;
    wire N__18454;
    wire N__18451;
    wire N__18448;
    wire N__18445;
    wire N__18442;
    wire N__18433;
    wire N__18430;
    wire N__18427;
    wire N__18424;
    wire N__18421;
    wire N__18420;
    wire N__18417;
    wire N__18414;
    wire N__18411;
    wire N__18408;
    wire N__18407;
    wire N__18406;
    wire N__18403;
    wire N__18400;
    wire N__18397;
    wire N__18394;
    wire N__18385;
    wire N__18382;
    wire N__18379;
    wire N__18376;
    wire N__18375;
    wire N__18374;
    wire N__18373;
    wire N__18370;
    wire N__18367;
    wire N__18364;
    wire N__18361;
    wire N__18352;
    wire N__18349;
    wire N__18346;
    wire N__18343;
    wire N__18340;
    wire N__18337;
    wire N__18334;
    wire N__18331;
    wire N__18328;
    wire N__18325;
    wire N__18322;
    wire N__18321;
    wire N__18320;
    wire N__18319;
    wire N__18316;
    wire N__18313;
    wire N__18310;
    wire N__18307;
    wire N__18302;
    wire N__18299;
    wire N__18292;
    wire N__18291;
    wire N__18288;
    wire N__18285;
    wire N__18282;
    wire N__18279;
    wire N__18274;
    wire N__18271;
    wire N__18268;
    wire N__18265;
    wire N__18262;
    wire N__18261;
    wire N__18258;
    wire N__18255;
    wire N__18252;
    wire N__18249;
    wire N__18246;
    wire N__18243;
    wire N__18240;
    wire N__18237;
    wire N__18234;
    wire N__18231;
    wire N__18228;
    wire N__18225;
    wire N__18222;
    wire N__18219;
    wire N__18216;
    wire N__18213;
    wire N__18210;
    wire N__18207;
    wire N__18204;
    wire N__18201;
    wire N__18198;
    wire N__18195;
    wire N__18192;
    wire N__18189;
    wire N__18186;
    wire N__18183;
    wire N__18180;
    wire N__18177;
    wire N__18174;
    wire N__18171;
    wire N__18168;
    wire N__18165;
    wire N__18162;
    wire N__18159;
    wire N__18156;
    wire N__18153;
    wire N__18150;
    wire N__18147;
    wire N__18144;
    wire N__18141;
    wire N__18138;
    wire N__18135;
    wire N__18132;
    wire N__18129;
    wire N__18126;
    wire N__18123;
    wire N__18120;
    wire N__18117;
    wire N__18114;
    wire N__18111;
    wire N__18108;
    wire N__18105;
    wire N__18102;
    wire N__18099;
    wire N__18096;
    wire N__18093;
    wire N__18090;
    wire N__18087;
    wire N__18084;
    wire N__18081;
    wire N__18078;
    wire N__18075;
    wire N__18072;
    wire N__18069;
    wire N__18066;
    wire N__18063;
    wire N__18060;
    wire N__18057;
    wire N__18052;
    wire N__18049;
    wire N__18046;
    wire N__18043;
    wire N__18040;
    wire N__18037;
    wire N__18034;
    wire N__18031;
    wire N__18028;
    wire N__18025;
    wire N__18022;
    wire N__18019;
    wire N__18016;
    wire N__18013;
    wire N__18010;
    wire N__18007;
    wire N__18004;
    wire N__18001;
    wire N__17998;
    wire N__17995;
    wire N__17992;
    wire N__17989;
    wire N__17986;
    wire N__17983;
    wire N__17980;
    wire N__17977;
    wire N__17974;
    wire N__17971;
    wire N__17968;
    wire N__17965;
    wire N__17962;
    wire N__17959;
    wire N__17956;
    wire N__17955;
    wire N__17952;
    wire N__17951;
    wire N__17948;
    wire N__17945;
    wire N__17944;
    wire N__17941;
    wire N__17938;
    wire N__17935;
    wire N__17932;
    wire N__17925;
    wire N__17920;
    wire N__17917;
    wire N__17914;
    wire N__17911;
    wire N__17908;
    wire N__17905;
    wire N__17902;
    wire N__17899;
    wire N__17896;
    wire N__17893;
    wire N__17890;
    wire N__17887;
    wire N__17886;
    wire N__17885;
    wire N__17884;
    wire N__17881;
    wire N__17878;
    wire N__17873;
    wire N__17866;
    wire N__17863;
    wire N__17860;
    wire N__17857;
    wire N__17854;
    wire N__17851;
    wire N__17848;
    wire N__17845;
    wire N__17842;
    wire N__17839;
    wire N__17838;
    wire N__17835;
    wire N__17832;
    wire N__17829;
    wire N__17824;
    wire N__17823;
    wire N__17822;
    wire N__17821;
    wire N__17818;
    wire N__17815;
    wire N__17812;
    wire N__17809;
    wire N__17804;
    wire N__17797;
    wire N__17794;
    wire N__17791;
    wire N__17788;
    wire N__17785;
    wire N__17782;
    wire N__17779;
    wire N__17776;
    wire N__17773;
    wire N__17770;
    wire N__17767;
    wire N__17764;
    wire N__17761;
    wire N__17758;
    wire N__17757;
    wire N__17756;
    wire N__17753;
    wire N__17750;
    wire N__17747;
    wire N__17742;
    wire N__17741;
    wire N__17738;
    wire N__17735;
    wire N__17732;
    wire N__17725;
    wire N__17722;
    wire N__17719;
    wire N__17716;
    wire N__17713;
    wire N__17712;
    wire N__17709;
    wire N__17708;
    wire N__17705;
    wire N__17704;
    wire N__17701;
    wire N__17698;
    wire N__17695;
    wire N__17692;
    wire N__17683;
    wire N__17680;
    wire N__17677;
    wire N__17674;
    wire N__17671;
    wire N__17668;
    wire N__17665;
    wire N__17662;
    wire N__17659;
    wire N__17656;
    wire N__17653;
    wire N__17650;
    wire N__17647;
    wire N__17644;
    wire N__17641;
    wire N__17638;
    wire N__17635;
    wire N__17632;
    wire N__17629;
    wire N__17626;
    wire N__17623;
    wire N__17620;
    wire N__17617;
    wire N__17614;
    wire N__17611;
    wire N__17608;
    wire N__17605;
    wire N__17602;
    wire N__17599;
    wire N__17596;
    wire N__17593;
    wire N__17590;
    wire N__17587;
    wire N__17584;
    wire N__17583;
    wire N__17582;
    wire N__17579;
    wire N__17578;
    wire N__17575;
    wire N__17572;
    wire N__17571;
    wire N__17568;
    wire N__17565;
    wire N__17562;
    wire N__17559;
    wire N__17556;
    wire N__17551;
    wire N__17548;
    wire N__17541;
    wire N__17536;
    wire N__17535;
    wire N__17532;
    wire N__17529;
    wire N__17526;
    wire N__17521;
    wire N__17518;
    wire N__17515;
    wire N__17512;
    wire N__17509;
    wire N__17506;
    wire N__17503;
    wire N__17502;
    wire N__17499;
    wire N__17498;
    wire N__17497;
    wire N__17494;
    wire N__17491;
    wire N__17488;
    wire N__17485;
    wire N__17476;
    wire N__17475;
    wire N__17472;
    wire N__17471;
    wire N__17470;
    wire N__17467;
    wire N__17464;
    wire N__17461;
    wire N__17458;
    wire N__17449;
    wire N__17446;
    wire N__17443;
    wire N__17442;
    wire N__17441;
    wire N__17438;
    wire N__17437;
    wire N__17434;
    wire N__17431;
    wire N__17426;
    wire N__17419;
    wire N__17416;
    wire N__17413;
    wire N__17412;
    wire N__17409;
    wire N__17408;
    wire N__17407;
    wire N__17404;
    wire N__17401;
    wire N__17398;
    wire N__17395;
    wire N__17386;
    wire N__17383;
    wire N__17380;
    wire N__17377;
    wire N__17374;
    wire N__17371;
    wire N__17370;
    wire N__17367;
    wire N__17364;
    wire N__17359;
    wire N__17356;
    wire N__17353;
    wire N__17350;
    wire N__17347;
    wire N__17344;
    wire N__17343;
    wire N__17340;
    wire N__17337;
    wire N__17332;
    wire N__17331;
    wire N__17328;
    wire N__17325;
    wire N__17320;
    wire N__17317;
    wire N__17314;
    wire N__17311;
    wire N__17308;
    wire N__17305;
    wire N__17302;
    wire N__17299;
    wire N__17296;
    wire N__17293;
    wire N__17290;
    wire N__17287;
    wire N__17284;
    wire N__17281;
    wire N__17278;
    wire N__17275;
    wire N__17272;
    wire N__17269;
    wire N__17266;
    wire N__17263;
    wire N__17260;
    wire N__17257;
    wire N__17254;
    wire N__17251;
    wire N__17248;
    wire N__17245;
    wire N__17242;
    wire N__17239;
    wire N__17236;
    wire N__17233;
    wire N__17230;
    wire N__17227;
    wire N__17224;
    wire N__17221;
    wire N__17218;
    wire N__17215;
    wire N__17212;
    wire N__17209;
    wire N__17206;
    wire N__17203;
    wire N__17200;
    wire N__17197;
    wire N__17194;
    wire N__17191;
    wire N__17188;
    wire N__17187;
    wire N__17184;
    wire N__17181;
    wire N__17176;
    wire N__17173;
    wire N__17172;
    wire N__17169;
    wire N__17166;
    wire N__17161;
    wire N__17158;
    wire N__17157;
    wire N__17154;
    wire N__17151;
    wire N__17146;
    wire N__17143;
    wire N__17140;
    wire N__17139;
    wire N__17136;
    wire N__17133;
    wire N__17128;
    wire N__17125;
    wire N__17122;
    wire N__17119;
    wire N__17118;
    wire N__17113;
    wire N__17110;
    wire N__17107;
    wire N__17106;
    wire N__17103;
    wire N__17100;
    wire N__17099;
    wire N__17098;
    wire N__17097;
    wire N__17094;
    wire N__17091;
    wire N__17084;
    wire N__17077;
    wire N__17074;
    wire N__17073;
    wire N__17072;
    wire N__17071;
    wire N__17068;
    wire N__17065;
    wire N__17062;
    wire N__17057;
    wire N__17050;
    wire N__17049;
    wire N__17048;
    wire N__17047;
    wire N__17044;
    wire N__17041;
    wire N__17036;
    wire N__17029;
    wire N__17028;
    wire N__17027;
    wire N__17026;
    wire N__17023;
    wire N__17020;
    wire N__17015;
    wire N__17008;
    wire N__17005;
    wire N__17004;
    wire N__17001;
    wire N__16998;
    wire N__16995;
    wire N__16992;
    wire N__16987;
    wire N__16986;
    wire N__16983;
    wire N__16980;
    wire N__16975;
    wire N__16974;
    wire N__16971;
    wire N__16968;
    wire N__16965;
    wire N__16962;
    wire N__16959;
    wire N__16956;
    wire N__16953;
    wire N__16950;
    wire N__16947;
    wire N__16944;
    wire N__16941;
    wire N__16938;
    wire N__16935;
    wire N__16932;
    wire N__16929;
    wire N__16926;
    wire N__16923;
    wire N__16920;
    wire N__16917;
    wire N__16914;
    wire N__16911;
    wire N__16908;
    wire N__16905;
    wire N__16902;
    wire N__16899;
    wire N__16896;
    wire N__16893;
    wire N__16890;
    wire N__16887;
    wire N__16884;
    wire N__16881;
    wire N__16878;
    wire N__16875;
    wire N__16872;
    wire N__16869;
    wire N__16866;
    wire N__16863;
    wire N__16860;
    wire N__16857;
    wire N__16854;
    wire N__16851;
    wire N__16848;
    wire N__16845;
    wire N__16842;
    wire N__16839;
    wire N__16836;
    wire N__16833;
    wire N__16830;
    wire N__16827;
    wire N__16824;
    wire N__16821;
    wire N__16818;
    wire N__16815;
    wire N__16812;
    wire N__16809;
    wire N__16806;
    wire N__16803;
    wire N__16800;
    wire N__16797;
    wire N__16794;
    wire N__16791;
    wire N__16788;
    wire N__16785;
    wire N__16782;
    wire N__16779;
    wire N__16776;
    wire N__16773;
    wire N__16770;
    wire N__16765;
    wire N__16762;
    wire N__16761;
    wire N__16760;
    wire N__16757;
    wire N__16756;
    wire N__16755;
    wire N__16752;
    wire N__16749;
    wire N__16746;
    wire N__16743;
    wire N__16740;
    wire N__16729;
    wire N__16726;
    wire N__16723;
    wire N__16720;
    wire N__16719;
    wire N__16718;
    wire N__16717;
    wire N__16714;
    wire N__16713;
    wire N__16712;
    wire N__16709;
    wire N__16706;
    wire N__16705;
    wire N__16702;
    wire N__16699;
    wire N__16694;
    wire N__16689;
    wire N__16686;
    wire N__16683;
    wire N__16678;
    wire N__16675;
    wire N__16668;
    wire N__16663;
    wire N__16660;
    wire N__16657;
    wire N__16654;
    wire N__16653;
    wire N__16650;
    wire N__16647;
    wire N__16642;
    wire N__16639;
    wire N__16638;
    wire N__16635;
    wire N__16632;
    wire N__16629;
    wire N__16626;
    wire N__16623;
    wire N__16620;
    wire N__16617;
    wire N__16614;
    wire N__16611;
    wire N__16608;
    wire N__16605;
    wire N__16602;
    wire N__16599;
    wire N__16596;
    wire N__16593;
    wire N__16590;
    wire N__16587;
    wire N__16584;
    wire N__16581;
    wire N__16578;
    wire N__16575;
    wire N__16572;
    wire N__16569;
    wire N__16566;
    wire N__16563;
    wire N__16560;
    wire N__16557;
    wire N__16554;
    wire N__16551;
    wire N__16548;
    wire N__16545;
    wire N__16542;
    wire N__16539;
    wire N__16536;
    wire N__16533;
    wire N__16530;
    wire N__16527;
    wire N__16524;
    wire N__16521;
    wire N__16518;
    wire N__16515;
    wire N__16512;
    wire N__16509;
    wire N__16506;
    wire N__16503;
    wire N__16500;
    wire N__16497;
    wire N__16494;
    wire N__16491;
    wire N__16488;
    wire N__16485;
    wire N__16482;
    wire N__16479;
    wire N__16476;
    wire N__16473;
    wire N__16470;
    wire N__16467;
    wire N__16464;
    wire N__16461;
    wire N__16458;
    wire N__16455;
    wire N__16452;
    wire N__16449;
    wire N__16446;
    wire N__16443;
    wire N__16440;
    wire N__16435;
    wire N__16432;
    wire N__16429;
    wire N__16426;
    wire N__16423;
    wire N__16420;
    wire N__16417;
    wire N__16414;
    wire N__16413;
    wire N__16410;
    wire N__16407;
    wire N__16404;
    wire N__16401;
    wire N__16398;
    wire N__16393;
    wire N__16392;
    wire N__16389;
    wire N__16386;
    wire N__16381;
    wire N__16378;
    wire N__16377;
    wire N__16374;
    wire N__16371;
    wire N__16366;
    wire N__16363;
    wire N__16360;
    wire N__16357;
    wire N__16354;
    wire N__16351;
    wire N__16348;
    wire N__16345;
    wire N__16342;
    wire N__16341;
    wire N__16338;
    wire N__16335;
    wire N__16332;
    wire N__16327;
    wire N__16324;
    wire N__16321;
    wire N__16320;
    wire N__16317;
    wire N__16314;
    wire N__16309;
    wire N__16308;
    wire N__16305;
    wire N__16302;
    wire N__16299;
    wire N__16296;
    wire N__16293;
    wire N__16290;
    wire N__16287;
    wire N__16284;
    wire N__16281;
    wire N__16278;
    wire N__16275;
    wire N__16272;
    wire N__16269;
    wire N__16266;
    wire N__16263;
    wire N__16260;
    wire N__16257;
    wire N__16254;
    wire N__16251;
    wire N__16248;
    wire N__16245;
    wire N__16242;
    wire N__16239;
    wire N__16236;
    wire N__16233;
    wire N__16230;
    wire N__16227;
    wire N__16224;
    wire N__16221;
    wire N__16218;
    wire N__16215;
    wire N__16212;
    wire N__16209;
    wire N__16206;
    wire N__16203;
    wire N__16200;
    wire N__16197;
    wire N__16194;
    wire N__16191;
    wire N__16188;
    wire N__16185;
    wire N__16182;
    wire N__16179;
    wire N__16176;
    wire N__16173;
    wire N__16170;
    wire N__16167;
    wire N__16164;
    wire N__16161;
    wire N__16158;
    wire N__16155;
    wire N__16152;
    wire N__16149;
    wire N__16146;
    wire N__16143;
    wire N__16140;
    wire N__16137;
    wire N__16134;
    wire N__16131;
    wire N__16128;
    wire N__16125;
    wire N__16122;
    wire N__16119;
    wire N__16116;
    wire N__16113;
    wire N__16110;
    wire N__16107;
    wire N__16104;
    wire N__16101;
    wire N__16098;
    wire N__16093;
    wire N__16090;
    wire N__16087;
    wire N__16084;
    wire N__16081;
    wire N__16078;
    wire N__16075;
    wire N__16072;
    wire N__16069;
    wire N__16066;
    wire N__16063;
    wire N__16060;
    wire N__16057;
    wire N__16054;
    wire N__16051;
    wire N__16048;
    wire N__16045;
    wire N__16042;
    wire N__16039;
    wire N__16038;
    wire N__16037;
    wire N__16036;
    wire N__16033;
    wire N__16030;
    wire N__16029;
    wire N__16026;
    wire N__16025;
    wire N__16022;
    wire N__16019;
    wire N__16016;
    wire N__16013;
    wire N__16010;
    wire N__16007;
    wire N__16004;
    wire N__16001;
    wire N__15996;
    wire N__15993;
    wire N__15990;
    wire N__15983;
    wire N__15978;
    wire N__15973;
    wire N__15970;
    wire N__15967;
    wire N__15964;
    wire N__15961;
    wire N__15958;
    wire N__15955;
    wire N__15952;
    wire N__15949;
    wire N__15948;
    wire N__15945;
    wire N__15942;
    wire N__15939;
    wire N__15934;
    wire N__15931;
    wire N__15930;
    wire N__15929;
    wire N__15928;
    wire N__15927;
    wire N__15924;
    wire N__15923;
    wire N__15922;
    wire N__15921;
    wire N__15918;
    wire N__15915;
    wire N__15908;
    wire N__15901;
    wire N__15892;
    wire N__15891;
    wire N__15890;
    wire N__15889;
    wire N__15888;
    wire N__15887;
    wire N__15886;
    wire N__15885;
    wire N__15882;
    wire N__15879;
    wire N__15872;
    wire N__15865;
    wire N__15856;
    wire N__15853;
    wire N__15852;
    wire N__15849;
    wire N__15848;
    wire N__15845;
    wire N__15844;
    wire N__15843;
    wire N__15842;
    wire N__15839;
    wire N__15836;
    wire N__15833;
    wire N__15830;
    wire N__15827;
    wire N__15824;
    wire N__15821;
    wire N__15818;
    wire N__15815;
    wire N__15808;
    wire N__15807;
    wire N__15806;
    wire N__15803;
    wire N__15796;
    wire N__15795;
    wire N__15792;
    wire N__15789;
    wire N__15786;
    wire N__15783;
    wire N__15776;
    wire N__15769;
    wire N__15766;
    wire N__15763;
    wire N__15762;
    wire N__15761;
    wire N__15760;
    wire N__15759;
    wire N__15758;
    wire N__15757;
    wire N__15756;
    wire N__15755;
    wire N__15752;
    wire N__15749;
    wire N__15746;
    wire N__15739;
    wire N__15732;
    wire N__15721;
    wire N__15720;
    wire N__15719;
    wire N__15716;
    wire N__15713;
    wire N__15712;
    wire N__15709;
    wire N__15704;
    wire N__15701;
    wire N__15698;
    wire N__15693;
    wire N__15690;
    wire N__15687;
    wire N__15684;
    wire N__15681;
    wire N__15678;
    wire N__15675;
    wire N__15670;
    wire N__15667;
    wire N__15664;
    wire N__15661;
    wire N__15658;
    wire N__15655;
    wire N__15652;
    wire N__15649;
    wire N__15648;
    wire N__15645;
    wire N__15642;
    wire N__15639;
    wire N__15636;
    wire N__15633;
    wire N__15630;
    wire N__15627;
    wire N__15624;
    wire N__15621;
    wire N__15618;
    wire N__15615;
    wire N__15612;
    wire N__15609;
    wire N__15606;
    wire N__15603;
    wire N__15600;
    wire N__15597;
    wire N__15594;
    wire N__15591;
    wire N__15588;
    wire N__15585;
    wire N__15582;
    wire N__15579;
    wire N__15576;
    wire N__15573;
    wire N__15570;
    wire N__15567;
    wire N__15564;
    wire N__15561;
    wire N__15558;
    wire N__15555;
    wire N__15552;
    wire N__15549;
    wire N__15546;
    wire N__15543;
    wire N__15540;
    wire N__15537;
    wire N__15534;
    wire N__15531;
    wire N__15528;
    wire N__15525;
    wire N__15522;
    wire N__15519;
    wire N__15516;
    wire N__15513;
    wire N__15510;
    wire N__15507;
    wire N__15504;
    wire N__15501;
    wire N__15498;
    wire N__15495;
    wire N__15492;
    wire N__15489;
    wire N__15486;
    wire N__15483;
    wire N__15480;
    wire N__15477;
    wire N__15474;
    wire N__15471;
    wire N__15468;
    wire N__15465;
    wire N__15462;
    wire N__15459;
    wire N__15456;
    wire N__15453;
    wire N__15450;
    wire N__15445;
    wire N__15442;
    wire N__15441;
    wire N__15440;
    wire N__15435;
    wire N__15432;
    wire N__15429;
    wire N__15426;
    wire N__15423;
    wire N__15420;
    wire N__15417;
    wire N__15414;
    wire N__15411;
    wire N__15408;
    wire N__15403;
    wire N__15400;
    wire N__15397;
    wire N__15396;
    wire N__15393;
    wire N__15390;
    wire N__15387;
    wire N__15384;
    wire N__15381;
    wire N__15378;
    wire N__15375;
    wire N__15372;
    wire N__15369;
    wire N__15366;
    wire N__15363;
    wire N__15360;
    wire N__15357;
    wire N__15354;
    wire N__15351;
    wire N__15348;
    wire N__15345;
    wire N__15342;
    wire N__15339;
    wire N__15336;
    wire N__15333;
    wire N__15330;
    wire N__15327;
    wire N__15324;
    wire N__15321;
    wire N__15318;
    wire N__15315;
    wire N__15312;
    wire N__15309;
    wire N__15306;
    wire N__15303;
    wire N__15300;
    wire N__15297;
    wire N__15294;
    wire N__15291;
    wire N__15288;
    wire N__15285;
    wire N__15282;
    wire N__15279;
    wire N__15276;
    wire N__15273;
    wire N__15270;
    wire N__15267;
    wire N__15264;
    wire N__15261;
    wire N__15258;
    wire N__15255;
    wire N__15252;
    wire N__15249;
    wire N__15246;
    wire N__15243;
    wire N__15240;
    wire N__15237;
    wire N__15234;
    wire N__15231;
    wire N__15228;
    wire N__15225;
    wire N__15222;
    wire N__15219;
    wire N__15216;
    wire N__15213;
    wire N__15210;
    wire N__15207;
    wire N__15204;
    wire N__15201;
    wire N__15198;
    wire N__15195;
    wire N__15192;
    wire N__15189;
    wire N__15186;
    wire N__15185;
    wire N__15182;
    wire N__15179;
    wire N__15176;
    wire N__15171;
    wire N__15166;
    wire N__15163;
    wire N__15162;
    wire N__15159;
    wire N__15156;
    wire N__15153;
    wire N__15150;
    wire N__15147;
    wire N__15144;
    wire N__15141;
    wire N__15138;
    wire N__15135;
    wire N__15132;
    wire N__15129;
    wire N__15126;
    wire N__15123;
    wire N__15120;
    wire N__15117;
    wire N__15114;
    wire N__15111;
    wire N__15108;
    wire N__15105;
    wire N__15102;
    wire N__15099;
    wire N__15096;
    wire N__15093;
    wire N__15090;
    wire N__15087;
    wire N__15084;
    wire N__15081;
    wire N__15078;
    wire N__15075;
    wire N__15072;
    wire N__15069;
    wire N__15066;
    wire N__15063;
    wire N__15060;
    wire N__15057;
    wire N__15054;
    wire N__15051;
    wire N__15048;
    wire N__15045;
    wire N__15042;
    wire N__15039;
    wire N__15036;
    wire N__15033;
    wire N__15030;
    wire N__15027;
    wire N__15024;
    wire N__15021;
    wire N__15018;
    wire N__15015;
    wire N__15012;
    wire N__15009;
    wire N__15006;
    wire N__15003;
    wire N__15000;
    wire N__14997;
    wire N__14994;
    wire N__14991;
    wire N__14988;
    wire N__14985;
    wire N__14982;
    wire N__14979;
    wire N__14976;
    wire N__14973;
    wire N__14970;
    wire N__14967;
    wire N__14964;
    wire N__14961;
    wire N__14958;
    wire N__14955;
    wire N__14954;
    wire N__14951;
    wire N__14948;
    wire N__14945;
    wire N__14942;
    wire N__14939;
    wire N__14932;
    wire N__14929;
    wire N__14926;
    wire N__14925;
    wire N__14922;
    wire N__14919;
    wire N__14916;
    wire N__14913;
    wire N__14910;
    wire N__14907;
    wire N__14904;
    wire N__14901;
    wire N__14898;
    wire N__14895;
    wire N__14892;
    wire N__14889;
    wire N__14886;
    wire N__14883;
    wire N__14880;
    wire N__14877;
    wire N__14874;
    wire N__14871;
    wire N__14868;
    wire N__14865;
    wire N__14862;
    wire N__14859;
    wire N__14856;
    wire N__14853;
    wire N__14850;
    wire N__14847;
    wire N__14844;
    wire N__14841;
    wire N__14838;
    wire N__14835;
    wire N__14832;
    wire N__14829;
    wire N__14826;
    wire N__14823;
    wire N__14820;
    wire N__14817;
    wire N__14814;
    wire N__14811;
    wire N__14808;
    wire N__14805;
    wire N__14802;
    wire N__14799;
    wire N__14796;
    wire N__14793;
    wire N__14790;
    wire N__14787;
    wire N__14784;
    wire N__14781;
    wire N__14778;
    wire N__14775;
    wire N__14772;
    wire N__14769;
    wire N__14766;
    wire N__14763;
    wire N__14760;
    wire N__14757;
    wire N__14754;
    wire N__14751;
    wire N__14748;
    wire N__14745;
    wire N__14742;
    wire N__14739;
    wire N__14736;
    wire N__14733;
    wire N__14730;
    wire N__14727;
    wire N__14724;
    wire N__14723;
    wire N__14720;
    wire N__14717;
    wire N__14714;
    wire N__14711;
    wire N__14708;
    wire N__14701;
    wire N__14698;
    wire N__14695;
    wire N__14692;
    wire N__14689;
    wire N__14686;
    wire N__14683;
    wire N__14680;
    wire N__14677;
    wire N__14674;
    wire N__14671;
    wire N__14668;
    wire N__14665;
    wire N__14662;
    wire N__14659;
    wire N__14656;
    wire N__14653;
    wire N__14650;
    wire N__14647;
    wire N__14644;
    wire N__14641;
    wire N__14638;
    wire N__14635;
    wire N__14632;
    wire N__14629;
    wire N__14626;
    wire N__14623;
    wire N__14620;
    wire N__14617;
    wire N__14614;
    wire N__14611;
    wire N__14608;
    wire N__14605;
    wire N__14604;
    wire N__14601;
    wire N__14598;
    wire N__14595;
    wire N__14592;
    wire N__14587;
    wire N__14584;
    wire N__14581;
    wire N__14578;
    wire N__14575;
    wire N__14572;
    wire N__14569;
    wire N__14566;
    wire N__14563;
    wire N__14560;
    wire N__14557;
    wire N__14554;
    wire N__14551;
    wire N__14548;
    wire N__14545;
    wire N__14542;
    wire N__14539;
    wire N__14536;
    wire N__14533;
    wire N__14530;
    wire N__14527;
    wire N__14524;
    wire N__14521;
    wire N__14520;
    wire N__14517;
    wire N__14514;
    wire N__14513;
    wire N__14508;
    wire N__14505;
    wire N__14502;
    wire N__14499;
    wire N__14496;
    wire N__14493;
    wire N__14490;
    wire N__14487;
    wire N__14482;
    wire N__14479;
    wire N__14476;
    wire N__14473;
    wire N__14470;
    wire N__14467;
    wire N__14464;
    wire N__14463;
    wire N__14462;
    wire N__14459;
    wire N__14456;
    wire N__14453;
    wire N__14450;
    wire N__14447;
    wire N__14444;
    wire N__14441;
    wire N__14438;
    wire N__14435;
    wire N__14432;
    wire N__14429;
    wire N__14426;
    wire N__14419;
    wire N__14416;
    wire N__14415;
    wire N__14412;
    wire N__14411;
    wire N__14408;
    wire N__14405;
    wire N__14402;
    wire N__14399;
    wire N__14396;
    wire N__14393;
    wire N__14390;
    wire N__14387;
    wire N__14384;
    wire N__14381;
    wire N__14378;
    wire N__14375;
    wire N__14372;
    wire N__14367;
    wire N__14364;
    wire N__14359;
    wire N__14356;
    wire N__14353;
    wire N__14352;
    wire N__14351;
    wire N__14348;
    wire N__14345;
    wire N__14342;
    wire N__14339;
    wire N__14336;
    wire N__14333;
    wire N__14330;
    wire N__14327;
    wire N__14324;
    wire N__14321;
    wire N__14318;
    wire N__14315;
    wire N__14310;
    wire N__14305;
    wire N__14304;
    wire N__14301;
    wire N__14300;
    wire N__14297;
    wire N__14294;
    wire N__14291;
    wire N__14288;
    wire N__14285;
    wire N__14282;
    wire N__14279;
    wire N__14276;
    wire N__14273;
    wire N__14270;
    wire N__14267;
    wire N__14264;
    wire N__14261;
    wire N__14254;
    wire N__14251;
    wire N__14248;
    wire N__14245;
    wire N__14244;
    wire N__14243;
    wire N__14240;
    wire N__14237;
    wire N__14234;
    wire N__14231;
    wire N__14228;
    wire N__14225;
    wire N__14222;
    wire N__14219;
    wire N__14216;
    wire N__14213;
    wire N__14210;
    wire N__14207;
    wire N__14204;
    wire N__14201;
    wire N__14198;
    wire N__14193;
    wire N__14188;
    wire N__14185;
    wire N__14182;
    wire N__14181;
    wire N__14178;
    wire N__14175;
    wire N__14172;
    wire N__14171;
    wire N__14168;
    wire N__14165;
    wire N__14162;
    wire N__14159;
    wire N__14156;
    wire N__14153;
    wire N__14150;
    wire N__14147;
    wire N__14144;
    wire N__14141;
    wire N__14138;
    wire N__14135;
    wire N__14132;
    wire N__14127;
    wire N__14122;
    wire N__14121;
    wire N__14118;
    wire N__14115;
    wire N__14110;
    wire N__14107;
    wire N__14106;
    wire N__14103;
    wire N__14100;
    wire N__14095;
    wire N__14094;
    wire N__14091;
    wire N__14088;
    wire N__14085;
    wire N__14082;
    wire N__14079;
    wire N__14076;
    wire N__14073;
    wire N__14070;
    wire N__14067;
    wire N__14064;
    wire N__14061;
    wire N__14058;
    wire N__14055;
    wire N__14052;
    wire N__14049;
    wire N__14046;
    wire N__14043;
    wire N__14040;
    wire N__14037;
    wire N__14034;
    wire N__14031;
    wire N__14028;
    wire N__14025;
    wire N__14022;
    wire N__14019;
    wire N__14016;
    wire N__14013;
    wire N__14010;
    wire N__14007;
    wire N__14004;
    wire N__14001;
    wire N__13998;
    wire N__13995;
    wire N__13992;
    wire N__13989;
    wire N__13986;
    wire N__13983;
    wire N__13980;
    wire N__13977;
    wire N__13974;
    wire N__13971;
    wire N__13968;
    wire N__13965;
    wire N__13962;
    wire N__13959;
    wire N__13956;
    wire N__13953;
    wire N__13950;
    wire N__13947;
    wire N__13944;
    wire N__13941;
    wire N__13938;
    wire N__13935;
    wire N__13932;
    wire N__13929;
    wire N__13926;
    wire N__13923;
    wire N__13920;
    wire N__13917;
    wire N__13914;
    wire N__13911;
    wire N__13908;
    wire N__13905;
    wire N__13902;
    wire N__13899;
    wire N__13896;
    wire N__13893;
    wire N__13890;
    wire N__13887;
    wire N__13884;
    wire N__13881;
    wire N__13876;
    wire N__13873;
    wire N__13870;
    wire N__13867;
    wire N__13864;
    wire N__13861;
    wire N__13858;
    wire N__13855;
    wire N__13852;
    wire N__13849;
    wire N__13846;
    wire N__13843;
    wire N__13840;
    wire N__13837;
    wire N__13836;
    wire N__13835;
    wire N__13834;
    wire N__13827;
    wire N__13824;
    wire N__13821;
    wire N__13816;
    wire N__13813;
    wire N__13812;
    wire N__13811;
    wire N__13808;
    wire N__13807;
    wire N__13804;
    wire N__13797;
    wire N__13792;
    wire N__13789;
    wire N__13786;
    wire N__13785;
    wire N__13784;
    wire N__13783;
    wire N__13780;
    wire N__13773;
    wire N__13768;
    wire N__13765;
    wire N__13762;
    wire N__13761;
    wire N__13758;
    wire N__13755;
    wire N__13754;
    wire N__13753;
    wire N__13748;
    wire N__13745;
    wire N__13742;
    wire N__13739;
    wire N__13736;
    wire N__13733;
    wire N__13726;
    wire N__13723;
    wire N__13720;
    wire N__13717;
    wire N__13714;
    wire N__13711;
    wire N__13708;
    wire N__13705;
    wire N__13702;
    wire N__13699;
    wire N__13696;
    wire N__13693;
    wire N__13690;
    wire N__13687;
    wire N__13684;
    wire N__13683;
    wire N__13682;
    wire N__13681;
    wire N__13678;
    wire N__13673;
    wire N__13670;
    wire N__13663;
    wire N__13660;
    wire N__13659;
    wire N__13656;
    wire N__13655;
    wire N__13654;
    wire N__13651;
    wire N__13646;
    wire N__13643;
    wire N__13636;
    wire N__13633;
    wire N__13632;
    wire N__13631;
    wire N__13630;
    wire N__13627;
    wire N__13624;
    wire N__13621;
    wire N__13618;
    wire N__13609;
    wire N__13606;
    wire N__13605;
    wire N__13604;
    wire N__13603;
    wire N__13600;
    wire N__13593;
    wire N__13588;
    wire N__13585;
    wire N__13584;
    wire N__13583;
    wire N__13582;
    wire N__13579;
    wire N__13574;
    wire N__13571;
    wire N__13564;
    wire N__13561;
    wire N__13560;
    wire N__13559;
    wire N__13558;
    wire N__13555;
    wire N__13550;
    wire N__13547;
    wire N__13540;
    wire N__13537;
    wire N__13536;
    wire N__13535;
    wire N__13534;
    wire N__13529;
    wire N__13526;
    wire N__13523;
    wire N__13516;
    wire N__13513;
    wire N__13510;
    wire N__13509;
    wire N__13508;
    wire N__13507;
    wire N__13504;
    wire N__13501;
    wire N__13496;
    wire N__13489;
    wire N__13486;
    wire N__13485;
    wire N__13482;
    wire N__13479;
    wire N__13476;
    wire N__13475;
    wire N__13474;
    wire N__13471;
    wire N__13468;
    wire N__13465;
    wire N__13462;
    wire N__13455;
    wire N__13452;
    wire N__13449;
    wire N__13446;
    wire N__13443;
    wire N__13440;
    wire N__13435;
    wire N__13432;
    wire N__13429;
    wire N__13426;
    wire N__13425;
    wire N__13424;
    wire N__13419;
    wire N__13416;
    wire N__13413;
    wire N__13408;
    wire N__13407;
    wire N__13404;
    wire N__13401;
    wire N__13396;
    wire N__13393;
    wire N__13390;
    wire N__13389;
    wire N__13388;
    wire N__13381;
    wire N__13378;
    wire N__13375;
    wire N__13374;
    wire N__13373;
    wire N__13366;
    wire N__13363;
    wire N__13360;
    wire N__13357;
    wire N__13356;
    wire N__13353;
    wire N__13350;
    wire N__13345;
    wire N__13344;
    wire N__13343;
    wire N__13342;
    wire N__13333;
    wire N__13330;
    wire N__13327;
    wire N__13326;
    wire N__13321;
    wire N__13318;
    wire N__13315;
    wire N__13312;
    wire N__13309;
    wire N__13306;
    wire N__13303;
    wire N__13300;
    wire N__13297;
    wire N__13294;
    wire N__13291;
    wire N__13288;
    wire N__13285;
    wire N__13282;
    wire N__13279;
    wire N__13276;
    wire N__13273;
    wire N__13270;
    wire N__13267;
    wire N__13264;
    wire N__13261;
    wire N__13258;
    wire N__13255;
    wire N__13254;
    wire N__13253;
    wire N__13250;
    wire N__13245;
    wire N__13240;
    wire N__13237;
    wire N__13234;
    wire N__13231;
    wire N__13228;
    wire N__13225;
    wire N__13222;
    wire N__13221;
    wire N__13220;
    wire N__13217;
    wire N__13212;
    wire N__13207;
    wire N__13206;
    wire N__13203;
    wire N__13200;
    wire N__13197;
    wire N__13194;
    wire N__13191;
    wire N__13188;
    wire N__13185;
    wire N__13182;
    wire N__13179;
    wire N__13176;
    wire N__13173;
    wire N__13170;
    wire N__13167;
    wire N__13164;
    wire N__13161;
    wire N__13158;
    wire N__13155;
    wire N__13152;
    wire N__13149;
    wire N__13146;
    wire N__13143;
    wire N__13140;
    wire N__13137;
    wire N__13134;
    wire N__13131;
    wire N__13128;
    wire N__13125;
    wire N__13122;
    wire N__13119;
    wire N__13116;
    wire N__13113;
    wire N__13110;
    wire N__13107;
    wire N__13104;
    wire N__13101;
    wire N__13098;
    wire N__13095;
    wire N__13092;
    wire N__13089;
    wire N__13086;
    wire N__13083;
    wire N__13080;
    wire N__13077;
    wire N__13074;
    wire N__13071;
    wire N__13068;
    wire N__13065;
    wire N__13062;
    wire N__13059;
    wire N__13056;
    wire N__13053;
    wire N__13050;
    wire N__13047;
    wire N__13044;
    wire N__13041;
    wire N__13038;
    wire N__13035;
    wire N__13032;
    wire N__13029;
    wire N__13026;
    wire N__13023;
    wire N__13020;
    wire N__13017;
    wire N__13014;
    wire N__13011;
    wire N__13008;
    wire N__13005;
    wire N__13002;
    wire N__12999;
    wire N__12996;
    wire N__12993;
    wire N__12990;
    wire N__12987;
    wire N__12982;
    wire N__12979;
    wire N__12976;
    wire N__12973;
    wire N__12970;
    wire N__12967;
    wire N__12964;
    wire N__12963;
    wire N__12960;
    wire N__12957;
    wire N__12952;
    wire N__12949;
    wire N__12948;
    wire N__12945;
    wire N__12942;
    wire N__12939;
    wire N__12936;
    wire N__12933;
    wire N__12930;
    wire N__12927;
    wire N__12924;
    wire N__12921;
    wire N__12918;
    wire N__12915;
    wire N__12912;
    wire N__12909;
    wire N__12906;
    wire N__12903;
    wire N__12900;
    wire N__12897;
    wire N__12894;
    wire N__12891;
    wire N__12888;
    wire N__12885;
    wire N__12882;
    wire N__12879;
    wire N__12876;
    wire N__12873;
    wire N__12870;
    wire N__12867;
    wire N__12864;
    wire N__12861;
    wire N__12858;
    wire N__12855;
    wire N__12852;
    wire N__12849;
    wire N__12846;
    wire N__12843;
    wire N__12840;
    wire N__12837;
    wire N__12834;
    wire N__12831;
    wire N__12828;
    wire N__12825;
    wire N__12822;
    wire N__12819;
    wire N__12816;
    wire N__12813;
    wire N__12810;
    wire N__12807;
    wire N__12804;
    wire N__12801;
    wire N__12798;
    wire N__12795;
    wire N__12792;
    wire N__12789;
    wire N__12786;
    wire N__12783;
    wire N__12780;
    wire N__12777;
    wire N__12774;
    wire N__12771;
    wire N__12768;
    wire N__12765;
    wire N__12762;
    wire N__12759;
    wire N__12756;
    wire N__12753;
    wire N__12750;
    wire N__12747;
    wire N__12744;
    wire N__12741;
    wire N__12736;
    wire N__12733;
    wire N__12730;
    wire N__12727;
    wire N__12724;
    wire N__12721;
    wire N__12718;
    wire N__12715;
    wire N__12712;
    wire N__12709;
    wire N__12706;
    wire N__12703;
    wire N__12700;
    wire N__12697;
    wire N__12694;
    wire N__12691;
    wire N__12688;
    wire N__12685;
    wire N__12682;
    wire N__12679;
    wire N__12676;
    wire N__12673;
    wire N__12670;
    wire N__12667;
    wire N__12664;
    wire N__12661;
    wire N__12658;
    wire N__12657;
    wire N__12656;
    wire N__12653;
    wire N__12650;
    wire N__12647;
    wire N__12646;
    wire N__12643;
    wire N__12638;
    wire N__12635;
    wire N__12632;
    wire N__12627;
    wire N__12624;
    wire N__12621;
    wire N__12618;
    wire N__12615;
    wire N__12610;
    wire N__12607;
    wire N__12606;
    wire N__12605;
    wire N__12602;
    wire N__12599;
    wire N__12598;
    wire N__12595;
    wire N__12592;
    wire N__12589;
    wire N__12586;
    wire N__12583;
    wire N__12578;
    wire N__12575;
    wire N__12570;
    wire N__12567;
    wire N__12562;
    wire N__12559;
    wire N__12556;
    wire N__12553;
    wire N__12550;
    wire N__12547;
    wire N__12546;
    wire N__12545;
    wire N__12544;
    wire N__12543;
    wire N__12532;
    wire N__12529;
    wire N__12526;
    wire N__12523;
    wire N__12520;
    wire N__12517;
    wire N__12516;
    wire N__12513;
    wire N__12512;
    wire N__12509;
    wire N__12508;
    wire N__12507;
    wire N__12506;
    wire N__12503;
    wire N__12500;
    wire N__12491;
    wire N__12484;
    wire N__12481;
    wire N__12478;
    wire N__12475;
    wire N__12472;
    wire N__12469;
    wire N__12468;
    wire N__12465;
    wire N__12462;
    wire N__12459;
    wire N__12456;
    wire N__12453;
    wire N__12450;
    wire N__12447;
    wire N__12444;
    wire N__12441;
    wire N__12438;
    wire N__12435;
    wire N__12432;
    wire N__12429;
    wire N__12426;
    wire N__12423;
    wire N__12420;
    wire N__12417;
    wire N__12414;
    wire N__12411;
    wire N__12408;
    wire N__12405;
    wire N__12402;
    wire N__12399;
    wire N__12396;
    wire N__12393;
    wire N__12390;
    wire N__12387;
    wire N__12384;
    wire N__12381;
    wire N__12378;
    wire N__12375;
    wire N__12372;
    wire N__12369;
    wire N__12366;
    wire N__12363;
    wire N__12360;
    wire N__12357;
    wire N__12354;
    wire N__12351;
    wire N__12348;
    wire N__12345;
    wire N__12342;
    wire N__12339;
    wire N__12336;
    wire N__12333;
    wire N__12330;
    wire N__12327;
    wire N__12324;
    wire N__12321;
    wire N__12318;
    wire N__12315;
    wire N__12312;
    wire N__12309;
    wire N__12306;
    wire N__12303;
    wire N__12300;
    wire N__12297;
    wire N__12294;
    wire N__12291;
    wire N__12288;
    wire N__12285;
    wire N__12282;
    wire N__12279;
    wire N__12276;
    wire N__12273;
    wire N__12270;
    wire N__12267;
    wire N__12264;
    wire N__12261;
    wire N__12258;
    wire N__12253;
    wire N__12250;
    wire N__12247;
    wire N__12244;
    wire N__12241;
    wire N__12238;
    wire N__12237;
    wire N__12236;
    wire N__12235;
    wire N__12234;
    wire N__12231;
    wire N__12222;
    wire N__12219;
    wire N__12214;
    wire N__12213;
    wire N__12210;
    wire N__12207;
    wire N__12204;
    wire N__12201;
    wire N__12198;
    wire N__12195;
    wire N__12192;
    wire N__12189;
    wire N__12186;
    wire N__12183;
    wire N__12180;
    wire N__12177;
    wire N__12174;
    wire N__12171;
    wire N__12168;
    wire N__12165;
    wire N__12162;
    wire N__12159;
    wire N__12156;
    wire N__12153;
    wire N__12150;
    wire N__12147;
    wire N__12144;
    wire N__12141;
    wire N__12138;
    wire N__12135;
    wire N__12132;
    wire N__12129;
    wire N__12126;
    wire N__12123;
    wire N__12120;
    wire N__12117;
    wire N__12114;
    wire N__12111;
    wire N__12108;
    wire N__12105;
    wire N__12102;
    wire N__12099;
    wire N__12096;
    wire N__12093;
    wire N__12090;
    wire N__12087;
    wire N__12084;
    wire N__12081;
    wire N__12078;
    wire N__12075;
    wire N__12072;
    wire N__12069;
    wire N__12066;
    wire N__12063;
    wire N__12060;
    wire N__12057;
    wire N__12054;
    wire N__12051;
    wire N__12048;
    wire N__12045;
    wire N__12042;
    wire N__12039;
    wire N__12036;
    wire N__12033;
    wire N__12030;
    wire N__12027;
    wire N__12024;
    wire N__12021;
    wire N__12018;
    wire N__12015;
    wire N__12012;
    wire N__12009;
    wire N__12006;
    wire N__12003;
    wire N__11998;
    wire N__11995;
    wire N__11992;
    wire N__11989;
    wire N__11988;
    wire N__11987;
    wire N__11986;
    wire N__11983;
    wire N__11978;
    wire N__11975;
    wire N__11968;
    wire N__11965;
    wire N__11962;
    wire N__11959;
    wire N__11958;
    wire N__11955;
    wire N__11952;
    wire N__11949;
    wire N__11946;
    wire N__11943;
    wire N__11940;
    wire N__11937;
    wire N__11934;
    wire N__11931;
    wire N__11928;
    wire N__11925;
    wire N__11922;
    wire N__11919;
    wire N__11916;
    wire N__11913;
    wire N__11910;
    wire N__11907;
    wire N__11904;
    wire N__11901;
    wire N__11898;
    wire N__11895;
    wire N__11892;
    wire N__11889;
    wire N__11886;
    wire N__11883;
    wire N__11880;
    wire N__11877;
    wire N__11874;
    wire N__11871;
    wire N__11868;
    wire N__11865;
    wire N__11862;
    wire N__11859;
    wire N__11856;
    wire N__11853;
    wire N__11850;
    wire N__11847;
    wire N__11844;
    wire N__11841;
    wire N__11838;
    wire N__11835;
    wire N__11832;
    wire N__11829;
    wire N__11826;
    wire N__11823;
    wire N__11820;
    wire N__11817;
    wire N__11814;
    wire N__11811;
    wire N__11808;
    wire N__11805;
    wire N__11802;
    wire N__11799;
    wire N__11796;
    wire N__11793;
    wire N__11790;
    wire N__11787;
    wire N__11784;
    wire N__11781;
    wire N__11778;
    wire N__11775;
    wire N__11772;
    wire N__11769;
    wire N__11766;
    wire N__11763;
    wire N__11760;
    wire N__11757;
    wire N__11754;
    wire N__11751;
    wire N__11748;
    wire N__11745;
    wire N__11742;
    wire N__11739;
    wire N__11734;
    wire N__11731;
    wire N__11728;
    wire N__11725;
    wire N__11722;
    wire N__11719;
    wire N__11716;
    wire N__11713;
    wire N__11710;
    wire N__11709;
    wire N__11706;
    wire N__11703;
    wire N__11700;
    wire N__11695;
    wire N__11692;
    wire N__11691;
    wire N__11688;
    wire N__11685;
    wire N__11682;
    wire N__11679;
    wire N__11676;
    wire N__11673;
    wire N__11668;
    wire N__11665;
    wire N__11662;
    wire N__11659;
    wire N__11656;
    wire N__11655;
    wire N__11652;
    wire N__11649;
    wire N__11646;
    wire N__11643;
    wire N__11640;
    wire N__11637;
    wire N__11634;
    wire N__11631;
    wire N__11628;
    wire N__11625;
    wire N__11622;
    wire N__11619;
    wire N__11616;
    wire N__11613;
    wire N__11610;
    wire N__11607;
    wire N__11604;
    wire N__11601;
    wire N__11598;
    wire N__11595;
    wire N__11592;
    wire N__11589;
    wire N__11586;
    wire N__11583;
    wire N__11580;
    wire N__11577;
    wire N__11574;
    wire N__11571;
    wire N__11568;
    wire N__11565;
    wire N__11562;
    wire N__11559;
    wire N__11556;
    wire N__11553;
    wire N__11550;
    wire N__11547;
    wire N__11544;
    wire N__11541;
    wire N__11538;
    wire N__11535;
    wire N__11532;
    wire N__11529;
    wire N__11526;
    wire N__11523;
    wire N__11520;
    wire N__11517;
    wire N__11514;
    wire N__11511;
    wire N__11508;
    wire N__11505;
    wire N__11502;
    wire N__11499;
    wire N__11496;
    wire N__11493;
    wire N__11490;
    wire N__11487;
    wire N__11484;
    wire N__11481;
    wire N__11478;
    wire N__11475;
    wire N__11472;
    wire N__11469;
    wire N__11466;
    wire N__11463;
    wire N__11460;
    wire N__11457;
    wire N__11454;
    wire N__11451;
    wire N__11448;
    wire N__11445;
    wire N__11440;
    wire N__11437;
    wire N__11434;
    wire N__11431;
    wire N__11428;
    wire N__11427;
    wire N__11424;
    wire N__11421;
    wire N__11418;
    wire N__11415;
    wire N__11412;
    wire N__11409;
    wire N__11406;
    wire N__11403;
    wire N__11400;
    wire N__11397;
    wire N__11394;
    wire N__11391;
    wire N__11388;
    wire N__11385;
    wire N__11382;
    wire N__11379;
    wire N__11376;
    wire N__11373;
    wire N__11370;
    wire N__11367;
    wire N__11364;
    wire N__11361;
    wire N__11358;
    wire N__11355;
    wire N__11352;
    wire N__11349;
    wire N__11346;
    wire N__11343;
    wire N__11340;
    wire N__11337;
    wire N__11334;
    wire N__11331;
    wire N__11328;
    wire N__11325;
    wire N__11322;
    wire N__11319;
    wire N__11316;
    wire N__11313;
    wire N__11310;
    wire N__11307;
    wire N__11304;
    wire N__11301;
    wire N__11298;
    wire N__11295;
    wire N__11292;
    wire N__11289;
    wire N__11286;
    wire N__11283;
    wire N__11280;
    wire N__11277;
    wire N__11274;
    wire N__11271;
    wire N__11268;
    wire N__11265;
    wire N__11262;
    wire N__11259;
    wire N__11256;
    wire N__11253;
    wire N__11250;
    wire N__11247;
    wire N__11244;
    wire N__11241;
    wire N__11238;
    wire N__11235;
    wire N__11232;
    wire N__11229;
    wire N__11226;
    wire N__11223;
    wire N__11220;
    wire N__11217;
    wire N__11212;
    wire N__11209;
    wire N__11208;
    wire N__11205;
    wire N__11202;
    wire N__11199;
    wire N__11196;
    wire N__11193;
    wire N__11190;
    wire N__11187;
    wire N__11184;
    wire N__11181;
    wire N__11178;
    wire N__11175;
    wire N__11172;
    wire N__11169;
    wire N__11166;
    wire N__11163;
    wire N__11160;
    wire N__11157;
    wire N__11154;
    wire N__11151;
    wire N__11148;
    wire N__11145;
    wire N__11142;
    wire N__11139;
    wire N__11136;
    wire N__11133;
    wire N__11130;
    wire N__11127;
    wire N__11124;
    wire N__11121;
    wire N__11118;
    wire N__11115;
    wire N__11112;
    wire N__11109;
    wire N__11106;
    wire N__11103;
    wire N__11100;
    wire N__11097;
    wire N__11094;
    wire N__11091;
    wire N__11088;
    wire N__11085;
    wire N__11082;
    wire N__11079;
    wire N__11076;
    wire N__11073;
    wire N__11070;
    wire N__11067;
    wire N__11064;
    wire N__11061;
    wire N__11058;
    wire N__11055;
    wire N__11052;
    wire N__11049;
    wire N__11046;
    wire N__11043;
    wire N__11040;
    wire N__11037;
    wire N__11034;
    wire N__11031;
    wire N__11028;
    wire N__11025;
    wire N__11022;
    wire N__11019;
    wire N__11016;
    wire N__11013;
    wire N__11010;
    wire N__11007;
    wire N__11004;
    wire N__10999;
    wire N__10996;
    wire N__10993;
    wire N__10990;
    wire N__10987;
    wire N__10984;
    wire N__10981;
    wire N__10978;
    wire N__10975;
    wire N__10972;
    wire N__10969;
    wire N__10966;
    wire N__10963;
    wire N__10960;
    wire N__10957;
    wire N__10954;
    wire N__10951;
    wire N__10948;
    wire N__10945;
    wire N__10942;
    wire N__10939;
    wire N__10936;
    wire N__10933;
    wire N__10930;
    wire N__10927;
    wire N__10924;
    wire N__10923;
    wire N__10922;
    wire N__10919;
    wire N__10916;
    wire N__10913;
    wire N__10910;
    wire N__10903;
    wire N__10902;
    wire N__10901;
    wire N__10898;
    wire N__10895;
    wire N__10892;
    wire N__10885;
    wire N__10882;
    wire N__10879;
    wire N__10876;
    wire N__10873;
    wire N__10870;
    wire N__10869;
    wire N__10866;
    wire N__10863;
    wire N__10860;
    wire N__10857;
    wire N__10854;
    wire N__10851;
    wire N__10848;
    wire N__10845;
    wire N__10842;
    wire N__10839;
    wire N__10836;
    wire N__10833;
    wire N__10830;
    wire N__10827;
    wire N__10824;
    wire N__10821;
    wire N__10818;
    wire N__10815;
    wire N__10812;
    wire N__10809;
    wire N__10806;
    wire N__10803;
    wire N__10800;
    wire N__10797;
    wire N__10794;
    wire N__10791;
    wire N__10788;
    wire N__10785;
    wire N__10782;
    wire N__10779;
    wire N__10776;
    wire N__10773;
    wire N__10770;
    wire N__10767;
    wire N__10764;
    wire N__10761;
    wire N__10758;
    wire N__10755;
    wire N__10752;
    wire N__10749;
    wire N__10746;
    wire N__10743;
    wire N__10740;
    wire N__10737;
    wire N__10734;
    wire N__10731;
    wire N__10728;
    wire N__10725;
    wire N__10722;
    wire N__10719;
    wire N__10716;
    wire N__10713;
    wire N__10710;
    wire N__10707;
    wire N__10704;
    wire N__10701;
    wire N__10698;
    wire N__10695;
    wire N__10692;
    wire N__10689;
    wire N__10686;
    wire N__10683;
    wire N__10680;
    wire N__10677;
    wire N__10674;
    wire N__10671;
    wire N__10668;
    wire N__10665;
    wire N__10660;
    wire N__10657;
    wire N__10654;
    wire N__10651;
    wire N__10648;
    wire N__10645;
    wire N__10642;
    wire N__10639;
    wire N__10636;
    wire N__10633;
    wire N__10630;
    wire N__10627;
    wire N__10624;
    wire N__10623;
    wire N__10620;
    wire N__10617;
    wire N__10612;
    wire N__10609;
    wire N__10608;
    wire N__10605;
    wire N__10602;
    wire N__10597;
    wire N__10594;
    wire N__10591;
    wire N__10588;
    wire N__10585;
    wire N__10584;
    wire N__10581;
    wire N__10578;
    wire N__10575;
    wire N__10572;
    wire N__10569;
    wire N__10566;
    wire N__10561;
    wire N__10560;
    wire N__10559;
    wire N__10556;
    wire N__10555;
    wire N__10552;
    wire N__10549;
    wire N__10546;
    wire N__10543;
    wire N__10534;
    wire N__10531;
    wire N__10528;
    wire N__10527;
    wire N__10524;
    wire N__10521;
    wire N__10520;
    wire N__10517;
    wire N__10516;
    wire N__10513;
    wire N__10510;
    wire N__10507;
    wire N__10504;
    wire N__10495;
    wire N__10494;
    wire N__10491;
    wire N__10488;
    wire N__10483;
    wire N__10482;
    wire N__10481;
    wire N__10478;
    wire N__10475;
    wire N__10472;
    wire N__10465;
    wire N__10462;
    wire N__10459;
    wire N__10456;
    wire N__10453;
    wire N__10450;
    wire N__10447;
    wire N__10444;
    wire N__10443;
    wire N__10440;
    wire N__10437;
    wire N__10432;
    wire N__10429;
    wire N__10428;
    wire N__10427;
    wire N__10424;
    wire N__10423;
    wire N__10420;
    wire N__10417;
    wire N__10412;
    wire N__10405;
    wire N__10402;
    wire N__10401;
    wire N__10400;
    wire N__10399;
    wire N__10396;
    wire N__10393;
    wire N__10388;
    wire N__10381;
    wire N__10378;
    wire N__10375;
    wire N__10372;
    wire N__10371;
    wire N__10370;
    wire N__10367;
    wire N__10364;
    wire N__10361;
    wire N__10354;
    wire N__10351;
    wire N__10350;
    wire N__10349;
    wire N__10346;
    wire N__10341;
    wire N__10336;
    wire N__10333;
    wire N__10330;
    wire N__10327;
    wire N__10324;
    wire N__10321;
    wire N__10318;
    wire N__10315;
    wire N__10312;
    wire N__10309;
    wire N__10306;
    wire N__10303;
    wire N__10300;
    wire N__10297;
    wire N__10294;
    wire N__10291;
    wire N__10290;
    wire N__10285;
    wire N__10282;
    wire N__10279;
    wire N__10276;
    wire N__10273;
    wire N__10270;
    wire N__10269;
    wire N__10266;
    wire N__10263;
    wire N__10262;
    wire N__10257;
    wire N__10254;
    wire N__10253;
    wire N__10248;
    wire N__10245;
    wire N__10240;
    wire N__10237;
    wire N__10234;
    wire N__10231;
    wire N__10228;
    wire N__10227;
    wire N__10226;
    wire N__10225;
    wire N__10222;
    wire N__10219;
    wire N__10216;
    wire N__10213;
    wire N__10206;
    wire N__10203;
    wire N__10198;
    wire N__10195;
    wire N__10192;
    wire N__10189;
    wire N__10188;
    wire N__10185;
    wire N__10182;
    wire N__10181;
    wire N__10180;
    wire N__10175;
    wire N__10172;
    wire N__10169;
    wire N__10164;
    wire N__10161;
    wire N__10158;
    wire N__10155;
    wire N__10152;
    wire N__10149;
    wire N__10146;
    wire N__10143;
    wire N__10140;
    wire N__10135;
    wire N__10132;
    wire N__10129;
    wire N__10126;
    wire N__10123;
    wire N__10120;
    wire N__10117;
    wire N__10114;
    wire N__10113;
    wire N__10112;
    wire N__10109;
    wire N__10106;
    wire N__10105;
    wire N__10102;
    wire N__10099;
    wire N__10096;
    wire N__10093;
    wire N__10090;
    wire N__10083;
    wire N__10078;
    wire N__10075;
    wire N__10072;
    wire N__10069;
    wire N__10066;
    wire N__10063;
    wire N__10060;
    wire N__10057;
    wire N__10054;
    wire N__10051;
    wire N__10048;
    wire N__10047;
    wire N__10044;
    wire N__10041;
    wire N__10040;
    wire N__10037;
    wire N__10034;
    wire N__10031;
    wire N__10026;
    wire N__10023;
    wire N__10020;
    wire N__10017;
    wire N__10012;
    wire N__10009;
    wire N__10006;
    wire N__10003;
    wire N__10000;
    wire N__9997;
    wire N__9994;
    wire N__9991;
    wire N__9988;
    wire N__9985;
    wire N__9982;
    wire N__9979;
    wire N__9976;
    wire N__9975;
    wire N__9972;
    wire N__9969;
    wire N__9966;
    wire N__9963;
    wire N__9960;
    wire N__9957;
    wire N__9954;
    wire N__9951;
    wire N__9948;
    wire N__9945;
    wire N__9942;
    wire N__9939;
    wire N__9936;
    wire N__9933;
    wire N__9930;
    wire N__9927;
    wire N__9924;
    wire N__9921;
    wire N__9918;
    wire N__9915;
    wire N__9912;
    wire N__9909;
    wire N__9906;
    wire N__9903;
    wire N__9900;
    wire N__9897;
    wire N__9894;
    wire N__9891;
    wire N__9888;
    wire N__9885;
    wire N__9882;
    wire N__9879;
    wire N__9876;
    wire N__9873;
    wire N__9870;
    wire N__9867;
    wire N__9864;
    wire N__9861;
    wire N__9858;
    wire N__9855;
    wire N__9852;
    wire N__9849;
    wire N__9846;
    wire N__9843;
    wire N__9840;
    wire N__9837;
    wire N__9834;
    wire N__9831;
    wire N__9828;
    wire N__9825;
    wire N__9822;
    wire N__9819;
    wire N__9816;
    wire N__9813;
    wire N__9810;
    wire N__9807;
    wire N__9804;
    wire N__9801;
    wire N__9798;
    wire N__9795;
    wire N__9792;
    wire N__9789;
    wire N__9786;
    wire N__9783;
    wire N__9780;
    wire N__9777;
    wire N__9772;
    wire N__9769;
    wire N__9768;
    wire N__9765;
    wire N__9762;
    wire N__9757;
    wire N__9754;
    wire N__9751;
    wire N__9748;
    wire N__9745;
    wire N__9742;
    wire N__9739;
    wire N__9736;
    wire N__9733;
    wire N__9730;
    wire N__9727;
    wire N__9724;
    wire N__9721;
    wire N__9718;
    wire N__9715;
    wire N__9712;
    wire N__9709;
    wire N__9706;
    wire N__9703;
    wire N__9700;
    wire N__9697;
    wire N__9694;
    wire N__9691;
    wire N__9688;
    wire N__9685;
    wire N__9682;
    wire N__9679;
    wire N__9676;
    wire N__9673;
    wire N__9672;
    wire N__9669;
    wire N__9666;
    wire N__9663;
    wire N__9660;
    wire N__9657;
    wire N__9654;
    wire N__9651;
    wire N__9648;
    wire N__9643;
    wire N__9640;
    wire N__9637;
    wire N__9634;
    wire N__9631;
    wire N__9628;
    wire N__9625;
    wire N__9622;
    wire N__9621;
    wire N__9620;
    wire N__9619;
    wire N__9616;
    wire N__9613;
    wire N__9610;
    wire N__9607;
    wire N__9598;
    wire N__9595;
    wire N__9594;
    wire N__9593;
    wire N__9592;
    wire N__9589;
    wire N__9586;
    wire N__9583;
    wire N__9580;
    wire N__9577;
    wire N__9568;
    wire N__9565;
    wire N__9564;
    wire N__9563;
    wire N__9562;
    wire N__9559;
    wire N__9556;
    wire N__9553;
    wire N__9550;
    wire N__9541;
    wire N__9538;
    wire N__9537;
    wire N__9536;
    wire N__9535;
    wire N__9532;
    wire N__9527;
    wire N__9524;
    wire N__9517;
    wire N__9514;
    wire N__9513;
    wire N__9512;
    wire N__9509;
    wire N__9506;
    wire N__9503;
    wire N__9496;
    wire N__9493;
    wire N__9492;
    wire N__9489;
    wire N__9488;
    wire N__9485;
    wire N__9482;
    wire N__9479;
    wire N__9472;
    wire N__9469;
    wire N__9468;
    wire N__9467;
    wire N__9466;
    wire N__9463;
    wire N__9458;
    wire N__9455;
    wire N__9448;
    wire N__9445;
    wire N__9444;
    wire N__9443;
    wire N__9442;
    wire N__9439;
    wire N__9436;
    wire N__9433;
    wire N__9430;
    wire N__9421;
    wire N__9418;
    wire N__9415;
    wire N__9412;
    wire N__9409;
    wire N__9406;
    wire N__9403;
    wire N__9400;
    wire N__9397;
    wire N__9394;
    wire N__9391;
    wire N__9388;
    wire N__9385;
    wire N__9382;
    wire N__9379;
    wire N__9376;
    wire N__9373;
    wire N__9370;
    wire N__9367;
    wire N__9364;
    wire N__9361;
    wire N__9358;
    wire N__9355;
    wire N__9352;
    wire N__9349;
    wire N__9346;
    wire N__9343;
    wire N__9340;
    wire N__9337;
    wire N__9334;
    wire N__9331;
    wire N__9328;
    wire N__9325;
    wire N__9322;
    wire N__9319;
    wire N__9316;
    wire N__9313;
    wire N__9310;
    wire N__9309;
    wire N__9308;
    wire N__9307;
    wire N__9304;
    wire N__9301;
    wire N__9298;
    wire N__9295;
    wire N__9286;
    wire N__9283;
    wire N__9280;
    wire N__9277;
    wire N__9274;
    wire N__9271;
    wire N__9268;
    wire N__9265;
    wire N__9262;
    wire N__9259;
    wire N__9256;
    wire N__9253;
    wire N__9250;
    wire N__9247;
    wire N__9244;
    wire N__9241;
    wire N__9238;
    wire N__9235;
    wire N__9232;
    wire N__9229;
    wire N__9226;
    wire N__9223;
    wire N__9220;
    wire N__9217;
    wire N__9214;
    wire N__9211;
    wire N__9208;
    wire N__9205;
    wire N__9202;
    wire N__9199;
    wire N__9196;
    wire N__9193;
    wire N__9190;
    wire N__9187;
    wire N__9184;
    wire N__9181;
    wire N__9178;
    wire N__9175;
    wire N__9172;
    wire N__9169;
    wire N__9166;
    wire N__9163;
    wire N__9160;
    wire N__9157;
    wire N__9154;
    wire N__9151;
    wire N__9148;
    wire N__9145;
    wire N__9142;
    wire N__9139;
    wire N__9136;
    wire N__9133;
    wire N__9130;
    wire N__9127;
    wire N__9124;
    wire N__9121;
    wire N__9118;
    wire N__9115;
    wire N__9112;
    wire N__9109;
    wire N__9106;
    wire N__9103;
    wire N__9100;
    wire N__9097;
    wire N__9094;
    wire N__9091;
    wire N__9088;
    wire N__9085;
    wire N__9082;
    wire N__9079;
    wire N__9076;
    wire N__9073;
    wire N__9070;
    wire N__9067;
    wire N__9064;
    wire N__9061;
    wire N__9058;
    wire N__9055;
    wire N__9052;
    wire N__9049;
    wire N__9046;
    wire N__9043;
    wire N__9040;
    wire N__9037;
    wire N__9034;
    wire N__9031;
    wire N__9028;
    wire N__9025;
    wire N__9022;
    wire N__9019;
    wire N__9016;
    wire N__9013;
    wire N__9010;
    wire N__9009;
    wire N__9006;
    wire N__9003;
    wire N__8998;
    wire N__8997;
    wire N__8994;
    wire N__8991;
    wire N__8990;
    wire N__8985;
    wire N__8982;
    wire N__8979;
    wire N__8976;
    wire N__8975;
    wire N__8974;
    wire N__8969;
    wire N__8966;
    wire N__8963;
    wire N__8958;
    wire N__8955;
    wire N__8954;
    wire N__8951;
    wire N__8948;
    wire N__8945;
    wire N__8942;
    wire N__8941;
    wire N__8938;
    wire N__8935;
    wire N__8932;
    wire N__8929;
    wire N__8924;
    wire N__8919;
    wire N__8916;
    wire N__8913;
    wire N__8910;
    wire N__8907;
    wire N__8902;
    wire N__8899;
    wire N__8896;
    wire N__8893;
    wire N__8890;
    wire N__8887;
    wire N__8884;
    wire N__8883;
    wire N__8880;
    wire N__8877;
    wire N__8876;
    wire N__8875;
    wire N__8870;
    wire N__8867;
    wire N__8864;
    wire N__8857;
    wire N__8856;
    wire N__8855;
    wire N__8852;
    wire N__8849;
    wire N__8846;
    wire N__8841;
    wire N__8840;
    wire N__8839;
    wire N__8836;
    wire N__8833;
    wire N__8830;
    wire N__8827;
    wire N__8824;
    wire N__8821;
    wire N__8818;
    wire N__8815;
    wire N__8812;
    wire N__8809;
    wire N__8806;
    wire N__8803;
    wire N__8800;
    wire N__8797;
    wire N__8794;
    wire N__8791;
    wire N__8788;
    wire N__8783;
    wire N__8780;
    wire N__8773;
    wire N__8772;
    wire N__8769;
    wire N__8766;
    wire N__8765;
    wire N__8760;
    wire N__8757;
    wire N__8752;
    wire N__8751;
    wire N__8750;
    wire N__8747;
    wire N__8744;
    wire N__8743;
    wire N__8740;
    wire N__8735;
    wire N__8732;
    wire N__8729;
    wire N__8726;
    wire N__8723;
    wire N__8722;
    wire N__8719;
    wire N__8716;
    wire N__8713;
    wire N__8710;
    wire N__8707;
    wire N__8704;
    wire N__8701;
    wire N__8698;
    wire N__8697;
    wire N__8694;
    wire N__8691;
    wire N__8688;
    wire N__8685;
    wire N__8682;
    wire N__8671;
    wire N__8668;
    wire N__8667;
    wire N__8666;
    wire N__8665;
    wire N__8662;
    wire N__8659;
    wire N__8656;
    wire N__8653;
    wire N__8650;
    wire N__8649;
    wire N__8646;
    wire N__8643;
    wire N__8642;
    wire N__8639;
    wire N__8636;
    wire N__8633;
    wire N__8630;
    wire N__8627;
    wire N__8626;
    wire N__8625;
    wire N__8622;
    wire N__8619;
    wire N__8616;
    wire N__8613;
    wire N__8610;
    wire N__8607;
    wire N__8604;
    wire N__8601;
    wire N__8598;
    wire N__8595;
    wire N__8588;
    wire N__8583;
    wire N__8580;
    wire N__8577;
    wire N__8574;
    wire N__8567;
    wire N__8564;
    wire N__8557;
    wire N__8556;
    wire N__8553;
    wire N__8550;
    wire N__8547;
    wire N__8546;
    wire N__8543;
    wire N__8540;
    wire N__8537;
    wire N__8536;
    wire N__8533;
    wire N__8528;
    wire N__8525;
    wire N__8522;
    wire N__8521;
    wire N__8516;
    wire N__8515;
    wire N__8512;
    wire N__8509;
    wire N__8508;
    wire N__8505;
    wire N__8502;
    wire N__8497;
    wire N__8494;
    wire N__8489;
    wire N__8484;
    wire N__8483;
    wire N__8480;
    wire N__8477;
    wire N__8474;
    wire N__8471;
    wire N__8466;
    wire N__8463;
    wire N__8460;
    wire N__8455;
    wire N__8452;
    wire N__8451;
    wire N__8448;
    wire N__8447;
    wire N__8444;
    wire N__8441;
    wire N__8440;
    wire N__8437;
    wire N__8434;
    wire N__8433;
    wire N__8430;
    wire N__8427;
    wire N__8424;
    wire N__8421;
    wire N__8418;
    wire N__8417;
    wire N__8412;
    wire N__8411;
    wire N__8408;
    wire N__8403;
    wire N__8400;
    wire N__8397;
    wire N__8394;
    wire N__8391;
    wire N__8386;
    wire N__8381;
    wire N__8380;
    wire N__8377;
    wire N__8374;
    wire N__8371;
    wire N__8368;
    wire N__8363;
    wire N__8358;
    wire N__8355;
    wire N__8352;
    wire N__8347;
    wire N__8346;
    wire N__8343;
    wire N__8340;
    wire N__8337;
    wire N__8336;
    wire N__8335;
    wire N__8332;
    wire N__8329;
    wire N__8326;
    wire N__8325;
    wire N__8322;
    wire N__8321;
    wire N__8318;
    wire N__8313;
    wire N__8310;
    wire N__8307;
    wire N__8304;
    wire N__8301;
    wire N__8296;
    wire N__8293;
    wire N__8290;
    wire N__8289;
    wire N__8286;
    wire N__8283;
    wire N__8280;
    wire N__8277;
    wire N__8274;
    wire N__8271;
    wire N__8268;
    wire N__8265;
    wire N__8262;
    wire N__8259;
    wire N__8258;
    wire N__8255;
    wire N__8252;
    wire N__8245;
    wire N__8242;
    wire N__8237;
    wire N__8234;
    wire N__8231;
    wire N__8228;
    wire N__8225;
    wire N__8222;
    wire N__8215;
    wire N__8214;
    wire N__8211;
    wire N__8208;
    wire N__8207;
    wire N__8206;
    wire N__8203;
    wire N__8200;
    wire N__8197;
    wire N__8194;
    wire N__8193;
    wire N__8190;
    wire N__8187;
    wire N__8184;
    wire N__8183;
    wire N__8182;
    wire N__8179;
    wire N__8176;
    wire N__8175;
    wire N__8172;
    wire N__8169;
    wire N__8166;
    wire N__8163;
    wire N__8160;
    wire N__8157;
    wire N__8154;
    wire N__8151;
    wire N__8146;
    wire N__8143;
    wire N__8140;
    wire N__8137;
    wire N__8130;
    wire N__8125;
    wire N__8122;
    wire N__8119;
    wire N__8116;
    wire N__8109;
    wire TVP_VIDEO_c_3;
    wire VCCG0;
    wire TVP_VIDEO_c_5;
    wire TVP_VIDEO_c_4;
    wire GNDG0;
    wire TVP_VIDEO_c_7;
    wire TVP_VIDEO_c_6;
    wire TVP_VIDEO_c_8;
    wire TVP_VIDEO_c_9;
    wire TVP_VIDEO_c_2;
    wire \receive_module.rx_counter.n12_cascade_ ;
    wire \receive_module.rx_counter.n3938_cascade_ ;
    wire \receive_module.rx_counter.n3938 ;
    wire \receive_module.rx_counter.n13 ;
    wire \receive_module.rx_counter.n3176_cascade_ ;
    wire \receive_module.rx_counter.n3208 ;
    wire \line_buffer.n675 ;
    wire \line_buffer.n683 ;
    wire \line_buffer.n611 ;
    wire \line_buffer.n4170_cascade_ ;
    wire \line_buffer.n619 ;
    wire \line_buffer.n643 ;
    wire \line_buffer.n651 ;
    wire \line_buffer.n687 ;
    wire \line_buffer.n679 ;
    wire \line_buffer.n4152 ;
    wire \line_buffer.n554 ;
    wire \line_buffer.n546 ;
    wire \line_buffer.n4155_cascade_ ;
    wire \line_buffer.n4173 ;
    wire \transmit_module.Y_DELTA_PATTERN_95 ;
    wire \line_buffer.n680 ;
    wire \line_buffer.n688 ;
    wire bfn_10_9_0_;
    wire \receive_module.rx_counter.n3669 ;
    wire \receive_module.rx_counter.n3670 ;
    wire \receive_module.rx_counter.n3671 ;
    wire \receive_module.rx_counter.n3672 ;
    wire \receive_module.rx_counter.n3673 ;
    wire \receive_module.rx_counter.n3674 ;
    wire \receive_module.rx_counter.n3675 ;
    wire \receive_module.rx_counter.n3676 ;
    wire bfn_10_10_0_;
    wire \transmit_module.Y_DELTA_PATTERN_84 ;
    wire \transmit_module.Y_DELTA_PATTERN_83 ;
    wire \transmit_module.Y_DELTA_PATTERN_90 ;
    wire \transmit_module.Y_DELTA_PATTERN_89 ;
    wire \transmit_module.Y_DELTA_PATTERN_88 ;
    wire \transmit_module.Y_DELTA_PATTERN_87 ;
    wire \transmit_module.Y_DELTA_PATTERN_92 ;
    wire \transmit_module.Y_DELTA_PATTERN_91 ;
    wire \transmit_module.Y_DELTA_PATTERN_86 ;
    wire \transmit_module.Y_DELTA_PATTERN_85 ;
    wire \transmit_module.Y_DELTA_PATTERN_94 ;
    wire \transmit_module.Y_DELTA_PATTERN_93 ;
    wire \transmit_module.Y_DELTA_PATTERN_96 ;
    wire \transmit_module.Y_DELTA_PATTERN_97 ;
    wire \line_buffer.n624 ;
    wire \line_buffer.n4122 ;
    wire \line_buffer.n616 ;
    wire \receive_module.rx_counter.Y_0 ;
    wire bfn_11_9_0_;
    wire \receive_module.rx_counter.Y_1 ;
    wire \receive_module.rx_counter.n3711 ;
    wire \receive_module.rx_counter.Y_2 ;
    wire \receive_module.rx_counter.n3712 ;
    wire \receive_module.rx_counter.Y_3 ;
    wire \receive_module.rx_counter.n3713 ;
    wire \receive_module.rx_counter.Y_4 ;
    wire \receive_module.rx_counter.n3714 ;
    wire \receive_module.rx_counter.Y_5 ;
    wire \receive_module.rx_counter.n3715 ;
    wire \receive_module.rx_counter.Y_6 ;
    wire \receive_module.rx_counter.n3716 ;
    wire \receive_module.rx_counter.Y_7 ;
    wire \receive_module.rx_counter.n3717 ;
    wire \receive_module.rx_counter.n3718 ;
    wire \receive_module.rx_counter.Y_8 ;
    wire bfn_11_10_0_;
    wire \receive_module.rx_counter.n3979 ;
    wire \receive_module.rx_counter.O_VISIBLE_N_89 ;
    wire DEBUG_c_6;
    wire \transmit_module.video_signal_controller.SYNC_BUFF1 ;
    wire \transmit_module.video_signal_controller.n3987_cascade_ ;
    wire \transmit_module.video_signal_controller.n4_cascade_ ;
    wire \transmit_module.video_signal_controller.n3935 ;
    wire \transmit_module.video_signal_controller.n3935_cascade_ ;
    wire \transmit_module.video_signal_controller.n6 ;
    wire \transmit_module.Y_DELTA_PATTERN_98 ;
    wire \transmit_module.Y_DELTA_PATTERN_76 ;
    wire \transmit_module.Y_DELTA_PATTERN_73 ;
    wire \transmit_module.Y_DELTA_PATTERN_82 ;
    wire \transmit_module.Y_DELTA_PATTERN_75 ;
    wire \transmit_module.Y_DELTA_PATTERN_74 ;
    wire \transmit_module.Y_DELTA_PATTERN_77 ;
    wire n1996;
    wire INVADV_R__i1C_net;
    wire \transmit_module.Y_DELTA_PATTERN_70 ;
    wire \transmit_module.Y_DELTA_PATTERN_72 ;
    wire \transmit_module.Y_DELTA_PATTERN_71 ;
    wire \transmit_module.Y_DELTA_PATTERN_63 ;
    wire n18;
    wire \receive_module.rx_counter.PULSE_1HZ_N_97 ;
    wire \receive_module.n4212_cascade_ ;
    wire \receive_module.n4213_cascade_ ;
    wire \receive_module.rx_counter.n3204 ;
    wire n659;
    wire DEBUG_c_0;
    wire n691;
    wire \line_buffer.n626 ;
    wire \line_buffer.n561 ;
    wire \transmit_module.video_signal_controller.n3978_cascade_ ;
    wire \transmit_module.video_signal_controller.n4052 ;
    wire \transmit_module.video_signal_controller.n4216_cascade_ ;
    wire \transmit_module.video_signal_controller.n12 ;
    wire \transmit_module.video_signal_controller.n2274_cascade_ ;
    wire \transmit_module.video_signal_controller.SYNC_BUFF2 ;
    wire \transmit_module.video_signal_controller.n3226 ;
    wire \transmit_module.video_signal_controller.n2260 ;
    wire \transmit_module.video_signal_controller.n3917 ;
    wire \transmit_module.video_signal_controller.n2260_cascade_ ;
    wire \transmit_module.video_signal_controller.n4217 ;
    wire \transmit_module.video_signal_controller.n18_cascade_ ;
    wire \transmit_module.video_signal_controller.n2219 ;
    wire \transmit_module.video_signal_controller.VGA_Y_0 ;
    wire bfn_12_16_0_;
    wire \transmit_module.video_signal_controller.VGA_Y_1 ;
    wire \transmit_module.video_signal_controller.n3677 ;
    wire \transmit_module.video_signal_controller.VGA_Y_2 ;
    wire \transmit_module.video_signal_controller.n3678 ;
    wire \transmit_module.video_signal_controller.n3679 ;
    wire \transmit_module.video_signal_controller.n3680 ;
    wire \transmit_module.video_signal_controller.VGA_Y_5 ;
    wire \transmit_module.video_signal_controller.n3681 ;
    wire \transmit_module.video_signal_controller.VGA_Y_6 ;
    wire \transmit_module.video_signal_controller.n3682 ;
    wire \transmit_module.video_signal_controller.VGA_Y_7 ;
    wire \transmit_module.video_signal_controller.n3683 ;
    wire \transmit_module.video_signal_controller.n3684 ;
    wire \transmit_module.video_signal_controller.VGA_Y_8 ;
    wire bfn_12_17_0_;
    wire \transmit_module.video_signal_controller.n3685 ;
    wire \transmit_module.video_signal_controller.n3686 ;
    wire \transmit_module.video_signal_controller.n3687 ;
    wire \transmit_module.video_signal_controller.n2594 ;
    wire \transmit_module.video_signal_controller.VGA_Y_3 ;
    wire \transmit_module.video_signal_controller.n4215 ;
    wire \transmit_module.video_signal_controller.VGA_Y_4 ;
    wire \transmit_module.video_signal_controller.n3892 ;
    wire \transmit_module.video_signal_controller.VGA_Y_9 ;
    wire \transmit_module.video_signal_controller.VGA_VISIBLE_Y_N_553_cascade_ ;
    wire \transmit_module.video_signal_controller.n3936 ;
    wire \transmit_module.n3926_cascade_ ;
    wire \transmit_module.video_signal_controller.VGA_Y_11 ;
    wire \transmit_module.video_signal_controller.VGA_Y_10 ;
    wire \transmit_module.video_signal_controller.n4218 ;
    wire \transmit_module.n219_cascade_ ;
    wire n28;
    wire n4210;
    wire n4210_cascade_;
    wire \transmit_module.Y_DELTA_PATTERN_64 ;
    wire \transmit_module.Y_DELTA_PATTERN_67 ;
    wire \transmit_module.Y_DELTA_PATTERN_81 ;
    wire \transmit_module.Y_DELTA_PATTERN_69 ;
    wire \transmit_module.Y_DELTA_PATTERN_68 ;
    wire \transmit_module.Y_DELTA_PATTERN_78 ;
    wire \transmit_module.Y_DELTA_PATTERN_62 ;
    wire \transmit_module.Y_DELTA_PATTERN_66 ;
    wire \transmit_module.Y_DELTA_PATTERN_65 ;
    wire \transmit_module.Y_DELTA_PATTERN_80 ;
    wire \transmit_module.Y_DELTA_PATTERN_79 ;
    wire \transmit_module.Y_DELTA_PATTERN_57 ;
    wire \transmit_module.ADDR_Y_COMPONENT_10 ;
    wire \transmit_module.n209 ;
    wire \transmit_module.n178 ;
    wire \transmit_module.n209_cascade_ ;
    wire n2283;
    wire old_HS;
    wire RX_ADDR_3;
    wire bfn_13_10_0_;
    wire RX_ADDR_4;
    wire \receive_module.rx_counter.n3650 ;
    wire RX_ADDR_5;
    wire \receive_module.rx_counter.n3651 ;
    wire \receive_module.rx_counter.n3652 ;
    wire \receive_module.rx_counter.n3653 ;
    wire \receive_module.rx_counter.n3654 ;
    wire \receive_module.rx_counter.n3655 ;
    wire \receive_module.O_X_9 ;
    wire \receive_module.rx_counter.n4 ;
    wire \receive_module.O_Y_0 ;
    wire \receive_module.O_X_6 ;
    wire RX_ADDR_6;
    wire bfn_13_11_0_;
    wire \receive_module.O_X_7 ;
    wire \receive_module.O_Y_1 ;
    wire RX_ADDR_7;
    wire \receive_module.n3699 ;
    wire \receive_module.O_Y_2 ;
    wire \receive_module.O_X_8 ;
    wire RX_ADDR_8;
    wire \receive_module.n3700 ;
    wire \receive_module.n7 ;
    wire \receive_module.O_Y_3 ;
    wire RX_ADDR_9;
    wire \receive_module.n3701 ;
    wire \receive_module.n6 ;
    wire \receive_module.O_Y_4 ;
    wire RX_ADDR_10;
    wire \receive_module.n3702 ;
    wire \receive_module.n5 ;
    wire \receive_module.O_Y_5 ;
    wire \receive_module.n3703 ;
    wire \receive_module.n4 ;
    wire \receive_module.O_Y_6 ;
    wire \receive_module.n3704 ;
    wire \receive_module.n3 ;
    wire \receive_module.O_Y_7 ;
    wire \receive_module.n3705 ;
    wire \line_buffer.n627 ;
    wire \line_buffer.n562 ;
    wire n690;
    wire \db5.COUNTER_3 ;
    wire \db5.NEXT_COUNTER_3 ;
    wire \db5.COUNTER_2 ;
    wire \db5.NEXT_COUNTER_2 ;
    wire \db5.COUNTER_1 ;
    wire \db5.NEXT_COUNTER_1 ;
    wire \db5.COUNTER_0 ;
    wire \db5.NEXT_COUNTER_0 ;
    wire \INVdb5.NEXT_COUNTER__i3C_net ;
    wire \db5.n4221 ;
    wire \transmit_module.video_signal_controller.n3997 ;
    wire \transmit_module.video_signal_controller.n3196 ;
    wire \line_buffer.n655 ;
    wire \line_buffer.n647 ;
    wire \transmit_module.video_signal_controller.VGA_X_0 ;
    wire bfn_13_15_0_;
    wire \transmit_module.video_signal_controller.VGA_X_1 ;
    wire \transmit_module.video_signal_controller.n3688 ;
    wire \transmit_module.video_signal_controller.VGA_X_2 ;
    wire \transmit_module.video_signal_controller.n3689 ;
    wire \transmit_module.video_signal_controller.VGA_X_3 ;
    wire \transmit_module.video_signal_controller.n3690 ;
    wire \transmit_module.video_signal_controller.VGA_X_4 ;
    wire \transmit_module.video_signal_controller.n3691 ;
    wire \transmit_module.video_signal_controller.VGA_X_5 ;
    wire \transmit_module.video_signal_controller.n3692 ;
    wire \transmit_module.video_signal_controller.VGA_X_6 ;
    wire \transmit_module.video_signal_controller.n3693 ;
    wire \transmit_module.video_signal_controller.VGA_X_7 ;
    wire \transmit_module.video_signal_controller.n3694 ;
    wire \transmit_module.video_signal_controller.n3695 ;
    wire \transmit_module.video_signal_controller.VGA_X_8 ;
    wire bfn_13_16_0_;
    wire \transmit_module.video_signal_controller.VGA_X_9 ;
    wire \transmit_module.video_signal_controller.n3696 ;
    wire \transmit_module.video_signal_controller.VGA_X_10 ;
    wire \transmit_module.video_signal_controller.n3697 ;
    wire \transmit_module.video_signal_controller.n3698 ;
    wire \transmit_module.video_signal_controller.VGA_X_11 ;
    wire \transmit_module.video_signal_controller.n2274 ;
    wire \line_buffer.n4102 ;
    wire \line_buffer.n648 ;
    wire \line_buffer.n656 ;
    wire \transmit_module.n186 ;
    wire \transmit_module.n4211_cascade_ ;
    wire \transmit_module.n217 ;
    wire n26;
    wire \line_buffer.n559 ;
    wire \line_buffer.n4182 ;
    wire \line_buffer.n551 ;
    wire \line_buffer.n4185_cascade_ ;
    wire \line_buffer.n4125 ;
    wire n1995;
    wire TX_DATA_2;
    wire n1994;
    wire n1993;
    wire n1992;
    wire n1991;
    wire TX_DATA_6;
    wire n1990;
    wire TX_DATA_7;
    wire ADV_B_c;
    wire INVADV_R__i2C_net;
    wire n2587;
    wire \transmit_module.Y_DELTA_PATTERN_43 ;
    wire \transmit_module.Y_DELTA_PATTERN_44 ;
    wire \transmit_module.Y_DELTA_PATTERN_46 ;
    wire \transmit_module.Y_DELTA_PATTERN_45 ;
    wire \transmit_module.Y_DELTA_PATTERN_47 ;
    wire \transmit_module.Y_DELTA_PATTERN_48 ;
    wire \transmit_module.Y_DELTA_PATTERN_53 ;
    wire \transmit_module.Y_DELTA_PATTERN_52 ;
    wire \transmit_module.Y_DELTA_PATTERN_49 ;
    wire \transmit_module.Y_DELTA_PATTERN_54 ;
    wire \transmit_module.Y_DELTA_PATTERN_51 ;
    wire \transmit_module.Y_DELTA_PATTERN_50 ;
    wire \transmit_module.Y_DELTA_PATTERN_56 ;
    wire \transmit_module.Y_DELTA_PATTERN_55 ;
    wire \transmit_module.Y_DELTA_PATTERN_59 ;
    wire \transmit_module.Y_DELTA_PATTERN_58 ;
    wire \transmit_module.Y_DELTA_PATTERN_61 ;
    wire \transmit_module.Y_DELTA_PATTERN_60 ;
    wire \line_buffer.n558 ;
    wire \line_buffer.n550 ;
    wire \line_buffer.n4101 ;
    wire n22;
    wire \receive_module.rx_counter.n5_cascade_ ;
    wire TVP_HSYNC_c;
    wire \receive_module.rx_counter.n4_adj_576 ;
    wire RX_ADDR_0;
    wire bfn_14_9_0_;
    wire RX_ADDR_1;
    wire \receive_module.rx_counter.n3720 ;
    wire RX_ADDR_2;
    wire \receive_module.rx_counter.n3721 ;
    wire \receive_module.rx_counter.n3722 ;
    wire \receive_module.rx_counter.n3723 ;
    wire \receive_module.rx_counter.n3724 ;
    wire \receive_module.rx_counter.n3725 ;
    wire \receive_module.rx_counter.n3726 ;
    wire \receive_module.rx_counter.n3727 ;
    wire bfn_14_10_0_;
    wire \receive_module.rx_counter.n3728 ;
    wire n4214;
    wire RX_ADDR_11;
    wire RX_ADDR_12;
    wire DEBUG_c_5;
    wire DEBUG_c_3;
    wire n658;
    wire \transmit_module.X_DELTA_PATTERN_13 ;
    wire \transmit_module.X_DELTA_PATTERN_9 ;
    wire \transmit_module.X_DELTA_PATTERN_12 ;
    wire \transmit_module.X_DELTA_PATTERN_11 ;
    wire \transmit_module.X_DELTA_PATTERN_10 ;
    wire \line_buffer.n4072 ;
    wire \line_buffer.n4134 ;
    wire \transmit_module.n2361 ;
    wire \transmit_module.ADDR_Y_COMPONENT_2 ;
    wire \transmit_module.n219 ;
    wire \transmit_module.n179_cascade_ ;
    wire \transmit_module.n213 ;
    wire \transmit_module.n179 ;
    wire \transmit_module.n210 ;
    wire n19;
    wire \transmit_module.n180 ;
    wire \transmit_module.n211 ;
    wire n20;
    wire \transmit_module.old_VGA_HS ;
    wire ADV_HSYNC_c;
    wire \transmit_module.n181 ;
    wire \transmit_module.n212 ;
    wire \transmit_module.n181_cascade_ ;
    wire n21;
    wire \transmit_module.ADDR_Y_COMPONENT_7 ;
    wire \transmit_module.ADDR_Y_COMPONENT_6 ;
    wire \transmit_module.n182 ;
    wire \receive_module.rx_counter.FRAME_COUNTER_0 ;
    wire bfn_15_8_0_;
    wire \receive_module.rx_counter.FRAME_COUNTER_1 ;
    wire \receive_module.rx_counter.n3706 ;
    wire \receive_module.rx_counter.FRAME_COUNTER_2 ;
    wire \receive_module.rx_counter.n3707 ;
    wire \receive_module.rx_counter.FRAME_COUNTER_3 ;
    wire \receive_module.rx_counter.n3708 ;
    wire \receive_module.rx_counter.FRAME_COUNTER_4 ;
    wire \receive_module.rx_counter.n3709 ;
    wire \receive_module.rx_counter.n3710 ;
    wire \receive_module.rx_counter.FRAME_COUNTER_5 ;
    wire \receive_module.rx_counter.n2605 ;
    wire \receive_module.rx_counter.old_VS ;
    wire TVP_VSYNC_c;
    wire \receive_module.rx_counter.X_5 ;
    wire \receive_module.rx_counter.X_4 ;
    wire \receive_module.rx_counter.X_3 ;
    wire \receive_module.rx_counter.X_8 ;
    wire \receive_module.rx_counter.X_9 ;
    wire \receive_module.rx_counter.n4219 ;
    wire \receive_module.rx_counter.X_7 ;
    wire \receive_module.rx_counter.n4_adj_575_cascade_ ;
    wire \receive_module.rx_counter.X_6 ;
    wire \receive_module.rx_counter.O_VISIBLE_N_86 ;
    wire \receive_module.rx_counter.n11 ;
    wire LED_c;
    wire \receive_module.rx_counter.n4222 ;
    wire \line_buffer.n623 ;
    wire \line_buffer.n615 ;
    wire \line_buffer.n4071 ;
    wire \line_buffer.n646 ;
    wire \line_buffer.n654 ;
    wire \line_buffer.n549 ;
    wire \line_buffer.n4176_cascade_ ;
    wire \line_buffer.n557 ;
    wire \transmit_module.X_DELTA_PATTERN_8 ;
    wire \transmit_module.X_DELTA_PATTERN_7 ;
    wire \transmit_module.X_DELTA_PATTERN_6 ;
    wire \transmit_module.X_DELTA_PATTERN_14 ;
    wire \transmit_module.X_DELTA_PATTERN_2 ;
    wire \transmit_module.X_DELTA_PATTERN_1 ;
    wire \transmit_module.X_DELTA_PATTERN_3 ;
    wire \transmit_module.X_DELTA_PATTERN_15 ;
    wire \transmit_module.X_DELTA_PATTERN_5 ;
    wire \transmit_module.X_DELTA_PATTERN_4 ;
    wire \transmit_module.n2315 ;
    wire \transmit_module.X_DELTA_PATTERN_0 ;
    wire \transmit_module.n204 ;
    wire bfn_15_17_0_;
    wire \transmit_module.n3656 ;
    wire \transmit_module.TX_ADDR_2 ;
    wire \transmit_module.n202 ;
    wire \transmit_module.n3657 ;
    wire \transmit_module.n201 ;
    wire \transmit_module.n3658 ;
    wire \transmit_module.n3659 ;
    wire \transmit_module.n3660 ;
    wire \transmit_module.TX_ADDR_6 ;
    wire \transmit_module.n198 ;
    wire \transmit_module.n3661 ;
    wire \transmit_module.TX_ADDR_7 ;
    wire \transmit_module.n197 ;
    wire \transmit_module.n3662 ;
    wire \transmit_module.n3663 ;
    wire \transmit_module.n196 ;
    wire bfn_15_18_0_;
    wire \transmit_module.n195 ;
    wire \transmit_module.n3664 ;
    wire \transmit_module.TX_ADDR_10 ;
    wire \transmit_module.n194 ;
    wire \transmit_module.n3665 ;
    wire \transmit_module.n3666 ;
    wire \transmit_module.n3667 ;
    wire \transmit_module.n3668 ;
    wire \transmit_module.TX_ADDR_8 ;
    wire \transmit_module.ADDR_Y_COMPONENT_8 ;
    wire \transmit_module.n203 ;
    wire \transmit_module.n218_cascade_ ;
    wire \transmit_module.n188 ;
    wire \transmit_module.TX_ADDR_0 ;
    wire \transmit_module.ADDR_Y_COMPONENT_0 ;
    wire \transmit_module.TX_ADDR_3 ;
    wire \transmit_module.ADDR_Y_COMPONENT_3 ;
    wire \transmit_module.n193 ;
    wire \transmit_module.ADDR_Y_COMPONENT_11 ;
    wire \transmit_module.ADDR_Y_COMPONENT_1 ;
    wire \transmit_module.TX_ADDR_1 ;
    wire \transmit_module.n187 ;
    wire \transmit_module.n218 ;
    wire n27;
    wire \line_buffer.n678 ;
    wire \line_buffer.n686 ;
    wire \line_buffer.n614 ;
    wire \line_buffer.n4188_cascade_ ;
    wire \line_buffer.n622 ;
    wire \line_buffer.n4191_cascade_ ;
    wire \line_buffer.n4179 ;
    wire TX_DATA_5;
    wire \transmit_module.Y_DELTA_PATTERN_18 ;
    wire \transmit_module.Y_DELTA_PATTERN_21 ;
    wire \transmit_module.Y_DELTA_PATTERN_20 ;
    wire \transmit_module.Y_DELTA_PATTERN_19 ;
    wire \transmit_module.Y_DELTA_PATTERN_1 ;
    wire \transmit_module.TX_ADDR_9 ;
    wire \transmit_module.ADDR_Y_COMPONENT_9 ;
    wire \transmit_module.n200 ;
    wire \transmit_module.n215_cascade_ ;
    wire \transmit_module.ADDR_Y_COMPONENT_5 ;
    wire \transmit_module.n191 ;
    wire \transmit_module.BRAM_ADDR_13_N_258_13 ;
    wire \transmit_module.n199 ;
    wire \transmit_module.n3910 ;
    wire \transmit_module.n214_cascade_ ;
    wire \transmit_module.TX_ADDR_5 ;
    wire \transmit_module.ADDR_Y_COMPONENT_4 ;
    wire \transmit_module.TX_ADDR_4 ;
    wire \transmit_module.n184 ;
    wire \transmit_module.n215 ;
    wire n24;
    wire \transmit_module.n183 ;
    wire \transmit_module.n214 ;
    wire n23;
    wire \transmit_module.n4220 ;
    wire \transmit_module.n192 ;
    wire \transmit_module.n3926 ;
    wire \transmit_module.n2277 ;
    wire \transmit_module.Y_DELTA_PATTERN_42 ;
    wire DEBUG_c_1_c;
    wire GB_BUFFER_DEBUG_c_1_c_THRU_CO;
    wire \transmit_module.Y_DELTA_PATTERN_29 ;
    wire \transmit_module.Y_DELTA_PATTERN_31 ;
    wire \transmit_module.Y_DELTA_PATTERN_30 ;
    wire \transmit_module.Y_DELTA_PATTERN_12 ;
    wire \transmit_module.Y_DELTA_PATTERN_32 ;
    wire \transmit_module.Y_DELTA_PATTERN_13 ;
    wire \transmit_module.Y_DELTA_PATTERN_14 ;
    wire \transmit_module.Y_DELTA_PATTERN_26 ;
    wire \transmit_module.Y_DELTA_PATTERN_25 ;
    wire \transmit_module.Y_DELTA_PATTERN_28 ;
    wire \transmit_module.Y_DELTA_PATTERN_27 ;
    wire \transmit_module.Y_DELTA_PATTERN_0 ;
    wire \transmit_module.Y_DELTA_PATTERN_99 ;
    wire \transmit_module.Y_DELTA_PATTERN_37 ;
    wire \transmit_module.Y_DELTA_PATTERN_36 ;
    wire \transmit_module.Y_DELTA_PATTERN_38 ;
    wire \transmit_module.n185 ;
    wire \transmit_module.n216 ;
    wire \transmit_module.n4211 ;
    wire n25;
    wire \transmit_module.ADDR_Y_COMPONENT_12 ;
    wire \transmit_module.ADDR_Y_COMPONENT_13 ;
    wire \transmit_module.n2305 ;
    wire \transmit_module.Y_DELTA_PATTERN_39 ;
    wire \transmit_module.Y_DELTA_PATTERN_41 ;
    wire \transmit_module.Y_DELTA_PATTERN_40 ;
    wire \line_buffer.n620 ;
    wire \line_buffer.n612 ;
    wire \transmit_module.Y_DELTA_PATTERN_6 ;
    wire \transmit_module.Y_DELTA_PATTERN_5 ;
    wire \transmit_module.Y_DELTA_PATTERN_7 ;
    wire \transmit_module.Y_DELTA_PATTERN_11 ;
    wire \transmit_module.Y_DELTA_PATTERN_10 ;
    wire \transmit_module.Y_DELTA_PATTERN_9 ;
    wire \transmit_module.Y_DELTA_PATTERN_8 ;
    wire \transmit_module.Y_DELTA_PATTERN_15 ;
    wire \transmit_module.Y_DELTA_PATTERN_4 ;
    wire \transmit_module.Y_DELTA_PATTERN_17 ;
    wire \transmit_module.Y_DELTA_PATTERN_16 ;
    wire \transmit_module.Y_DELTA_PATTERN_3 ;
    wire \transmit_module.Y_DELTA_PATTERN_2 ;
    wire \transmit_module.Y_DELTA_PATTERN_22 ;
    wire \transmit_module.Y_DELTA_PATTERN_24 ;
    wire \transmit_module.Y_DELTA_PATTERN_23 ;
    wire \transmit_module.n4224 ;
    wire \line_buffer.n642 ;
    wire \line_buffer.n650 ;
    wire \line_buffer.n545 ;
    wire \line_buffer.n4164_cascade_ ;
    wire \line_buffer.n553 ;
    wire \line_buffer.n4167_cascade_ ;
    wire TX_DATA_1;
    wire \line_buffer.n4065 ;
    wire \line_buffer.n684 ;
    wire \line_buffer.n676 ;
    wire \line_buffer.n4066 ;
    wire \line_buffer.n555 ;
    wire \line_buffer.n547 ;
    wire \line_buffer.n4074_cascade_ ;
    wire \line_buffer.n4128 ;
    wire TX_DATA_3;
    wire \line_buffer.n652 ;
    wire \line_buffer.n644 ;
    wire \line_buffer.n4075 ;
    wire \transmit_module.Y_DELTA_PATTERN_33 ;
    wire \transmit_module.Y_DELTA_PATTERN_35 ;
    wire \transmit_module.Y_DELTA_PATTERN_34 ;
    wire \transmit_module.n4225 ;
    wire ADV_VSYNC_c;
    wire \line_buffer.n617 ;
    wire \line_buffer.n609 ;
    wire \line_buffer.n610 ;
    wire \line_buffer.n618 ;
    wire \line_buffer.n4161 ;
    wire \line_buffer.n673 ;
    wire \line_buffer.n681 ;
    wire \line_buffer.n4146 ;
    wire \line_buffer.n4149 ;
    wire TX_DATA_0;
    wire \line_buffer.n621 ;
    wire \line_buffer.n613 ;
    wire \line_buffer.n653 ;
    wire \line_buffer.n645 ;
    wire \line_buffer.n4062 ;
    wire \line_buffer.n4078 ;
    wire DEBUG_c_2;
    wire \line_buffer.n4140 ;
    wire TX_DATA_4;
    wire ADV_CLK_c;
    wire \line_buffer.n641 ;
    wire \line_buffer.n649 ;
    wire \line_buffer.n552 ;
    wire \line_buffer.n4116 ;
    wire \line_buffer.n544 ;
    wire \line_buffer.n4119 ;
    wire \line_buffer.n548 ;
    wire \line_buffer.n556 ;
    wire \line_buffer.n4077 ;
    wire \line_buffer.n674 ;
    wire TX_ADDR_12;
    wire \line_buffer.n682 ;
    wire \line_buffer.n4158 ;
    wire \line_buffer.n685 ;
    wire \line_buffer.n677 ;
    wire TX_ADDR_11;
    wire \line_buffer.n4063 ;
    wire CONSTANT_ONE_NET;
    wire _gnd_net_;

    defparam \tx_pll.TX_PLL_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \tx_pll.TX_PLL_inst .TEST_MODE=1'b0;
    defparam \tx_pll.TX_PLL_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \tx_pll.TX_PLL_inst .PLLOUT_SELECT="GENCLK";
    defparam \tx_pll.TX_PLL_inst .FILTER_RANGE=3'b010;
    defparam \tx_pll.TX_PLL_inst .FEEDBACK_PATH="SIMPLE";
    defparam \tx_pll.TX_PLL_inst .FDA_RELATIVE=4'b0000;
    defparam \tx_pll.TX_PLL_inst .FDA_FEEDBACK=4'b0000;
    defparam \tx_pll.TX_PLL_inst .ENABLE_ICEGATE=1'b0;
    defparam \tx_pll.TX_PLL_inst .DIVR=4'b0000;
    defparam \tx_pll.TX_PLL_inst .DIVQ=3'b100;
    defparam \tx_pll.TX_PLL_inst .DIVF=7'b0100110;
    defparam \tx_pll.TX_PLL_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE \tx_pll.TX_PLL_inst  (
            .EXTFEEDBACK(),
            .LATCHINPUTVALUE(),
            .SCLK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(ADV_CLK_c),
            .REFERENCECLK(N__19215),
            .RESETB(N__23324),
            .BYPASS(GNDG0),
            .SDI(),
            .DYNAMICDELAY({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,dangling_wire_4,dangling_wire_5,dangling_wire_6,dangling_wire_7}),
            .PLLOUTGLOBAL());
    defparam \line_buffer.mem2_physical .WRITE_MODE=3;
    defparam \line_buffer.mem2_physical .READ_MODE=3;
    defparam \line_buffer.mem2_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem2_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem2_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem2_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem2_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem2_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem2_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem2_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem2_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem2_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem2_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem2_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem2_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem2_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem2_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem2_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem2_physical  (
            .RDATA({dangling_wire_8,dangling_wire_9,dangling_wire_10,dangling_wire_11,\line_buffer.n559 ,dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,\line_buffer.n558 ,dangling_wire_19,dangling_wire_20,dangling_wire_21}),
            .RADDR({N__9840,N__16167,N__16833,N__16497,N__15513,N__18567,N__18801,N__19971,N__13950,N__18126,N__10740}),
            .WADDR({N__12804,N__13062,N__11814,N__12072,N__12339,N__11067,N__11292,N__11526,N__14790,N__15021,N__15252}),
            .MASK({dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29,dangling_wire_30,dangling_wire_31,dangling_wire_32,dangling_wire_33,dangling_wire_34,dangling_wire_35,dangling_wire_36,dangling_wire_37}),
            .WDATA({dangling_wire_38,dangling_wire_39,dangling_wire_40,dangling_wire_41,N__8743,dangling_wire_42,dangling_wire_43,dangling_wire_44,dangling_wire_45,dangling_wire_46,dangling_wire_47,dangling_wire_48,N__8855,dangling_wire_49,dangling_wire_50,dangling_wire_51}),
            .RCLKE(),
            .RCLK(N__22387),
            .RE(N__23189),
            .WCLKE(),
            .WCLK(N__19361),
            .WE(N__12610));
    defparam \line_buffer.mem14_physical .WRITE_MODE=3;
    defparam \line_buffer.mem14_physical .READ_MODE=3;
    defparam \line_buffer.mem14_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem14_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem14_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem14_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem14_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem14_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem14_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem14_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem14_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem14_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem14_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem14_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem14_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem14_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem14_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem14_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem14_physical  (
            .RDATA({dangling_wire_52,dangling_wire_53,dangling_wire_54,dangling_wire_55,\line_buffer.n646 ,dangling_wire_56,dangling_wire_57,dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,\line_buffer.n645 ,dangling_wire_63,dangling_wire_64,dangling_wire_65}),
            .RADDR({N__9912,N__16239,N__16905,N__16569,N__15585,N__18639,N__18873,N__20043,N__14022,N__18198,N__10812}),
            .WADDR({N__12876,N__13134,N__11886,N__12144,N__12411,N__11139,N__11364,N__11598,N__14862,N__15093,N__15324}),
            .MASK({dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73,dangling_wire_74,dangling_wire_75,dangling_wire_76,dangling_wire_77,dangling_wire_78,dangling_wire_79,dangling_wire_80,dangling_wire_81}),
            .WDATA({dangling_wire_82,dangling_wire_83,dangling_wire_84,dangling_wire_85,N__8666,dangling_wire_86,dangling_wire_87,dangling_wire_88,dangling_wire_89,dangling_wire_90,dangling_wire_91,dangling_wire_92,N__8536,dangling_wire_93,dangling_wire_94,dangling_wire_95}),
            .RCLKE(),
            .RCLK(N__22623),
            .RE(N__23261),
            .WCLKE(),
            .WCLK(N__19346),
            .WE(N__15712));
    defparam \line_buffer.mem5_physical .WRITE_MODE=3;
    defparam \line_buffer.mem5_physical .READ_MODE=3;
    defparam \line_buffer.mem5_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem5_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem5_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem5_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem5_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem5_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem5_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem5_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem5_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem5_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem5_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem5_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem5_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem5_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem5_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem5_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem5_physical  (
            .RDATA({dangling_wire_96,dangling_wire_97,dangling_wire_98,dangling_wire_99,\line_buffer.n656 ,dangling_wire_100,dangling_wire_101,dangling_wire_102,dangling_wire_103,dangling_wire_104,dangling_wire_105,dangling_wire_106,\line_buffer.n655 ,dangling_wire_107,dangling_wire_108,dangling_wire_109}),
            .RADDR({N__9843,N__16176,N__16842,N__16506,N__15516,N__18582,N__18810,N__19986,N__13965,N__18129,N__10737}),
            .WADDR({N__12825,N__13077,N__11829,N__12081,N__12336,N__11076,N__11295,N__11523,N__14793,N__15030,N__15267}),
            .MASK({dangling_wire_110,dangling_wire_111,dangling_wire_112,dangling_wire_113,dangling_wire_114,dangling_wire_115,dangling_wire_116,dangling_wire_117,dangling_wire_118,dangling_wire_119,dangling_wire_120,dangling_wire_121,dangling_wire_122,dangling_wire_123,dangling_wire_124,dangling_wire_125}),
            .WDATA({dangling_wire_126,dangling_wire_127,dangling_wire_128,dangling_wire_129,N__8765,dangling_wire_130,dangling_wire_131,dangling_wire_132,dangling_wire_133,dangling_wire_134,dangling_wire_135,dangling_wire_136,N__8876,dangling_wire_137,dangling_wire_138,dangling_wire_139}),
            .RCLKE(),
            .RCLK(N__21959),
            .RE(N__23281),
            .WCLKE(),
            .WCLK(N__19360),
            .WE(N__10120));
    defparam \line_buffer.mem11_physical .WRITE_MODE=3;
    defparam \line_buffer.mem11_physical .READ_MODE=3;
    defparam \line_buffer.mem11_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem11_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem11_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem11_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem11_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem11_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem11_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem11_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem11_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem11_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem11_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem11_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem11_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem11_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem11_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem11_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem11_physical  (
            .RDATA({dangling_wire_140,dangling_wire_141,dangling_wire_142,dangling_wire_143,\line_buffer.n614 ,dangling_wire_144,dangling_wire_145,dangling_wire_146,dangling_wire_147,dangling_wire_148,dangling_wire_149,dangling_wire_150,\line_buffer.n613 ,dangling_wire_151,dangling_wire_152,dangling_wire_153}),
            .RADDR({N__9948,N__16275,N__16941,N__16605,N__15621,N__18675,N__18909,N__20079,N__14058,N__18234,N__10848}),
            .WADDR({N__12912,N__13170,N__11922,N__12180,N__12447,N__11175,N__11400,N__11634,N__14898,N__15129,N__15360}),
            .MASK({dangling_wire_154,dangling_wire_155,dangling_wire_156,dangling_wire_157,dangling_wire_158,dangling_wire_159,dangling_wire_160,dangling_wire_161,dangling_wire_162,dangling_wire_163,dangling_wire_164,dangling_wire_165,dangling_wire_166,dangling_wire_167,dangling_wire_168,dangling_wire_169}),
            .WDATA({dangling_wire_170,dangling_wire_171,dangling_wire_172,dangling_wire_173,N__8626,dangling_wire_174,dangling_wire_175,dangling_wire_176,dangling_wire_177,dangling_wire_178,dangling_wire_179,dangling_wire_180,N__8515,dangling_wire_181,dangling_wire_182,dangling_wire_183}),
            .RCLKE(),
            .RCLK(N__22676),
            .RE(N__23344),
            .WCLKE(),
            .WCLK(N__19333),
            .WE(N__10227));
    defparam \line_buffer.mem21_physical .WRITE_MODE=3;
    defparam \line_buffer.mem21_physical .READ_MODE=3;
    defparam \line_buffer.mem21_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem21_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem21_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem21_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem21_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem21_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem21_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem21_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem21_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem21_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem21_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem21_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem21_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem21_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem21_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem21_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem21_physical  (
            .RDATA({dangling_wire_184,dangling_wire_185,dangling_wire_186,dangling_wire_187,\line_buffer.n676 ,dangling_wire_188,dangling_wire_189,dangling_wire_190,dangling_wire_191,dangling_wire_192,dangling_wire_193,dangling_wire_194,\line_buffer.n675 ,dangling_wire_195,dangling_wire_196,dangling_wire_197}),
            .RADDR({N__9816,N__16143,N__16809,N__16473,N__15489,N__18543,N__18777,N__19947,N__13926,N__18102,N__10716}),
            .WADDR({N__12780,N__13038,N__11790,N__12048,N__12315,N__11043,N__11268,N__11502,N__14766,N__14997,N__15228}),
            .MASK({dangling_wire_198,dangling_wire_199,dangling_wire_200,dangling_wire_201,dangling_wire_202,dangling_wire_203,dangling_wire_204,dangling_wire_205,dangling_wire_206,dangling_wire_207,dangling_wire_208,dangling_wire_209,dangling_wire_210,dangling_wire_211,dangling_wire_212,dangling_wire_213}),
            .WDATA({dangling_wire_214,dangling_wire_215,dangling_wire_216,dangling_wire_217,N__8447,dangling_wire_218,dangling_wire_219,dangling_wire_220,dangling_wire_221,dangling_wire_222,dangling_wire_223,dangling_wire_224,N__8347,dangling_wire_225,dangling_wire_226,dangling_wire_227}),
            .RCLKE(),
            .RCLK(N__22386),
            .RE(N__23138),
            .WCLKE(),
            .WCLK(N__19365),
            .WE(N__13486));
    defparam \line_buffer.mem12_physical .WRITE_MODE=3;
    defparam \line_buffer.mem12_physical .READ_MODE=3;
    defparam \line_buffer.mem12_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem12_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem12_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem12_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem12_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem12_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem12_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem12_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem12_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem12_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem12_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem12_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem12_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem12_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem12_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem12_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem12_physical  (
            .RDATA({dangling_wire_228,dangling_wire_229,dangling_wire_230,dangling_wire_231,\line_buffer.n612 ,dangling_wire_232,dangling_wire_233,dangling_wire_234,dangling_wire_235,dangling_wire_236,dangling_wire_237,dangling_wire_238,\line_buffer.n611 ,dangling_wire_239,dangling_wire_240,dangling_wire_241}),
            .RADDR({N__9936,N__16263,N__16929,N__16593,N__15609,N__18663,N__18897,N__20067,N__14046,N__18222,N__10836}),
            .WADDR({N__12900,N__13158,N__11910,N__12168,N__12435,N__11163,N__11388,N__11622,N__14886,N__15117,N__15348}),
            .MASK({dangling_wire_242,dangling_wire_243,dangling_wire_244,dangling_wire_245,dangling_wire_246,dangling_wire_247,dangling_wire_248,dangling_wire_249,dangling_wire_250,dangling_wire_251,dangling_wire_252,dangling_wire_253,dangling_wire_254,dangling_wire_255,dangling_wire_256,dangling_wire_257}),
            .WDATA({dangling_wire_258,dangling_wire_259,dangling_wire_260,dangling_wire_261,N__8417,dangling_wire_262,dangling_wire_263,dangling_wire_264,dangling_wire_265,dangling_wire_266,dangling_wire_267,dangling_wire_268,N__8335,dangling_wire_269,dangling_wire_270,dangling_wire_271}),
            .RCLKE(),
            .RCLK(N__22655),
            .RE(N__23311),
            .WCLKE(),
            .WCLK(N__19341),
            .WE(N__10226));
    defparam \line_buffer.mem18_physical .WRITE_MODE=3;
    defparam \line_buffer.mem18_physical .READ_MODE=3;
    defparam \line_buffer.mem18_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem18_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem18_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem18_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem18_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem18_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem18_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem18_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem18_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem18_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem18_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem18_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem18_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem18_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem18_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem18_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem18_physical  (
            .RDATA({dangling_wire_272,dangling_wire_273,dangling_wire_274,dangling_wire_275,\line_buffer.n555 ,dangling_wire_276,dangling_wire_277,dangling_wire_278,dangling_wire_279,dangling_wire_280,dangling_wire_281,dangling_wire_282,\line_buffer.n554 ,dangling_wire_283,dangling_wire_284,dangling_wire_285}),
            .RADDR({N__9864,N__16191,N__16857,N__16521,N__15537,N__18591,N__18825,N__19995,N__13974,N__18150,N__10764}),
            .WADDR({N__12828,N__13086,N__11838,N__12096,N__12363,N__11091,N__11316,N__11550,N__14814,N__15045,N__15276}),
            .MASK({dangling_wire_286,dangling_wire_287,dangling_wire_288,dangling_wire_289,dangling_wire_290,dangling_wire_291,dangling_wire_292,dangling_wire_293,dangling_wire_294,dangling_wire_295,dangling_wire_296,dangling_wire_297,dangling_wire_298,dangling_wire_299,dangling_wire_300,dangling_wire_301}),
            .WDATA({dangling_wire_302,dangling_wire_303,dangling_wire_304,dangling_wire_305,N__8451,dangling_wire_306,dangling_wire_307,dangling_wire_308,dangling_wire_309,dangling_wire_310,dangling_wire_311,dangling_wire_312,N__8336,dangling_wire_313,dangling_wire_314,dangling_wire_315}),
            .RCLKE(),
            .RCLK(N__22516),
            .RE(N__23124),
            .WCLKE(),
            .WCLK(N__19354),
            .WE(N__12606));
    defparam \line_buffer.mem24_physical .WRITE_MODE=3;
    defparam \line_buffer.mem24_physical .READ_MODE=3;
    defparam \line_buffer.mem24_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem24_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem24_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem24_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem24_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem24_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem24_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem24_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem24_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem24_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem24_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem24_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem24_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem24_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem24_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem24_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem24_physical  (
            .RDATA({dangling_wire_316,dangling_wire_317,dangling_wire_318,dangling_wire_319,\line_buffer.n620 ,dangling_wire_320,dangling_wire_321,dangling_wire_322,dangling_wire_323,dangling_wire_324,dangling_wire_325,dangling_wire_326,\line_buffer.n619 ,dangling_wire_327,dangling_wire_328,dangling_wire_329}),
            .RADDR({N__9963,N__16296,N__16962,N__16626,N__15636,N__18702,N__18930,N__20106,N__14085,N__18249,N__10857}),
            .WADDR({N__12945,N__13197,N__11949,N__12201,N__12456,N__11196,N__11415,N__11643,N__14913,N__15150,N__15387}),
            .MASK({dangling_wire_330,dangling_wire_331,dangling_wire_332,dangling_wire_333,dangling_wire_334,dangling_wire_335,dangling_wire_336,dangling_wire_337,dangling_wire_338,dangling_wire_339,dangling_wire_340,dangling_wire_341,dangling_wire_342,dangling_wire_343,dangling_wire_344,dangling_wire_345}),
            .WDATA({dangling_wire_346,dangling_wire_347,dangling_wire_348,dangling_wire_349,N__8380,dangling_wire_350,dangling_wire_351,dangling_wire_352,dangling_wire_353,dangling_wire_354,dangling_wire_355,dangling_wire_356,N__8258,dangling_wire_357,dangling_wire_358,dangling_wire_359}),
            .RCLKE(),
            .RCLK(N__22407),
            .RE(N__23394),
            .WCLKE(),
            .WCLK(N__19328),
            .WE(N__12656));
    defparam \line_buffer.mem1_physical .WRITE_MODE=3;
    defparam \line_buffer.mem1_physical .READ_MODE=3;
    defparam \line_buffer.mem1_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem1_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem1_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem1_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem1_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem1_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem1_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem1_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem1_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem1_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem1_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem1_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem1_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem1_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem1_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem1_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem1_physical  (
            .RDATA({dangling_wire_360,dangling_wire_361,dangling_wire_362,dangling_wire_363,\line_buffer.n648 ,dangling_wire_364,dangling_wire_365,dangling_wire_366,dangling_wire_367,dangling_wire_368,dangling_wire_369,dangling_wire_370,\line_buffer.n647 ,dangling_wire_371,dangling_wire_372,dangling_wire_373}),
            .RADDR({N__9972,N__16299,N__16965,N__16629,N__15645,N__18699,N__18933,N__20103,N__14082,N__18258,N__10870}),
            .WADDR({N__12936,N__13194,N__11946,N__12204,N__12469,N__11199,N__11424,N__11656,N__14922,N__15153,N__15384}),
            .MASK({dangling_wire_374,dangling_wire_375,dangling_wire_376,dangling_wire_377,dangling_wire_378,dangling_wire_379,dangling_wire_380,dangling_wire_381,dangling_wire_382,dangling_wire_383,dangling_wire_384,dangling_wire_385,dangling_wire_386,dangling_wire_387,dangling_wire_388,dangling_wire_389}),
            .WDATA({dangling_wire_390,dangling_wire_391,dangling_wire_392,dangling_wire_393,N__8722,dangling_wire_394,dangling_wire_395,dangling_wire_396,dangling_wire_397,dangling_wire_398,dangling_wire_399,dangling_wire_400,N__8840,dangling_wire_401,dangling_wire_402,dangling_wire_403}),
            .RCLKE(),
            .RCLK(N__22688),
            .RE(N__23370),
            .WCLKE(),
            .WCLK(N__19325),
            .WE(N__15719));
    defparam \line_buffer.mem15_physical .WRITE_MODE=3;
    defparam \line_buffer.mem15_physical .READ_MODE=3;
    defparam \line_buffer.mem15_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem15_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem15_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem15_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem15_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem15_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem15_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem15_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem15_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem15_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem15_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem15_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem15_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem15_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem15_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem15_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem15_physical  (
            .RDATA({dangling_wire_404,dangling_wire_405,dangling_wire_406,dangling_wire_407,\line_buffer.n644 ,dangling_wire_408,dangling_wire_409,dangling_wire_410,dangling_wire_411,dangling_wire_412,dangling_wire_413,dangling_wire_414,\line_buffer.n643 ,dangling_wire_415,dangling_wire_416,dangling_wire_417}),
            .RADDR({N__9900,N__16227,N__16893,N__16557,N__15573,N__18627,N__18861,N__20031,N__14010,N__18186,N__10800}),
            .WADDR({N__12864,N__13122,N__11874,N__12132,N__12399,N__11127,N__11352,N__11586,N__14850,N__15081,N__15312}),
            .MASK({dangling_wire_418,dangling_wire_419,dangling_wire_420,dangling_wire_421,dangling_wire_422,dangling_wire_423,dangling_wire_424,dangling_wire_425,dangling_wire_426,dangling_wire_427,dangling_wire_428,dangling_wire_429,dangling_wire_430,dangling_wire_431,dangling_wire_432,dangling_wire_433}),
            .WDATA({dangling_wire_434,dangling_wire_435,dangling_wire_436,dangling_wire_437,N__8433,dangling_wire_438,dangling_wire_439,dangling_wire_440,dangling_wire_441,dangling_wire_442,dangling_wire_443,dangling_wire_444,N__8325,dangling_wire_445,dangling_wire_446,dangling_wire_447}),
            .RCLKE(),
            .RCLK(N__22622),
            .RE(N__23260),
            .WCLKE(),
            .WCLK(N__19348),
            .WE(N__15720));
    defparam \line_buffer.mem27_physical .WRITE_MODE=3;
    defparam \line_buffer.mem27_physical .READ_MODE=3;
    defparam \line_buffer.mem27_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem27_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem27_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem27_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem27_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem27_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem27_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem27_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem27_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem27_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem27_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem27_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem27_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem27_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem27_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem27_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem27_physical  (
            .RDATA({dangling_wire_448,dangling_wire_449,dangling_wire_450,dangling_wire_451,\line_buffer.n652 ,dangling_wire_452,dangling_wire_453,dangling_wire_454,dangling_wire_455,dangling_wire_456,dangling_wire_457,dangling_wire_458,\line_buffer.n651 ,dangling_wire_459,dangling_wire_460,dangling_wire_461}),
            .RADDR({N__9927,N__16260,N__16926,N__16590,N__15600,N__18666,N__18894,N__20070,N__14049,N__18213,N__10821}),
            .WADDR({N__12909,N__13161,N__11913,N__12165,N__12420,N__11160,N__11379,N__11607,N__14877,N__15114,N__15351}),
            .MASK({dangling_wire_462,dangling_wire_463,dangling_wire_464,dangling_wire_465,dangling_wire_466,dangling_wire_467,dangling_wire_468,dangling_wire_469,dangling_wire_470,dangling_wire_471,dangling_wire_472,dangling_wire_473,dangling_wire_474,dangling_wire_475,dangling_wire_476,dangling_wire_477}),
            .WDATA({dangling_wire_478,dangling_wire_479,dangling_wire_480,dangling_wire_481,N__8411,dangling_wire_482,dangling_wire_483,dangling_wire_484,dangling_wire_485,dangling_wire_486,dangling_wire_487,dangling_wire_488,N__8289,dangling_wire_489,dangling_wire_490,dangling_wire_491}),
            .RCLKE(),
            .RCLK(N__22640),
            .RE(N__23373),
            .WCLKE(),
            .WCLK(N__19343),
            .WE(N__10113));
    defparam \line_buffer.mem4_physical .WRITE_MODE=3;
    defparam \line_buffer.mem4_physical .READ_MODE=3;
    defparam \line_buffer.mem4_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem4_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem4_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem4_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem4_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem4_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem4_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem4_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem4_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem4_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem4_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem4_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem4_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem4_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem4_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem4_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem4_physical  (
            .RDATA({dangling_wire_492,dangling_wire_493,dangling_wire_494,dangling_wire_495,\line_buffer.n624 ,dangling_wire_496,dangling_wire_497,dangling_wire_498,dangling_wire_499,dangling_wire_500,dangling_wire_501,dangling_wire_502,\line_buffer.n623 ,dangling_wire_503,dangling_wire_504,dangling_wire_505}),
            .RADDR({N__9855,N__16188,N__16854,N__16518,N__15528,N__18594,N__18822,N__19998,N__13977,N__18141,N__10749}),
            .WADDR({N__12837,N__13089,N__11841,N__12093,N__12348,N__11088,N__11307,N__11535,N__14805,N__15042,N__15279}),
            .MASK({dangling_wire_506,dangling_wire_507,dangling_wire_508,dangling_wire_509,dangling_wire_510,dangling_wire_511,dangling_wire_512,dangling_wire_513,dangling_wire_514,dangling_wire_515,dangling_wire_516,dangling_wire_517,dangling_wire_518,dangling_wire_519,dangling_wire_520,dangling_wire_521}),
            .WDATA({dangling_wire_522,dangling_wire_523,dangling_wire_524,dangling_wire_525,N__8750,dangling_wire_526,dangling_wire_527,dangling_wire_528,dangling_wire_529,dangling_wire_530,dangling_wire_531,dangling_wire_532,N__8875,dangling_wire_533,dangling_wire_534,dangling_wire_535}),
            .RCLKE(),
            .RCLK(N__22488),
            .RE(N__23282),
            .WCLKE(),
            .WCLK(N__19355),
            .WE(N__12658));
    defparam \line_buffer.mem16_physical .WRITE_MODE=3;
    defparam \line_buffer.mem16_physical .READ_MODE=3;
    defparam \line_buffer.mem16_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem16_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem16_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem16_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem16_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem16_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem16_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem16_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem16_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem16_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem16_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem16_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem16_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem16_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem16_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem16_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem16_physical  (
            .RDATA({dangling_wire_536,dangling_wire_537,dangling_wire_538,dangling_wire_539,\line_buffer.n642 ,dangling_wire_540,dangling_wire_541,dangling_wire_542,dangling_wire_543,dangling_wire_544,dangling_wire_545,dangling_wire_546,\line_buffer.n641 ,dangling_wire_547,dangling_wire_548,dangling_wire_549}),
            .RADDR({N__9888,N__16215,N__16881,N__16545,N__15561,N__18615,N__18849,N__20019,N__13998,N__18174,N__10788}),
            .WADDR({N__12852,N__13110,N__11862,N__12120,N__12387,N__11115,N__11340,N__11574,N__14838,N__15069,N__15300}),
            .MASK({dangling_wire_550,dangling_wire_551,dangling_wire_552,dangling_wire_553,dangling_wire_554,dangling_wire_555,dangling_wire_556,dangling_wire_557,dangling_wire_558,dangling_wire_559,dangling_wire_560,dangling_wire_561,dangling_wire_562,dangling_wire_563,dangling_wire_564,dangling_wire_565}),
            .WDATA({dangling_wire_566,dangling_wire_567,dangling_wire_568,dangling_wire_569,N__8214,dangling_wire_570,dangling_wire_571,dangling_wire_572,dangling_wire_573,dangling_wire_574,dangling_wire_575,dangling_wire_576,N__8997,dangling_wire_577,dangling_wire_578,dangling_wire_579}),
            .RCLKE(),
            .RCLK(N__22583),
            .RE(N__23192),
            .WCLKE(),
            .WCLK(N__19350),
            .WE(N__15721));
    defparam \line_buffer.mem30_physical .WRITE_MODE=3;
    defparam \line_buffer.mem30_physical .READ_MODE=3;
    defparam \line_buffer.mem30_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem30_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem30_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem30_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem30_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem30_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem30_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem30_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem30_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem30_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem30_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem30_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem30_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem30_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem30_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem30_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem30_physical  (
            .RDATA({dangling_wire_580,dangling_wire_581,dangling_wire_582,dangling_wire_583,\line_buffer.n684 ,dangling_wire_584,dangling_wire_585,dangling_wire_586,dangling_wire_587,dangling_wire_588,dangling_wire_589,dangling_wire_590,\line_buffer.n683 ,dangling_wire_591,dangling_wire_592,dangling_wire_593}),
            .RADDR({N__9879,N__16212,N__16878,N__16542,N__15552,N__18618,N__18846,N__20022,N__14001,N__18165,N__10773}),
            .WADDR({N__12861,N__13113,N__11865,N__12117,N__12372,N__11112,N__11331,N__11559,N__14829,N__15066,N__15303}),
            .MASK({dangling_wire_594,dangling_wire_595,dangling_wire_596,dangling_wire_597,dangling_wire_598,dangling_wire_599,dangling_wire_600,dangling_wire_601,dangling_wire_602,dangling_wire_603,dangling_wire_604,dangling_wire_605,dangling_wire_606,dangling_wire_607,dangling_wire_608,dangling_wire_609}),
            .WDATA({dangling_wire_610,dangling_wire_611,dangling_wire_612,dangling_wire_613,N__8440,dangling_wire_614,dangling_wire_615,dangling_wire_616,dangling_wire_617,dangling_wire_618,dangling_wire_619,dangling_wire_620,N__8321,dangling_wire_621,dangling_wire_622,dangling_wire_623}),
            .RCLKE(),
            .RCLK(N__22579),
            .RE(N__23326),
            .WCLKE(),
            .WCLK(N__19351),
            .WE(N__10262));
    defparam \line_buffer.mem7_physical .WRITE_MODE=3;
    defparam \line_buffer.mem7_physical .READ_MODE=3;
    defparam \line_buffer.mem7_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem7_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem7_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem7_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem7_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem7_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem7_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem7_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem7_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem7_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem7_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem7_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem7_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem7_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem7_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem7_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem7_physical  (
            .RDATA({dangling_wire_624,dangling_wire_625,dangling_wire_626,dangling_wire_627,\line_buffer.n551 ,dangling_wire_628,dangling_wire_629,dangling_wire_630,dangling_wire_631,dangling_wire_632,dangling_wire_633,dangling_wire_634,\line_buffer.n550 ,dangling_wire_635,dangling_wire_636,dangling_wire_637}),
            .RADDR({N__9819,N__16152,N__16818,N__16482,N__15492,N__18558,N__18786,N__19962,N__13941,N__18105,N__10713}),
            .WADDR({N__12801,N__13053,N__11805,N__12057,N__12312,N__11052,N__11271,N__11499,N__14769,N__15006,N__15243}),
            .MASK({dangling_wire_638,dangling_wire_639,dangling_wire_640,dangling_wire_641,dangling_wire_642,dangling_wire_643,dangling_wire_644,dangling_wire_645,dangling_wire_646,dangling_wire_647,dangling_wire_648,dangling_wire_649,dangling_wire_650,dangling_wire_651,dangling_wire_652,dangling_wire_653}),
            .WDATA({dangling_wire_654,dangling_wire_655,dangling_wire_656,dangling_wire_657,N__8773,dangling_wire_658,dangling_wire_659,dangling_wire_660,dangling_wire_661,dangling_wire_662,dangling_wire_663,dangling_wire_664,N__8884,dangling_wire_665,dangling_wire_666,dangling_wire_667}),
            .RCLKE(),
            .RCLK(N__22020),
            .RE(N__23228),
            .WCLKE(),
            .WCLK(N__19364),
            .WE(N__10181));
    defparam \line_buffer.mem20_physical .WRITE_MODE=3;
    defparam \line_buffer.mem20_physical .READ_MODE=3;
    defparam \line_buffer.mem20_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem20_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem20_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem20_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem20_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem20_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem20_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem20_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem20_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem20_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem20_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem20_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem20_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem20_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem20_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem20_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem20_physical  (
            .RDATA({dangling_wire_668,dangling_wire_669,dangling_wire_670,dangling_wire_671,\line_buffer.n678 ,dangling_wire_672,dangling_wire_673,dangling_wire_674,dangling_wire_675,dangling_wire_676,dangling_wire_677,dangling_wire_678,\line_buffer.n677 ,dangling_wire_679,dangling_wire_680,dangling_wire_681}),
            .RADDR({N__9828,N__16155,N__16821,N__16485,N__15501,N__18555,N__18789,N__19959,N__13938,N__18114,N__10728}),
            .WADDR({N__12792,N__13050,N__11802,N__12060,N__12327,N__11055,N__11280,N__11514,N__14778,N__15009,N__15240}),
            .MASK({dangling_wire_682,dangling_wire_683,dangling_wire_684,dangling_wire_685,dangling_wire_686,dangling_wire_687,dangling_wire_688,dangling_wire_689,dangling_wire_690,dangling_wire_691,dangling_wire_692,dangling_wire_693,dangling_wire_694,dangling_wire_695,dangling_wire_696,dangling_wire_697}),
            .WDATA({dangling_wire_698,dangling_wire_699,dangling_wire_700,dangling_wire_701,N__8665,dangling_wire_702,dangling_wire_703,dangling_wire_704,dangling_wire_705,dangling_wire_706,dangling_wire_707,dangling_wire_708,N__8557,dangling_wire_709,dangling_wire_710,dangling_wire_711}),
            .RCLKE(),
            .RCLK(N__22205),
            .RE(N__23190),
            .WCLKE(),
            .WCLK(N__19363),
            .WE(N__13475));
    defparam \line_buffer.mem13_physical .WRITE_MODE=3;
    defparam \line_buffer.mem13_physical .READ_MODE=3;
    defparam \line_buffer.mem13_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem13_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem13_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem13_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem13_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem13_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem13_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem13_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem13_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem13_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem13_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem13_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem13_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem13_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem13_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem13_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem13_physical  (
            .RDATA({dangling_wire_712,dangling_wire_713,dangling_wire_714,dangling_wire_715,\line_buffer.n610 ,dangling_wire_716,dangling_wire_717,dangling_wire_718,dangling_wire_719,dangling_wire_720,dangling_wire_721,dangling_wire_722,\line_buffer.n609 ,dangling_wire_723,dangling_wire_724,dangling_wire_725}),
            .RADDR({N__9924,N__16251,N__16917,N__16581,N__15597,N__18651,N__18885,N__20055,N__14034,N__18210,N__10824}),
            .WADDR({N__12888,N__13146,N__11898,N__12156,N__12423,N__11151,N__11376,N__11610,N__14874,N__15105,N__15336}),
            .MASK({dangling_wire_726,dangling_wire_727,dangling_wire_728,dangling_wire_729,dangling_wire_730,dangling_wire_731,dangling_wire_732,dangling_wire_733,dangling_wire_734,dangling_wire_735,dangling_wire_736,dangling_wire_737,dangling_wire_738,dangling_wire_739,dangling_wire_740,dangling_wire_741}),
            .WDATA({dangling_wire_742,dangling_wire_743,dangling_wire_744,dangling_wire_745,N__8193,dangling_wire_746,dangling_wire_747,dangling_wire_748,dangling_wire_749,dangling_wire_750,dangling_wire_751,dangling_wire_752,N__8990,dangling_wire_753,dangling_wire_754,dangling_wire_755}),
            .RCLKE(),
            .RCLK(N__22654),
            .RE(N__23310),
            .WCLKE(),
            .WCLK(N__19344),
            .WE(N__10225));
    defparam \line_buffer.mem19_physical .WRITE_MODE=3;
    defparam \line_buffer.mem19_physical .READ_MODE=3;
    defparam \line_buffer.mem19_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem19_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem19_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem19_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem19_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem19_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem19_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem19_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem19_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem19_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem19_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem19_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem19_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem19_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem19_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem19_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem19_physical  (
            .RDATA({dangling_wire_756,dangling_wire_757,dangling_wire_758,dangling_wire_759,\line_buffer.n553 ,dangling_wire_760,dangling_wire_761,dangling_wire_762,dangling_wire_763,dangling_wire_764,dangling_wire_765,dangling_wire_766,\line_buffer.n552 ,dangling_wire_767,dangling_wire_768,dangling_wire_769}),
            .RADDR({N__9852,N__16179,N__16845,N__16509,N__15525,N__18579,N__18813,N__19983,N__13962,N__18138,N__10752}),
            .WADDR({N__12816,N__13074,N__11826,N__12084,N__12351,N__11079,N__11304,N__11538,N__14802,N__15033,N__15264}),
            .MASK({dangling_wire_770,dangling_wire_771,dangling_wire_772,dangling_wire_773,dangling_wire_774,dangling_wire_775,dangling_wire_776,dangling_wire_777,dangling_wire_778,dangling_wire_779,dangling_wire_780,dangling_wire_781,dangling_wire_782,dangling_wire_783,dangling_wire_784,dangling_wire_785}),
            .WDATA({dangling_wire_786,dangling_wire_787,dangling_wire_788,dangling_wire_789,N__8206,dangling_wire_790,dangling_wire_791,dangling_wire_792,dangling_wire_793,dangling_wire_794,dangling_wire_795,dangling_wire_796,N__9009,dangling_wire_797,dangling_wire_798,dangling_wire_799}),
            .RCLKE(),
            .RCLK(N__22515),
            .RE(N__23117),
            .WCLKE(),
            .WCLK(N__19359),
            .WE(N__12605));
    defparam \line_buffer.mem23_physical .WRITE_MODE=3;
    defparam \line_buffer.mem23_physical .READ_MODE=3;
    defparam \line_buffer.mem23_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem23_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem23_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem23_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem23_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem23_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem23_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem23_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem23_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem23_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem23_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem23_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem23_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem23_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem23_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem23_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem23_physical  (
            .RDATA({dangling_wire_800,dangling_wire_801,dangling_wire_802,dangling_wire_803,\line_buffer.n622 ,dangling_wire_804,dangling_wire_805,dangling_wire_806,dangling_wire_807,dangling_wire_808,dangling_wire_809,dangling_wire_810,\line_buffer.n621 ,dangling_wire_811,dangling_wire_812,dangling_wire_813}),
            .RADDR({N__9975,N__16308,N__16974,N__16638,N__15648,N__18712,N__18942,N__20116,N__14095,N__18261,N__10869}),
            .WADDR({N__12952,N__13207,N__11959,N__12213,N__12468,N__11208,N__11427,N__11655,N__14925,N__15162,N__15397}),
            .MASK({dangling_wire_814,dangling_wire_815,dangling_wire_816,dangling_wire_817,dangling_wire_818,dangling_wire_819,dangling_wire_820,dangling_wire_821,dangling_wire_822,dangling_wire_823,dangling_wire_824,dangling_wire_825,dangling_wire_826,dangling_wire_827,dangling_wire_828,dangling_wire_829}),
            .WDATA({dangling_wire_830,dangling_wire_831,dangling_wire_832,dangling_wire_833,N__8642,dangling_wire_834,dangling_wire_835,dangling_wire_836,dangling_wire_837,dangling_wire_838,dangling_wire_839,dangling_wire_840,N__8483,dangling_wire_841,dangling_wire_842,dangling_wire_843}),
            .RCLKE(),
            .RCLK(N__22690),
            .RE(N__23395),
            .WCLKE(),
            .WCLK(N__19323),
            .WE(N__12657));
    defparam \line_buffer.mem0_physical .WRITE_MODE=3;
    defparam \line_buffer.mem0_physical .READ_MODE=3;
    defparam \line_buffer.mem0_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem0_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem0_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem0_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem0_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem0_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem0_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem0_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem0_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem0_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem0_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem0_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem0_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem0_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem0_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem0_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem0_physical  (
            .RDATA({dangling_wire_844,dangling_wire_845,dangling_wire_846,dangling_wire_847,\line_buffer.n616 ,dangling_wire_848,dangling_wire_849,dangling_wire_850,dangling_wire_851,dangling_wire_852,dangling_wire_853,dangling_wire_854,\line_buffer.n615 ,dangling_wire_855,dangling_wire_856,dangling_wire_857}),
            .RADDR({N__9979,N__16309,N__16975,N__16639,N__15652,N__18711,N__18943,N__20115,N__14094,N__18265,N__10876}),
            .WADDR({N__12948,N__13206,N__11958,N__12214,N__12475,N__11209,N__11431,N__11662,N__14929,N__15163,N__15396}),
            .MASK({dangling_wire_858,dangling_wire_859,dangling_wire_860,dangling_wire_861,dangling_wire_862,dangling_wire_863,dangling_wire_864,dangling_wire_865,dangling_wire_866,dangling_wire_867,dangling_wire_868,dangling_wire_869,dangling_wire_870,dangling_wire_871,dangling_wire_872,dangling_wire_873}),
            .WDATA({dangling_wire_874,dangling_wire_875,dangling_wire_876,dangling_wire_877,N__8697,dangling_wire_878,dangling_wire_879,dangling_wire_880,dangling_wire_881,dangling_wire_882,dangling_wire_883,dangling_wire_884,N__8839,dangling_wire_885,dangling_wire_886,dangling_wire_887}),
            .RCLKE(),
            .RCLK(N__22689),
            .RE(N__23371),
            .WCLKE(),
            .WCLK(N__19321),
            .WE(N__10234));
    defparam \line_buffer.mem26_physical .WRITE_MODE=3;
    defparam \line_buffer.mem26_physical .READ_MODE=3;
    defparam \line_buffer.mem26_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem26_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem26_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem26_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem26_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem26_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem26_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem26_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem26_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem26_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem26_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem26_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem26_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem26_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem26_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem26_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem26_physical  (
            .RDATA({dangling_wire_888,dangling_wire_889,dangling_wire_890,dangling_wire_891,\line_buffer.n654 ,dangling_wire_892,dangling_wire_893,dangling_wire_894,dangling_wire_895,dangling_wire_896,dangling_wire_897,dangling_wire_898,\line_buffer.n653 ,dangling_wire_899,dangling_wire_900,dangling_wire_901}),
            .RADDR({N__9939,N__16272,N__16938,N__16602,N__15612,N__18678,N__18906,N__20082,N__14061,N__18225,N__10833}),
            .WADDR({N__12921,N__13173,N__11925,N__12177,N__12432,N__11172,N__11391,N__11619,N__14889,N__15126,N__15363}),
            .MASK({dangling_wire_902,dangling_wire_903,dangling_wire_904,dangling_wire_905,dangling_wire_906,dangling_wire_907,dangling_wire_908,dangling_wire_909,dangling_wire_910,dangling_wire_911,dangling_wire_912,dangling_wire_913,dangling_wire_914,dangling_wire_915,dangling_wire_916,dangling_wire_917}),
            .WDATA({dangling_wire_918,dangling_wire_919,dangling_wire_920,dangling_wire_921,N__8625,dangling_wire_922,dangling_wire_923,dangling_wire_924,dangling_wire_925,dangling_wire_926,dangling_wire_927,dangling_wire_928,N__8508,dangling_wire_929,dangling_wire_930,dangling_wire_931}),
            .RCLKE(),
            .RCLK(N__22668),
            .RE(N__23386),
            .WCLKE(),
            .WCLK(N__19337),
            .WE(N__10112));
    defparam \line_buffer.mem3_physical .WRITE_MODE=3;
    defparam \line_buffer.mem3_physical .READ_MODE=3;
    defparam \line_buffer.mem3_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem3_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem3_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem3_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem3_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem3_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem3_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem3_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem3_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem3_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem3_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem3_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem3_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem3_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem3_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem3_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem3_physical  (
            .RDATA({dangling_wire_932,dangling_wire_933,dangling_wire_934,dangling_wire_935,\line_buffer.n680 ,dangling_wire_936,dangling_wire_937,dangling_wire_938,dangling_wire_939,dangling_wire_940,dangling_wire_941,dangling_wire_942,\line_buffer.n679 ,dangling_wire_943,dangling_wire_944,dangling_wire_945}),
            .RADDR({N__9891,N__16224,N__16890,N__16554,N__15564,N__18630,N__18858,N__20034,N__14013,N__18177,N__10785}),
            .WADDR({N__12873,N__13125,N__11877,N__12129,N__12384,N__11124,N__11343,N__11571,N__14841,N__15078,N__15315}),
            .MASK({dangling_wire_946,dangling_wire_947,dangling_wire_948,dangling_wire_949,dangling_wire_950,dangling_wire_951,dangling_wire_952,dangling_wire_953,dangling_wire_954,dangling_wire_955,dangling_wire_956,dangling_wire_957,dangling_wire_958,dangling_wire_959,dangling_wire_960,dangling_wire_961}),
            .WDATA({dangling_wire_962,dangling_wire_963,dangling_wire_964,dangling_wire_965,N__8751,dangling_wire_966,dangling_wire_967,dangling_wire_968,dangling_wire_969,dangling_wire_970,dangling_wire_971,dangling_wire_972,N__8856,dangling_wire_973,dangling_wire_974,dangling_wire_975}),
            .RCLKE(),
            .RCLK(N__22538),
            .RE(N__23352),
            .WCLKE(),
            .WCLK(N__19349),
            .WE(N__13474));
    defparam \line_buffer.mem17_physical .WRITE_MODE=3;
    defparam \line_buffer.mem17_physical .READ_MODE=3;
    defparam \line_buffer.mem17_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem17_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem17_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem17_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem17_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem17_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem17_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem17_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem17_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem17_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem17_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem17_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem17_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem17_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem17_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem17_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem17_physical  (
            .RDATA({dangling_wire_976,dangling_wire_977,dangling_wire_978,dangling_wire_979,\line_buffer.n557 ,dangling_wire_980,dangling_wire_981,dangling_wire_982,dangling_wire_983,dangling_wire_984,dangling_wire_985,dangling_wire_986,\line_buffer.n556 ,dangling_wire_987,dangling_wire_988,dangling_wire_989}),
            .RADDR({N__9876,N__16203,N__16869,N__16533,N__15549,N__18603,N__18837,N__20007,N__13986,N__18162,N__10776}),
            .WADDR({N__12840,N__13098,N__11850,N__12108,N__12375,N__11103,N__11328,N__11562,N__14826,N__15057,N__15288}),
            .MASK({dangling_wire_990,dangling_wire_991,dangling_wire_992,dangling_wire_993,dangling_wire_994,dangling_wire_995,dangling_wire_996,dangling_wire_997,dangling_wire_998,dangling_wire_999,dangling_wire_1000,dangling_wire_1001,dangling_wire_1002,dangling_wire_1003,dangling_wire_1004,dangling_wire_1005}),
            .WDATA({dangling_wire_1006,dangling_wire_1007,dangling_wire_1008,dangling_wire_1009,N__8649,dangling_wire_1010,dangling_wire_1011,dangling_wire_1012,dangling_wire_1013,dangling_wire_1014,dangling_wire_1015,dangling_wire_1016,N__8546,dangling_wire_1017,dangling_wire_1018,dangling_wire_1019}),
            .RCLKE(),
            .RCLK(N__22582),
            .RE(N__23191),
            .WCLKE(),
            .WCLK(N__19352),
            .WE(N__12598));
    defparam \line_buffer.mem31_physical .WRITE_MODE=3;
    defparam \line_buffer.mem31_physical .READ_MODE=3;
    defparam \line_buffer.mem31_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem31_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem31_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem31_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem31_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem31_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem31_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem31_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem31_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem31_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem31_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem31_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem31_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem31_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem31_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem31_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem31_physical  (
            .RDATA({dangling_wire_1020,dangling_wire_1021,dangling_wire_1022,dangling_wire_1023,\line_buffer.n682 ,dangling_wire_1024,dangling_wire_1025,dangling_wire_1026,dangling_wire_1027,dangling_wire_1028,dangling_wire_1029,dangling_wire_1030,\line_buffer.n681 ,dangling_wire_1031,dangling_wire_1032,dangling_wire_1033}),
            .RADDR({N__9867,N__16200,N__16866,N__16530,N__15540,N__18606,N__18834,N__20010,N__13989,N__18153,N__10761}),
            .WADDR({N__12849,N__13101,N__11853,N__12105,N__12360,N__11100,N__11319,N__11547,N__14817,N__15054,N__15291}),
            .MASK({dangling_wire_1034,dangling_wire_1035,dangling_wire_1036,dangling_wire_1037,dangling_wire_1038,dangling_wire_1039,dangling_wire_1040,dangling_wire_1041,dangling_wire_1042,dangling_wire_1043,dangling_wire_1044,dangling_wire_1045,dangling_wire_1046,dangling_wire_1047,dangling_wire_1048,dangling_wire_1049}),
            .WDATA({dangling_wire_1050,dangling_wire_1051,dangling_wire_1052,dangling_wire_1053,N__8183,dangling_wire_1054,dangling_wire_1055,dangling_wire_1056,dangling_wire_1057,dangling_wire_1058,dangling_wire_1059,dangling_wire_1060,N__8974,dangling_wire_1061,dangling_wire_1062,dangling_wire_1063}),
            .RCLKE(),
            .RCLK(N__22436),
            .RE(N__23325),
            .WCLKE(),
            .WCLK(N__19353),
            .WE(N__10269));
    defparam \line_buffer.mem9_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem9_physical .WRITE_MODE=3;
    defparam \line_buffer.mem9_physical .READ_MODE=3;
    defparam \line_buffer.mem9_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem9_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem9_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem9_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem9_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem9_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem9_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem9_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem9_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem9_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem9_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem9_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem9_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem9_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem9_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem9_physical  (
            .RDATA({dangling_wire_1064,dangling_wire_1065,dangling_wire_1066,dangling_wire_1067,\line_buffer.n547 ,dangling_wire_1068,dangling_wire_1069,dangling_wire_1070,dangling_wire_1071,dangling_wire_1072,dangling_wire_1073,dangling_wire_1074,\line_buffer.n546 ,dangling_wire_1075,dangling_wire_1076,dangling_wire_1077}),
            .RADDR({N__9795,N__16128,N__16794,N__16458,N__15468,N__18534,N__18762,N__19938,N__13917,N__18081,N__10689}),
            .WADDR({N__12777,N__13029,N__11781,N__12033,N__12288,N__11028,N__11247,N__11475,N__14745,N__14982,N__15219}),
            .MASK({dangling_wire_1078,dangling_wire_1079,dangling_wire_1080,dangling_wire_1081,dangling_wire_1082,dangling_wire_1083,dangling_wire_1084,dangling_wire_1085,dangling_wire_1086,dangling_wire_1087,dangling_wire_1088,dangling_wire_1089,dangling_wire_1090,dangling_wire_1091,dangling_wire_1092,dangling_wire_1093}),
            .WDATA({dangling_wire_1094,dangling_wire_1095,dangling_wire_1096,dangling_wire_1097,N__8455,dangling_wire_1098,dangling_wire_1099,dangling_wire_1100,dangling_wire_1101,dangling_wire_1102,dangling_wire_1103,dangling_wire_1104,N__8346,dangling_wire_1105,dangling_wire_1106,dangling_wire_1107}),
            .RCLKE(),
            .RCLK(N__22037),
            .RE(N__23343),
            .WCLKE(),
            .WCLK(N__19368),
            .WE(N__10189));
    defparam \line_buffer.mem29_physical .WRITE_MODE=3;
    defparam \line_buffer.mem29_physical .READ_MODE=3;
    defparam \line_buffer.mem29_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem29_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem29_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem29_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem29_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem29_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem29_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem29_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem29_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem29_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem29_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem29_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem29_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem29_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem29_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem29_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem29_physical  (
            .RDATA({dangling_wire_1108,dangling_wire_1109,dangling_wire_1110,dangling_wire_1111,\line_buffer.n686 ,dangling_wire_1112,dangling_wire_1113,dangling_wire_1114,dangling_wire_1115,dangling_wire_1116,dangling_wire_1117,dangling_wire_1118,\line_buffer.n685 ,dangling_wire_1119,dangling_wire_1120,dangling_wire_1121}),
            .RADDR({N__9903,N__16236,N__16902,N__16566,N__15576,N__18642,N__18870,N__20046,N__14025,N__18189,N__10797}),
            .WADDR({N__12885,N__13137,N__11889,N__12141,N__12396,N__11136,N__11355,N__11583,N__14853,N__15090,N__15327}),
            .MASK({dangling_wire_1122,dangling_wire_1123,dangling_wire_1124,dangling_wire_1125,dangling_wire_1126,dangling_wire_1127,dangling_wire_1128,dangling_wire_1129,dangling_wire_1130,dangling_wire_1131,dangling_wire_1132,dangling_wire_1133,dangling_wire_1134,dangling_wire_1135,dangling_wire_1136,dangling_wire_1137}),
            .WDATA({dangling_wire_1138,dangling_wire_1139,dangling_wire_1140,dangling_wire_1141,N__8667,dangling_wire_1142,dangling_wire_1143,dangling_wire_1144,dangling_wire_1145,dangling_wire_1146,dangling_wire_1147,dangling_wire_1148,N__8521,dangling_wire_1149,dangling_wire_1150,dangling_wire_1151}),
            .RCLKE(),
            .RCLK(N__22675),
            .RE(N__23353),
            .WCLKE(),
            .WCLK(N__19347),
            .WE(N__10253));
    defparam \line_buffer.mem6_physical .WRITE_MODE=3;
    defparam \line_buffer.mem6_physical .READ_MODE=3;
    defparam \line_buffer.mem6_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem6_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem6_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem6_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem6_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem6_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem6_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem6_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem6_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem6_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem6_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem6_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem6_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem6_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem6_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem6_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem6_physical  (
            .RDATA({dangling_wire_1152,dangling_wire_1153,dangling_wire_1154,dangling_wire_1155,\line_buffer.n688 ,dangling_wire_1156,dangling_wire_1157,dangling_wire_1158,dangling_wire_1159,dangling_wire_1160,dangling_wire_1161,dangling_wire_1162,\line_buffer.n687 ,dangling_wire_1163,dangling_wire_1164,dangling_wire_1165}),
            .RADDR({N__9831,N__16164,N__16830,N__16494,N__15504,N__18570,N__18798,N__19974,N__13953,N__18117,N__10725}),
            .WADDR({N__12813,N__13065,N__11817,N__12069,N__12324,N__11064,N__11283,N__11511,N__14781,N__15018,N__15255}),
            .MASK({dangling_wire_1166,dangling_wire_1167,dangling_wire_1168,dangling_wire_1169,dangling_wire_1170,dangling_wire_1171,dangling_wire_1172,dangling_wire_1173,dangling_wire_1174,dangling_wire_1175,dangling_wire_1176,dangling_wire_1177,dangling_wire_1178,dangling_wire_1179,dangling_wire_1180,dangling_wire_1181}),
            .WDATA({dangling_wire_1182,dangling_wire_1183,dangling_wire_1184,dangling_wire_1185,N__8772,dangling_wire_1186,dangling_wire_1187,dangling_wire_1188,dangling_wire_1189,dangling_wire_1190,dangling_wire_1191,dangling_wire_1192,N__8883,dangling_wire_1193,dangling_wire_1194,dangling_wire_1195}),
            .RCLKE(),
            .RCLK(N__22408),
            .RE(N__23227),
            .WCLKE(),
            .WCLK(N__19362),
            .WE(N__10273));
    defparam \line_buffer.mem10_physical .WRITE_MODE=3;
    defparam \line_buffer.mem10_physical .READ_MODE=3;
    defparam \line_buffer.mem10_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem10_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem10_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem10_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem10_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem10_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem10_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem10_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem10_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem10_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem10_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem10_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem10_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem10_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem10_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem10_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem10_physical  (
            .RDATA({dangling_wire_1196,dangling_wire_1197,dangling_wire_1198,dangling_wire_1199,\line_buffer.n545 ,dangling_wire_1200,dangling_wire_1201,dangling_wire_1202,dangling_wire_1203,dangling_wire_1204,dangling_wire_1205,dangling_wire_1206,\line_buffer.n544 ,dangling_wire_1207,dangling_wire_1208,dangling_wire_1209}),
            .RADDR({N__9960,N__16287,N__16953,N__16617,N__15633,N__18687,N__18921,N__20091,N__14070,N__18246,N__10860}),
            .WADDR({N__12924,N__13182,N__11934,N__12192,N__12459,N__11187,N__11412,N__11646,N__14910,N__15141,N__15372}),
            .MASK({dangling_wire_1210,dangling_wire_1211,dangling_wire_1212,dangling_wire_1213,dangling_wire_1214,dangling_wire_1215,dangling_wire_1216,dangling_wire_1217,dangling_wire_1218,dangling_wire_1219,dangling_wire_1220,dangling_wire_1221,dangling_wire_1222,dangling_wire_1223,dangling_wire_1224,dangling_wire_1225}),
            .WDATA({dangling_wire_1226,dangling_wire_1227,dangling_wire_1228,dangling_wire_1229,N__8207,dangling_wire_1230,dangling_wire_1231,dangling_wire_1232,dangling_wire_1233,dangling_wire_1234,dangling_wire_1235,dangling_wire_1236,N__8975,dangling_wire_1237,dangling_wire_1238,dangling_wire_1239}),
            .RCLKE(),
            .RCLK(N__22677),
            .RE(N__23345),
            .WCLKE(),
            .WCLK(N__19331),
            .WE(N__10180));
    defparam \line_buffer.mem22_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem22_physical .WRITE_MODE=3;
    defparam \line_buffer.mem22_physical .READ_MODE=3;
    defparam \line_buffer.mem22_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem22_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem22_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem22_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem22_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem22_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem22_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem22_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem22_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem22_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem22_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem22_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem22_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem22_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem22_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem22_physical  (
            .RDATA({dangling_wire_1240,dangling_wire_1241,dangling_wire_1242,dangling_wire_1243,\line_buffer.n674 ,dangling_wire_1244,dangling_wire_1245,dangling_wire_1246,dangling_wire_1247,dangling_wire_1248,dangling_wire_1249,dangling_wire_1250,\line_buffer.n673 ,dangling_wire_1251,dangling_wire_1252,dangling_wire_1253}),
            .RADDR({N__9804,N__16131,N__16797,N__16461,N__15477,N__18531,N__18765,N__19935,N__13914,N__18090,N__10704}),
            .WADDR({N__12768,N__13026,N__11778,N__12036,N__12303,N__11031,N__11256,N__11490,N__14754,N__14985,N__15216}),
            .MASK({dangling_wire_1254,dangling_wire_1255,dangling_wire_1256,dangling_wire_1257,dangling_wire_1258,dangling_wire_1259,dangling_wire_1260,dangling_wire_1261,dangling_wire_1262,dangling_wire_1263,dangling_wire_1264,dangling_wire_1265,dangling_wire_1266,dangling_wire_1267,dangling_wire_1268,dangling_wire_1269}),
            .WDATA({dangling_wire_1270,dangling_wire_1271,dangling_wire_1272,dangling_wire_1273,N__8215,dangling_wire_1274,dangling_wire_1275,dangling_wire_1276,dangling_wire_1277,dangling_wire_1278,dangling_wire_1279,dangling_wire_1280,N__9016,dangling_wire_1281,dangling_wire_1282,dangling_wire_1283}),
            .RCLKE(),
            .RCLK(N__22239),
            .RE(N__23139),
            .WCLKE(),
            .WCLK(N__19367),
            .WE(N__13485));
    defparam \line_buffer.mem25_physical .WRITE_MODE=3;
    defparam \line_buffer.mem25_physical .READ_MODE=3;
    defparam \line_buffer.mem25_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem25_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem25_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem25_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem25_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem25_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem25_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem25_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem25_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem25_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem25_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem25_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem25_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem25_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem25_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem25_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem25_physical  (
            .RDATA({dangling_wire_1284,dangling_wire_1285,dangling_wire_1286,dangling_wire_1287,\line_buffer.n618 ,dangling_wire_1288,dangling_wire_1289,dangling_wire_1290,dangling_wire_1291,dangling_wire_1292,dangling_wire_1293,dangling_wire_1294,\line_buffer.n617 ,dangling_wire_1295,dangling_wire_1296,dangling_wire_1297}),
            .RADDR({N__9951,N__16284,N__16950,N__16614,N__15624,N__18690,N__18918,N__20094,N__14073,N__18237,N__10845}),
            .WADDR({N__12933,N__13185,N__11937,N__12189,N__12444,N__11184,N__11403,N__11631,N__14901,N__15138,N__15375}),
            .MASK({dangling_wire_1298,dangling_wire_1299,dangling_wire_1300,dangling_wire_1301,dangling_wire_1302,dangling_wire_1303,dangling_wire_1304,dangling_wire_1305,dangling_wire_1306,dangling_wire_1307,dangling_wire_1308,dangling_wire_1309,dangling_wire_1310,dangling_wire_1311,dangling_wire_1312,dangling_wire_1313}),
            .WDATA({dangling_wire_1314,dangling_wire_1315,dangling_wire_1316,dangling_wire_1317,N__8182,dangling_wire_1318,dangling_wire_1319,dangling_wire_1320,dangling_wire_1321,dangling_wire_1322,dangling_wire_1323,dangling_wire_1324,N__8941,dangling_wire_1325,dangling_wire_1326,dangling_wire_1327}),
            .RCLKE(),
            .RCLK(N__22684),
            .RE(N__23387),
            .WCLKE(),
            .WCLK(N__19332),
            .WE(N__12646));
    defparam \line_buffer.mem8_physical .WRITE_MODE=3;
    defparam \line_buffer.mem8_physical .READ_MODE=3;
    defparam \line_buffer.mem8_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem8_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem8_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem8_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem8_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem8_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem8_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem8_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem8_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem8_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem8_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem8_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem8_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem8_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem8_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem8_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem8_physical  (
            .RDATA({dangling_wire_1328,dangling_wire_1329,dangling_wire_1330,dangling_wire_1331,\line_buffer.n549 ,dangling_wire_1332,dangling_wire_1333,dangling_wire_1334,dangling_wire_1335,dangling_wire_1336,dangling_wire_1337,dangling_wire_1338,\line_buffer.n548 ,dangling_wire_1339,dangling_wire_1340,dangling_wire_1341}),
            .RADDR({N__9807,N__16140,N__16806,N__16470,N__15480,N__18546,N__18774,N__19950,N__13929,N__18093,N__10701}),
            .WADDR({N__12789,N__13041,N__11793,N__12045,N__12300,N__11040,N__11259,N__11487,N__14757,N__14994,N__15231}),
            .MASK({dangling_wire_1342,dangling_wire_1343,dangling_wire_1344,dangling_wire_1345,dangling_wire_1346,dangling_wire_1347,dangling_wire_1348,dangling_wire_1349,dangling_wire_1350,dangling_wire_1351,dangling_wire_1352,dangling_wire_1353,dangling_wire_1354,dangling_wire_1355,dangling_wire_1356,dangling_wire_1357}),
            .WDATA({dangling_wire_1358,dangling_wire_1359,dangling_wire_1360,dangling_wire_1361,N__8671,dangling_wire_1362,dangling_wire_1363,dangling_wire_1364,dangling_wire_1365,dangling_wire_1366,dangling_wire_1367,dangling_wire_1368,N__8556,dangling_wire_1369,dangling_wire_1370,dangling_wire_1371}),
            .RCLKE(),
            .RCLK(N__22225),
            .RE(N__23299),
            .WCLKE(),
            .WCLK(N__19366),
            .WE(N__10188));
    defparam \line_buffer.mem28_physical .WRITE_MODE=3;
    defparam \line_buffer.mem28_physical .READ_MODE=3;
    defparam \line_buffer.mem28_physical .INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem28_physical .INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem28_physical .INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem28_physical .INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem28_physical .INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem28_physical .INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem28_physical .INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem28_physical .INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem28_physical .INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem28_physical .INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem28_physical .INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem28_physical .INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem28_physical .INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem28_physical .INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem28_physical .INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam \line_buffer.mem28_physical .INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K \line_buffer.mem28_physical  (
            .RDATA({dangling_wire_1372,dangling_wire_1373,dangling_wire_1374,dangling_wire_1375,\line_buffer.n650 ,dangling_wire_1376,dangling_wire_1377,dangling_wire_1378,dangling_wire_1379,dangling_wire_1380,dangling_wire_1381,dangling_wire_1382,\line_buffer.n649 ,dangling_wire_1383,dangling_wire_1384,dangling_wire_1385}),
            .RADDR({N__9915,N__16248,N__16914,N__16578,N__15588,N__18654,N__18882,N__20058,N__14037,N__18201,N__10809}),
            .WADDR({N__12897,N__13149,N__11901,N__12153,N__12408,N__11148,N__11367,N__11595,N__14865,N__15102,N__15339}),
            .MASK({dangling_wire_1386,dangling_wire_1387,dangling_wire_1388,dangling_wire_1389,dangling_wire_1390,dangling_wire_1391,dangling_wire_1392,dangling_wire_1393,dangling_wire_1394,dangling_wire_1395,dangling_wire_1396,dangling_wire_1397,dangling_wire_1398,dangling_wire_1399,dangling_wire_1400,dangling_wire_1401}),
            .WDATA({dangling_wire_1402,dangling_wire_1403,dangling_wire_1404,dangling_wire_1405,N__8175,dangling_wire_1406,dangling_wire_1407,dangling_wire_1408,dangling_wire_1409,dangling_wire_1410,dangling_wire_1411,dangling_wire_1412,N__8954,dangling_wire_1413,dangling_wire_1414,dangling_wire_1415}),
            .RCLKE(),
            .RCLK(N__22600),
            .RE(N__23372),
            .WCLKE(),
            .WCLK(N__19345),
            .WE(N__10105));
    PRE_IO_GBUF DEBUG_c_1_pad_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__24374),
            .GLOBALBUFFEROUTPUT(DEBUG_c_1_c));
    defparam DEBUG_c_1_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_c_1_pad_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_c_1_pad_iopad (
            .OE(N__24376),
            .DIN(N__24375),
            .DOUT(N__24374),
            .PACKAGEPIN(TVP_CLK));
    defparam DEBUG_c_1_pad_preio.PIN_TYPE=6'b000001;
    defparam DEBUG_c_1_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_c_1_pad_preio (
            .PADOEN(N__24376),
            .PADOUT(N__24375),
            .PADIN(N__24374),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_CLK_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_CLK_pad_iopad.PULLUP=1'b0;
    IO_PAD ADV_CLK_pad_iopad (
            .OE(N__24365),
            .DIN(N__24364),
            .DOUT(N__24363),
            .PACKAGEPIN(ADV_CLK));
    defparam ADV_CLK_pad_preio.PIN_TYPE=6'b011001;
    defparam ADV_CLK_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_CLK_pad_preio (
            .PADOEN(N__24365),
            .PADOUT(N__24364),
            .PADIN(N__24363),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__22536),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_3_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_3_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_3_iopad (
            .OE(N__24356),
            .DIN(N__24355),
            .DOUT(N__24354),
            .PACKAGEPIN(DEBUG[3]));
    defparam DEBUG_pad_3_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_3_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_3_preio (
            .PADOEN(N__24356),
            .PADOUT(N__24355),
            .PADIN(N__24354),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__15769),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_VIDEO_pad_2_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_VIDEO_pad_2_iopad.PULLUP=1'b1;
    IO_PAD TVP_VIDEO_pad_2_iopad (
            .OE(N__24347),
            .DIN(N__24346),
            .DOUT(N__24345),
            .PACKAGEPIN(TVP_VIDEO[2]));
    defparam TVP_VIDEO_pad_2_preio.PIN_TYPE=6'b000001;
    defparam TVP_VIDEO_pad_2_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_VIDEO_pad_2_preio (
            .PADOEN(N__24347),
            .PADOUT(N__24346),
            .PADIN(N__24345),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_VIDEO_c_2),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_5_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_5_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_5_iopad (
            .OE(N__24338),
            .DIN(N__24337),
            .DOUT(N__24336),
            .PACKAGEPIN(ADV_G[5]));
    defparam ADV_G_pad_5_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_5_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_5_preio (
            .PADOEN(N__24338),
            .PADOUT(N__24337),
            .PADIN(N__24336),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__14304),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_3_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_3_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_3_iopad (
            .OE(N__24329),
            .DIN(N__24328),
            .DOUT(N__24327),
            .PACKAGEPIN(ADV_R[3]));
    defparam ADV_R_pad_3_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_3_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_3_preio (
            .PADOEN(N__24329),
            .PADOUT(N__24328),
            .PADIN(N__24327),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__14415),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_1_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_1_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_1_iopad (
            .OE(N__24320),
            .DIN(N__24319),
            .DOUT(N__24318),
            .PACKAGEPIN(ADV_G[1]));
    defparam ADV_G_pad_1_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_1_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_1_preio (
            .PADOEN(N__24320),
            .PADOUT(N__24319),
            .PADIN(N__24318),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__14524),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_0_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_0_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_0_iopad (
            .OE(N__24311),
            .DIN(N__24310),
            .DOUT(N__24309),
            .PACKAGEPIN(ADV_R[0]));
    defparam ADV_R_pad_0_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_0_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_0_preio (
            .PADOEN(N__24311),
            .PADOUT(N__24310),
            .PADIN(N__24309),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10047),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_2_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_2_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_2_iopad (
            .OE(N__24302),
            .DIN(N__24301),
            .DOUT(N__24300),
            .PACKAGEPIN(DEBUG[2]));
    defparam DEBUG_pad_2_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_2_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_2_preio (
            .PADOEN(N__24302),
            .PADOUT(N__24301),
            .PADIN(N__24300),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__22873),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_VIDEO_pad_3_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_VIDEO_pad_3_iopad.PULLUP=1'b1;
    IO_PAD TVP_VIDEO_pad_3_iopad (
            .OE(N__24293),
            .DIN(N__24292),
            .DOUT(N__24291),
            .PACKAGEPIN(TVP_VIDEO[3]));
    defparam TVP_VIDEO_pad_3_preio.PIN_TYPE=6'b000001;
    defparam TVP_VIDEO_pad_3_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_VIDEO_pad_3_preio (
            .PADOEN(N__24293),
            .PADOUT(N__24292),
            .PADIN(N__24291),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_VIDEO_c_3),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_4_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_4_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_4_iopad (
            .OE(N__24284),
            .DIN(N__24283),
            .DOUT(N__24282),
            .PACKAGEPIN(ADV_G[4]));
    defparam ADV_G_pad_4_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_4_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_4_preio (
            .PADOEN(N__24284),
            .PADOUT(N__24283),
            .PADIN(N__24282),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__14351),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_5_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_5_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_5_iopad (
            .OE(N__24275),
            .DIN(N__24274),
            .DOUT(N__24273),
            .PACKAGEPIN(ADV_R[5]));
    defparam ADV_R_pad_5_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_5_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_5_preio (
            .PADOEN(N__24275),
            .PADOUT(N__24274),
            .PADIN(N__24273),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__14300),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_VIDEO_pad_9_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_VIDEO_pad_9_iopad.PULLUP=1'b1;
    IO_PAD TVP_VIDEO_pad_9_iopad (
            .OE(N__24266),
            .DIN(N__24265),
            .DOUT(N__24264),
            .PACKAGEPIN(TVP_VIDEO[9]));
    defparam TVP_VIDEO_pad_9_preio.PIN_TYPE=6'b000001;
    defparam TVP_VIDEO_pad_9_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_VIDEO_pad_9_preio (
            .PADOEN(N__24266),
            .PADOUT(N__24265),
            .PADIN(N__24264),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_VIDEO_c_9),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_1_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_1_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_1_iopad (
            .OE(N__24257),
            .DIN(N__24256),
            .DOUT(N__24255),
            .PACKAGEPIN(DEBUG[1]));
    defparam DEBUG_pad_1_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_1_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_1_preio (
            .PADOEN(N__24257),
            .PADOUT(N__24256),
            .PADIN(N__24255),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__19222),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_1_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_1_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_1_iopad (
            .OE(N__24248),
            .DIN(N__24247),
            .DOUT(N__24246),
            .PACKAGEPIN(ADV_B[1]));
    defparam ADV_B_pad_1_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_1_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_1_preio (
            .PADOEN(N__24248),
            .PADOUT(N__24247),
            .PADIN(N__24246),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__14513),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_SYNC_N_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_SYNC_N_pad_iopad.PULLUP=1'b1;
    IO_PAD ADV_SYNC_N_pad_iopad (
            .OE(N__24239),
            .DIN(N__24238),
            .DOUT(N__24237),
            .PACKAGEPIN(ADV_SYNC_N));
    defparam ADV_SYNC_N_pad_preio.PIN_TYPE=6'b011001;
    defparam ADV_SYNC_N_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_SYNC_N_pad_preio (
            .PADOEN(N__24239),
            .PADOUT(N__24238),
            .PADIN(N__24237),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_6_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_6_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_6_iopad (
            .OE(N__24230),
            .DIN(N__24229),
            .DOUT(N__24228),
            .PACKAGEPIN(ADV_B[6]));
    defparam ADV_B_pad_6_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_6_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_6_preio (
            .PADOEN(N__24230),
            .PADOUT(N__24229),
            .PADIN(N__24228),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__14245),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_6_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_6_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_6_iopad (
            .OE(N__24221),
            .DIN(N__24220),
            .DOUT(N__24219),
            .PACKAGEPIN(DEBUG[6]));
    defparam DEBUG_pad_6_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_6_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_6_preio (
            .PADOEN(N__24221),
            .PADOUT(N__24220),
            .PADIN(N__24219),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9676),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_VIDEO_pad_7_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_VIDEO_pad_7_iopad.PULLUP=1'b1;
    IO_PAD TVP_VIDEO_pad_7_iopad (
            .OE(N__24212),
            .DIN(N__24211),
            .DOUT(N__24210),
            .PACKAGEPIN(TVP_VIDEO[7]));
    defparam TVP_VIDEO_pad_7_preio.PIN_TYPE=6'b000001;
    defparam TVP_VIDEO_pad_7_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_VIDEO_pad_7_preio (
            .PADOEN(N__24212),
            .PADOUT(N__24211),
            .PADIN(N__24210),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_VIDEO_c_7),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_0_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_0_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_0_iopad (
            .OE(N__24203),
            .DIN(N__24202),
            .DOUT(N__24201),
            .PACKAGEPIN(ADV_G[0]));
    defparam ADV_G_pad_0_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_0_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_0_preio (
            .PADOEN(N__24203),
            .PADOUT(N__24202),
            .PADIN(N__24201),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10054),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_1_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_1_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_1_iopad (
            .OE(N__24194),
            .DIN(N__24193),
            .DOUT(N__24192),
            .PACKAGEPIN(ADV_R[1]));
    defparam ADV_R_pad_1_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_1_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_1_preio (
            .PADOEN(N__24194),
            .PADOUT(N__24193),
            .PADIN(N__24192),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__14520),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_5_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_5_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_5_iopad (
            .OE(N__24185),
            .DIN(N__24184),
            .DOUT(N__24183),
            .PACKAGEPIN(DEBUG[5]));
    defparam DEBUG_pad_5_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_5_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_5_preio (
            .PADOEN(N__24185),
            .PADOUT(N__24184),
            .PADIN(N__24183),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__15856),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_HSYNC_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_HSYNC_pad_iopad.PULLUP=1'b1;
    IO_PAD TVP_HSYNC_pad_iopad (
            .OE(N__24176),
            .DIN(N__24175),
            .DOUT(N__24174),
            .PACKAGEPIN(TVP_HSYNC));
    defparam TVP_HSYNC_pad_preio.PIN_TYPE=6'b000001;
    defparam TVP_HSYNC_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_HSYNC_pad_preio (
            .PADOEN(N__24176),
            .PADOUT(N__24175),
            .PADIN(N__24174),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_HSYNC_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_7_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_7_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_7_iopad (
            .OE(N__24167),
            .DIN(N__24166),
            .DOUT(N__24165),
            .PACKAGEPIN(ADV_G[7]));
    defparam ADV_G_pad_7_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_7_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_7_preio (
            .PADOEN(N__24167),
            .PADOUT(N__24166),
            .PADIN(N__24165),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__14171),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_6_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_6_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_6_iopad (
            .OE(N__24158),
            .DIN(N__24157),
            .DOUT(N__24156),
            .PACKAGEPIN(ADV_R[6]));
    defparam ADV_R_pad_6_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_6_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_6_preio (
            .PADOEN(N__24158),
            .PADOUT(N__24157),
            .PADIN(N__24156),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__14243),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_VSYNC_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_VSYNC_pad_iopad.PULLUP=1'b1;
    IO_PAD TVP_VSYNC_pad_iopad (
            .OE(N__24149),
            .DIN(N__24148),
            .DOUT(N__24147),
            .PACKAGEPIN(TVP_VSYNC));
    defparam TVP_VSYNC_pad_preio.PIN_TYPE=6'b000001;
    defparam TVP_VSYNC_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_VSYNC_pad_preio (
            .PADOEN(N__24149),
            .PADOUT(N__24148),
            .PADIN(N__24147),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_VSYNC_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_BLANK_N_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_BLANK_N_pad_iopad.PULLUP=1'b1;
    IO_PAD ADV_BLANK_N_pad_iopad (
            .OE(N__24140),
            .DIN(N__24139),
            .DOUT(N__24138),
            .PACKAGEPIN(ADV_BLANK_N));
    defparam ADV_BLANK_N_pad_preio.PIN_TYPE=6'b011001;
    defparam ADV_BLANK_N_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_BLANK_N_pad_preio (
            .PADOEN(N__24140),
            .PADOUT(N__24139),
            .PADIN(N__24138),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__23323),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_0_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_0_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_0_iopad (
            .OE(N__24131),
            .DIN(N__24130),
            .DOUT(N__24129),
            .PACKAGEPIN(DEBUG[0]));
    defparam DEBUG_pad_0_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_0_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_0_preio (
            .PADOEN(N__24131),
            .PADOUT(N__24130),
            .PADIN(N__24129),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10075),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_2_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_2_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_2_iopad (
            .OE(N__24122),
            .DIN(N__24121),
            .DOUT(N__24120),
            .PACKAGEPIN(ADV_B[2]));
    defparam ADV_B_pad_2_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_2_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_2_preio (
            .PADOEN(N__24122),
            .PADOUT(N__24121),
            .PADIN(N__24120),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__14463),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_7_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_7_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_7_iopad (
            .OE(N__24113),
            .DIN(N__24112),
            .DOUT(N__24111),
            .PACKAGEPIN(ADV_B[7]));
    defparam ADV_B_pad_7_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_7_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_7_preio (
            .PADOEN(N__24113),
            .PADOUT(N__24112),
            .PADIN(N__24111),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__14182),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam LED_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam LED_pad_iopad.PULLUP=1'b0;
    IO_PAD LED_pad_iopad (
            .OE(N__24104),
            .DIN(N__24103),
            .DOUT(N__24102),
            .PACKAGEPIN(LED));
    defparam LED_pad_preio.PIN_TYPE=6'b011001;
    defparam LED_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO LED_pad_preio (
            .PADOEN(N__24104),
            .PADOUT(N__24103),
            .PADIN(N__24102),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__17359),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_VIDEO_pad_4_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_VIDEO_pad_4_iopad.PULLUP=1'b1;
    IO_PAD TVP_VIDEO_pad_4_iopad (
            .OE(N__24095),
            .DIN(N__24094),
            .DOUT(N__24093),
            .PACKAGEPIN(TVP_VIDEO[4]));
    defparam TVP_VIDEO_pad_4_preio.PIN_TYPE=6'b000001;
    defparam TVP_VIDEO_pad_4_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_VIDEO_pad_4_preio (
            .PADOEN(N__24095),
            .PADOUT(N__24094),
            .PADIN(N__24093),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_VIDEO_c_4),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_3_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_3_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_3_iopad (
            .OE(N__24086),
            .DIN(N__24085),
            .DOUT(N__24084),
            .PACKAGEPIN(ADV_G[3]));
    defparam ADV_G_pad_3_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_3_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_3_preio (
            .PADOEN(N__24086),
            .PADOUT(N__24085),
            .PADIN(N__24084),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__14411),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_HSYNC_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_HSYNC_pad_iopad.PULLUP=1'b0;
    IO_PAD ADV_HSYNC_pad_iopad (
            .OE(N__24077),
            .DIN(N__24076),
            .DOUT(N__24075),
            .PACKAGEPIN(ADV_HSYNC));
    defparam ADV_HSYNC_pad_preio.PIN_TYPE=6'b011001;
    defparam ADV_HSYNC_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_HSYNC_pad_preio (
            .PADOEN(N__24077),
            .PADOUT(N__24076),
            .PADIN(N__24075),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__16729),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_2_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_2_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_2_iopad (
            .OE(N__24068),
            .DIN(N__24067),
            .DOUT(N__24066),
            .PACKAGEPIN(ADV_R[2]));
    defparam ADV_R_pad_2_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_2_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_2_preio (
            .PADOEN(N__24068),
            .PADOUT(N__24067),
            .PADIN(N__24066),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__14462),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_4_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_4_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_4_iopad (
            .OE(N__24059),
            .DIN(N__24058),
            .DOUT(N__24057),
            .PACKAGEPIN(ADV_B[4]));
    defparam ADV_B_pad_4_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_4_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_4_preio (
            .PADOEN(N__24059),
            .PADOUT(N__24058),
            .PADIN(N__24057),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__14359),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_4_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_4_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_4_iopad (
            .OE(N__24050),
            .DIN(N__24049),
            .DOUT(N__24048),
            .PACKAGEPIN(DEBUG[4]));
    defparam DEBUG_pad_4_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_4_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_4_preio (
            .PADOEN(N__24050),
            .PADOUT(N__24049),
            .PADIN(N__24048),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10657),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_6_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_6_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_6_iopad (
            .OE(N__24041),
            .DIN(N__24040),
            .DOUT(N__24039),
            .PACKAGEPIN(ADV_G[6]));
    defparam ADV_G_pad_6_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_6_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_6_preio (
            .PADOEN(N__24041),
            .PADOUT(N__24040),
            .PADIN(N__24039),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__14244),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_7_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_7_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_7_iopad (
            .OE(N__24032),
            .DIN(N__24031),
            .DOUT(N__24030),
            .PACKAGEPIN(ADV_R[7]));
    defparam ADV_R_pad_7_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_7_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_7_preio (
            .PADOEN(N__24032),
            .PADOUT(N__24031),
            .PADIN(N__24030),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__14181),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_3_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_3_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_3_iopad (
            .OE(N__24023),
            .DIN(N__24022),
            .DOUT(N__24021),
            .PACKAGEPIN(ADV_B[3]));
    defparam ADV_B_pad_3_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_3_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_3_preio (
            .PADOEN(N__24023),
            .PADOUT(N__24022),
            .PADIN(N__24021),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__14416),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_R_pad_4_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_R_pad_4_iopad.PULLUP=1'b0;
    IO_PAD ADV_R_pad_4_iopad (
            .OE(N__24014),
            .DIN(N__24013),
            .DOUT(N__24012),
            .PACKAGEPIN(ADV_R[4]));
    defparam ADV_R_pad_4_preio.PIN_TYPE=6'b011001;
    defparam ADV_R_pad_4_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_R_pad_4_preio (
            .PADOEN(N__24014),
            .PADOUT(N__24013),
            .PADIN(N__24012),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__14352),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_VIDEO_pad_8_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_VIDEO_pad_8_iopad.PULLUP=1'b1;
    IO_PAD TVP_VIDEO_pad_8_iopad (
            .OE(N__24005),
            .DIN(N__24004),
            .DOUT(N__24003),
            .PACKAGEPIN(TVP_VIDEO[8]));
    defparam TVP_VIDEO_pad_8_preio.PIN_TYPE=6'b000001;
    defparam TVP_VIDEO_pad_8_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_VIDEO_pad_8_preio (
            .PADOEN(N__24005),
            .PADOUT(N__24004),
            .PADIN(N__24003),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_VIDEO_c_8),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_0_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_0_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_0_iopad (
            .OE(N__23996),
            .DIN(N__23995),
            .DOUT(N__23994),
            .PACKAGEPIN(ADV_B[0]));
    defparam ADV_B_pad_0_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_0_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_0_preio (
            .PADOEN(N__23996),
            .PADOUT(N__23995),
            .PADIN(N__23994),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__10040),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_VIDEO_pad_5_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_VIDEO_pad_5_iopad.PULLUP=1'b1;
    IO_PAD TVP_VIDEO_pad_5_iopad (
            .OE(N__23987),
            .DIN(N__23986),
            .DOUT(N__23985),
            .PACKAGEPIN(TVP_VIDEO[5]));
    defparam TVP_VIDEO_pad_5_preio.PIN_TYPE=6'b000001;
    defparam TVP_VIDEO_pad_5_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_VIDEO_pad_5_preio (
            .PADOEN(N__23987),
            .PADOUT(N__23986),
            .PADIN(N__23985),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_VIDEO_c_5),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_G_pad_2_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_G_pad_2_iopad.PULLUP=1'b0;
    IO_PAD ADV_G_pad_2_iopad (
            .OE(N__23978),
            .DIN(N__23977),
            .DOUT(N__23976),
            .PACKAGEPIN(ADV_G[2]));
    defparam ADV_G_pad_2_preio.PIN_TYPE=6'b011001;
    defparam ADV_G_pad_2_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_G_pad_2_preio (
            .PADOEN(N__23978),
            .PADOUT(N__23977),
            .PADIN(N__23976),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__14464),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_VSYNC_pad_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_VSYNC_pad_iopad.PULLUP=1'b0;
    IO_PAD ADV_VSYNC_pad_iopad (
            .OE(N__23969),
            .DIN(N__23968),
            .DOUT(N__23967),
            .PACKAGEPIN(ADV_VSYNC));
    defparam ADV_VSYNC_pad_preio.PIN_TYPE=6'b011001;
    defparam ADV_VSYNC_pad_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_VSYNC_pad_preio (
            .PADOEN(N__23969),
            .PADOUT(N__23968),
            .PADIN(N__23967),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__21171),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam ADV_B_pad_5_iopad.IO_STANDARD="SB_LVCMOS";
    defparam ADV_B_pad_5_iopad.PULLUP=1'b0;
    IO_PAD ADV_B_pad_5_iopad (
            .OE(N__23960),
            .DIN(N__23959),
            .DOUT(N__23958),
            .PACKAGEPIN(ADV_B[5]));
    defparam ADV_B_pad_5_preio.PIN_TYPE=6'b011001;
    defparam ADV_B_pad_5_preio.NEG_TRIGGER=1'b0;
    PRE_IO ADV_B_pad_5_preio (
            .PADOEN(N__23960),
            .PADOUT(N__23959),
            .PADIN(N__23958),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__14305),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam DEBUG_pad_7_iopad.IO_STANDARD="SB_LVCMOS";
    defparam DEBUG_pad_7_iopad.PULLUP=1'b1;
    IO_PAD DEBUG_pad_7_iopad (
            .OE(N__23951),
            .DIN(N__23950),
            .DOUT(N__23949),
            .PACKAGEPIN(DEBUG[7]));
    defparam DEBUG_pad_7_preio.PIN_TYPE=6'b011001;
    defparam DEBUG_pad_7_preio.NEG_TRIGGER=1'b0;
    PRE_IO DEBUG_pad_7_preio (
            .PADOEN(N__23951),
            .PADOUT(N__23950),
            .PADIN(N__23949),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__23385),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam TVP_VIDEO_pad_6_iopad.IO_STANDARD="SB_LVCMOS";
    defparam TVP_VIDEO_pad_6_iopad.PULLUP=1'b1;
    IO_PAD TVP_VIDEO_pad_6_iopad (
            .OE(N__23942),
            .DIN(N__23941),
            .DOUT(N__23940),
            .PACKAGEPIN(TVP_VIDEO[6]));
    defparam TVP_VIDEO_pad_6_preio.PIN_TYPE=6'b000001;
    defparam TVP_VIDEO_pad_6_preio.NEG_TRIGGER=1'b0;
    PRE_IO TVP_VIDEO_pad_6_preio (
            .PADOEN(N__23942),
            .PADOUT(N__23941),
            .PADIN(N__23940),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(TVP_VIDEO_c_6),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__5782 (
            .O(N__23923),
            .I(N__23920));
    LocalMux I__5781 (
            .O(N__23920),
            .I(N__23917));
    Span12Mux_h I__5780 (
            .O(N__23917),
            .I(N__23914));
    Span12Mux_v I__5779 (
            .O(N__23914),
            .I(N__23911));
    Odrv12 I__5778 (
            .O(N__23911),
            .I(\line_buffer.n548 ));
    InMux I__5777 (
            .O(N__23908),
            .I(N__23905));
    LocalMux I__5776 (
            .O(N__23905),
            .I(N__23902));
    Span4Mux_h I__5775 (
            .O(N__23902),
            .I(N__23899));
    Span4Mux_h I__5774 (
            .O(N__23899),
            .I(N__23896));
    Odrv4 I__5773 (
            .O(N__23896),
            .I(\line_buffer.n556 ));
    CascadeMux I__5772 (
            .O(N__23893),
            .I(N__23890));
    InMux I__5771 (
            .O(N__23890),
            .I(N__23887));
    LocalMux I__5770 (
            .O(N__23887),
            .I(N__23884));
    Odrv12 I__5769 (
            .O(N__23884),
            .I(\line_buffer.n4077 ));
    InMux I__5768 (
            .O(N__23881),
            .I(N__23878));
    LocalMux I__5767 (
            .O(N__23878),
            .I(N__23875));
    Span4Mux_v I__5766 (
            .O(N__23875),
            .I(N__23872));
    Span4Mux_h I__5765 (
            .O(N__23872),
            .I(N__23869));
    Sp12to4 I__5764 (
            .O(N__23869),
            .I(N__23866));
    Odrv12 I__5763 (
            .O(N__23866),
            .I(\line_buffer.n674 ));
    InMux I__5762 (
            .O(N__23863),
            .I(N__23860));
    LocalMux I__5761 (
            .O(N__23860),
            .I(N__23856));
    InMux I__5760 (
            .O(N__23859),
            .I(N__23852));
    Span4Mux_v I__5759 (
            .O(N__23856),
            .I(N__23833));
    InMux I__5758 (
            .O(N__23855),
            .I(N__23830));
    LocalMux I__5757 (
            .O(N__23852),
            .I(N__23825));
    InMux I__5756 (
            .O(N__23851),
            .I(N__23822));
    InMux I__5755 (
            .O(N__23850),
            .I(N__23819));
    InMux I__5754 (
            .O(N__23849),
            .I(N__23813));
    InMux I__5753 (
            .O(N__23848),
            .I(N__23813));
    InMux I__5752 (
            .O(N__23847),
            .I(N__23808));
    InMux I__5751 (
            .O(N__23846),
            .I(N__23808));
    InMux I__5750 (
            .O(N__23845),
            .I(N__23803));
    InMux I__5749 (
            .O(N__23844),
            .I(N__23800));
    InMux I__5748 (
            .O(N__23843),
            .I(N__23795));
    InMux I__5747 (
            .O(N__23842),
            .I(N__23795));
    InMux I__5746 (
            .O(N__23841),
            .I(N__23790));
    InMux I__5745 (
            .O(N__23840),
            .I(N__23790));
    InMux I__5744 (
            .O(N__23839),
            .I(N__23783));
    InMux I__5743 (
            .O(N__23838),
            .I(N__23783));
    InMux I__5742 (
            .O(N__23837),
            .I(N__23783));
    InMux I__5741 (
            .O(N__23836),
            .I(N__23780));
    Span4Mux_h I__5740 (
            .O(N__23833),
            .I(N__23775));
    LocalMux I__5739 (
            .O(N__23830),
            .I(N__23775));
    InMux I__5738 (
            .O(N__23829),
            .I(N__23772));
    InMux I__5737 (
            .O(N__23828),
            .I(N__23769));
    Span4Mux_v I__5736 (
            .O(N__23825),
            .I(N__23762));
    LocalMux I__5735 (
            .O(N__23822),
            .I(N__23762));
    LocalMux I__5734 (
            .O(N__23819),
            .I(N__23762));
    InMux I__5733 (
            .O(N__23818),
            .I(N__23759));
    LocalMux I__5732 (
            .O(N__23813),
            .I(N__23756));
    LocalMux I__5731 (
            .O(N__23808),
            .I(N__23753));
    InMux I__5730 (
            .O(N__23807),
            .I(N__23750));
    CascadeMux I__5729 (
            .O(N__23806),
            .I(N__23747));
    LocalMux I__5728 (
            .O(N__23803),
            .I(N__23742));
    LocalMux I__5727 (
            .O(N__23800),
            .I(N__23742));
    LocalMux I__5726 (
            .O(N__23795),
            .I(N__23736));
    LocalMux I__5725 (
            .O(N__23790),
            .I(N__23736));
    LocalMux I__5724 (
            .O(N__23783),
            .I(N__23731));
    LocalMux I__5723 (
            .O(N__23780),
            .I(N__23731));
    Span4Mux_h I__5722 (
            .O(N__23775),
            .I(N__23720));
    LocalMux I__5721 (
            .O(N__23772),
            .I(N__23720));
    LocalMux I__5720 (
            .O(N__23769),
            .I(N__23720));
    Span4Mux_v I__5719 (
            .O(N__23762),
            .I(N__23720));
    LocalMux I__5718 (
            .O(N__23759),
            .I(N__23720));
    Span4Mux_h I__5717 (
            .O(N__23756),
            .I(N__23715));
    Span4Mux_h I__5716 (
            .O(N__23753),
            .I(N__23715));
    LocalMux I__5715 (
            .O(N__23750),
            .I(N__23712));
    InMux I__5714 (
            .O(N__23747),
            .I(N__23709));
    Span4Mux_h I__5713 (
            .O(N__23742),
            .I(N__23706));
    InMux I__5712 (
            .O(N__23741),
            .I(N__23703));
    Span4Mux_h I__5711 (
            .O(N__23736),
            .I(N__23700));
    Span12Mux_h I__5710 (
            .O(N__23731),
            .I(N__23697));
    Span4Mux_h I__5709 (
            .O(N__23720),
            .I(N__23694));
    Span4Mux_v I__5708 (
            .O(N__23715),
            .I(N__23685));
    Span4Mux_h I__5707 (
            .O(N__23712),
            .I(N__23685));
    LocalMux I__5706 (
            .O(N__23709),
            .I(N__23685));
    Span4Mux_h I__5705 (
            .O(N__23706),
            .I(N__23685));
    LocalMux I__5704 (
            .O(N__23703),
            .I(TX_ADDR_12));
    Odrv4 I__5703 (
            .O(N__23700),
            .I(TX_ADDR_12));
    Odrv12 I__5702 (
            .O(N__23697),
            .I(TX_ADDR_12));
    Odrv4 I__5701 (
            .O(N__23694),
            .I(TX_ADDR_12));
    Odrv4 I__5700 (
            .O(N__23685),
            .I(TX_ADDR_12));
    CascadeMux I__5699 (
            .O(N__23674),
            .I(N__23671));
    InMux I__5698 (
            .O(N__23671),
            .I(N__23668));
    LocalMux I__5697 (
            .O(N__23668),
            .I(N__23665));
    Span12Mux_h I__5696 (
            .O(N__23665),
            .I(N__23662));
    Odrv12 I__5695 (
            .O(N__23662),
            .I(\line_buffer.n682 ));
    InMux I__5694 (
            .O(N__23659),
            .I(N__23656));
    LocalMux I__5693 (
            .O(N__23656),
            .I(\line_buffer.n4158 ));
    InMux I__5692 (
            .O(N__23653),
            .I(N__23650));
    LocalMux I__5691 (
            .O(N__23650),
            .I(N__23647));
    Span4Mux_v I__5690 (
            .O(N__23647),
            .I(N__23644));
    Sp12to4 I__5689 (
            .O(N__23644),
            .I(N__23641));
    Span12Mux_h I__5688 (
            .O(N__23641),
            .I(N__23638));
    Odrv12 I__5687 (
            .O(N__23638),
            .I(\line_buffer.n685 ));
    InMux I__5686 (
            .O(N__23635),
            .I(N__23632));
    LocalMux I__5685 (
            .O(N__23632),
            .I(N__23629));
    Span4Mux_v I__5684 (
            .O(N__23629),
            .I(N__23626));
    Span4Mux_v I__5683 (
            .O(N__23626),
            .I(N__23623));
    Span4Mux_v I__5682 (
            .O(N__23623),
            .I(N__23620));
    Span4Mux_h I__5681 (
            .O(N__23620),
            .I(N__23617));
    Odrv4 I__5680 (
            .O(N__23617),
            .I(\line_buffer.n677 ));
    InMux I__5679 (
            .O(N__23614),
            .I(N__23608));
    CascadeMux I__5678 (
            .O(N__23613),
            .I(N__23605));
    InMux I__5677 (
            .O(N__23612),
            .I(N__23595));
    InMux I__5676 (
            .O(N__23611),
            .I(N__23592));
    LocalMux I__5675 (
            .O(N__23608),
            .I(N__23587));
    InMux I__5674 (
            .O(N__23605),
            .I(N__23583));
    InMux I__5673 (
            .O(N__23604),
            .I(N__23578));
    InMux I__5672 (
            .O(N__23603),
            .I(N__23578));
    InMux I__5671 (
            .O(N__23602),
            .I(N__23573));
    InMux I__5670 (
            .O(N__23601),
            .I(N__23570));
    InMux I__5669 (
            .O(N__23600),
            .I(N__23563));
    InMux I__5668 (
            .O(N__23599),
            .I(N__23563));
    InMux I__5667 (
            .O(N__23598),
            .I(N__23563));
    LocalMux I__5666 (
            .O(N__23595),
            .I(N__23560));
    LocalMux I__5665 (
            .O(N__23592),
            .I(N__23557));
    InMux I__5664 (
            .O(N__23591),
            .I(N__23554));
    InMux I__5663 (
            .O(N__23590),
            .I(N__23550));
    Span4Mux_v I__5662 (
            .O(N__23587),
            .I(N__23547));
    InMux I__5661 (
            .O(N__23586),
            .I(N__23544));
    LocalMux I__5660 (
            .O(N__23583),
            .I(N__23540));
    LocalMux I__5659 (
            .O(N__23578),
            .I(N__23537));
    InMux I__5658 (
            .O(N__23577),
            .I(N__23532));
    InMux I__5657 (
            .O(N__23576),
            .I(N__23529));
    LocalMux I__5656 (
            .O(N__23573),
            .I(N__23522));
    LocalMux I__5655 (
            .O(N__23570),
            .I(N__23522));
    LocalMux I__5654 (
            .O(N__23563),
            .I(N__23522));
    Span4Mux_h I__5653 (
            .O(N__23560),
            .I(N__23519));
    Span4Mux_h I__5652 (
            .O(N__23557),
            .I(N__23513));
    LocalMux I__5651 (
            .O(N__23554),
            .I(N__23513));
    InMux I__5650 (
            .O(N__23553),
            .I(N__23510));
    LocalMux I__5649 (
            .O(N__23550),
            .I(N__23503));
    Span4Mux_v I__5648 (
            .O(N__23547),
            .I(N__23503));
    LocalMux I__5647 (
            .O(N__23544),
            .I(N__23503));
    InMux I__5646 (
            .O(N__23543),
            .I(N__23500));
    Span4Mux_h I__5645 (
            .O(N__23540),
            .I(N__23497));
    Span4Mux_h I__5644 (
            .O(N__23537),
            .I(N__23494));
    InMux I__5643 (
            .O(N__23536),
            .I(N__23489));
    InMux I__5642 (
            .O(N__23535),
            .I(N__23486));
    LocalMux I__5641 (
            .O(N__23532),
            .I(N__23482));
    LocalMux I__5640 (
            .O(N__23529),
            .I(N__23479));
    Span4Mux_v I__5639 (
            .O(N__23522),
            .I(N__23474));
    Span4Mux_v I__5638 (
            .O(N__23519),
            .I(N__23474));
    InMux I__5637 (
            .O(N__23518),
            .I(N__23471));
    Span4Mux_v I__5636 (
            .O(N__23513),
            .I(N__23468));
    LocalMux I__5635 (
            .O(N__23510),
            .I(N__23465));
    Span4Mux_v I__5634 (
            .O(N__23503),
            .I(N__23462));
    LocalMux I__5633 (
            .O(N__23500),
            .I(N__23459));
    Span4Mux_v I__5632 (
            .O(N__23497),
            .I(N__23454));
    Span4Mux_v I__5631 (
            .O(N__23494),
            .I(N__23454));
    InMux I__5630 (
            .O(N__23493),
            .I(N__23449));
    InMux I__5629 (
            .O(N__23492),
            .I(N__23449));
    LocalMux I__5628 (
            .O(N__23489),
            .I(N__23444));
    LocalMux I__5627 (
            .O(N__23486),
            .I(N__23444));
    InMux I__5626 (
            .O(N__23485),
            .I(N__23441));
    Span12Mux_h I__5625 (
            .O(N__23482),
            .I(N__23438));
    Span4Mux_h I__5624 (
            .O(N__23479),
            .I(N__23431));
    Span4Mux_h I__5623 (
            .O(N__23474),
            .I(N__23431));
    LocalMux I__5622 (
            .O(N__23471),
            .I(N__23431));
    Span4Mux_v I__5621 (
            .O(N__23468),
            .I(N__23422));
    Span4Mux_v I__5620 (
            .O(N__23465),
            .I(N__23422));
    Span4Mux_h I__5619 (
            .O(N__23462),
            .I(N__23422));
    Span4Mux_h I__5618 (
            .O(N__23459),
            .I(N__23422));
    Span4Mux_h I__5617 (
            .O(N__23454),
            .I(N__23419));
    LocalMux I__5616 (
            .O(N__23449),
            .I(N__23414));
    Span12Mux_h I__5615 (
            .O(N__23444),
            .I(N__23414));
    LocalMux I__5614 (
            .O(N__23441),
            .I(TX_ADDR_11));
    Odrv12 I__5613 (
            .O(N__23438),
            .I(TX_ADDR_11));
    Odrv4 I__5612 (
            .O(N__23431),
            .I(TX_ADDR_11));
    Odrv4 I__5611 (
            .O(N__23422),
            .I(TX_ADDR_11));
    Odrv4 I__5610 (
            .O(N__23419),
            .I(TX_ADDR_11));
    Odrv12 I__5609 (
            .O(N__23414),
            .I(TX_ADDR_11));
    InMux I__5608 (
            .O(N__23401),
            .I(N__23398));
    LocalMux I__5607 (
            .O(N__23398),
            .I(\line_buffer.n4063 ));
    SRMux I__5606 (
            .O(N__23395),
            .I(N__23391));
    SRMux I__5605 (
            .O(N__23394),
            .I(N__23388));
    LocalMux I__5604 (
            .O(N__23391),
            .I(N__23380));
    LocalMux I__5603 (
            .O(N__23388),
            .I(N__23380));
    SRMux I__5602 (
            .O(N__23387),
            .I(N__23377));
    SRMux I__5601 (
            .O(N__23386),
            .I(N__23374));
    IoInMux I__5600 (
            .O(N__23385),
            .I(N__23367));
    Span4Mux_s3_v I__5599 (
            .O(N__23380),
            .I(N__23360));
    LocalMux I__5598 (
            .O(N__23377),
            .I(N__23360));
    LocalMux I__5597 (
            .O(N__23374),
            .I(N__23360));
    SRMux I__5596 (
            .O(N__23373),
            .I(N__23357));
    SRMux I__5595 (
            .O(N__23372),
            .I(N__23354));
    SRMux I__5594 (
            .O(N__23371),
            .I(N__23349));
    SRMux I__5593 (
            .O(N__23370),
            .I(N__23346));
    LocalMux I__5592 (
            .O(N__23367),
            .I(N__23340));
    Span4Mux_v I__5591 (
            .O(N__23360),
            .I(N__23333));
    LocalMux I__5590 (
            .O(N__23357),
            .I(N__23333));
    LocalMux I__5589 (
            .O(N__23354),
            .I(N__23333));
    SRMux I__5588 (
            .O(N__23353),
            .I(N__23330));
    SRMux I__5587 (
            .O(N__23352),
            .I(N__23327));
    LocalMux I__5586 (
            .O(N__23349),
            .I(N__23318));
    LocalMux I__5585 (
            .O(N__23346),
            .I(N__23318));
    SRMux I__5584 (
            .O(N__23345),
            .I(N__23315));
    SRMux I__5583 (
            .O(N__23344),
            .I(N__23312));
    SRMux I__5582 (
            .O(N__23343),
            .I(N__23300));
    Span4Mux_s0_h I__5581 (
            .O(N__23340),
            .I(N__23296));
    Span4Mux_v I__5580 (
            .O(N__23333),
            .I(N__23289));
    LocalMux I__5579 (
            .O(N__23330),
            .I(N__23289));
    LocalMux I__5578 (
            .O(N__23327),
            .I(N__23289));
    SRMux I__5577 (
            .O(N__23326),
            .I(N__23286));
    SRMux I__5576 (
            .O(N__23325),
            .I(N__23283));
    IoInMux I__5575 (
            .O(N__23324),
            .I(N__23278));
    IoInMux I__5574 (
            .O(N__23323),
            .I(N__23275));
    Span4Mux_s3_v I__5573 (
            .O(N__23318),
            .I(N__23268));
    LocalMux I__5572 (
            .O(N__23315),
            .I(N__23268));
    LocalMux I__5571 (
            .O(N__23312),
            .I(N__23268));
    SRMux I__5570 (
            .O(N__23311),
            .I(N__23265));
    SRMux I__5569 (
            .O(N__23310),
            .I(N__23262));
    CascadeMux I__5568 (
            .O(N__23309),
            .I(N__23257));
    CascadeMux I__5567 (
            .O(N__23308),
            .I(N__23253));
    CascadeMux I__5566 (
            .O(N__23307),
            .I(N__23249));
    CascadeMux I__5565 (
            .O(N__23306),
            .I(N__23246));
    CascadeMux I__5564 (
            .O(N__23305),
            .I(N__23242));
    CascadeMux I__5563 (
            .O(N__23304),
            .I(N__23239));
    CascadeMux I__5562 (
            .O(N__23303),
            .I(N__23235));
    LocalMux I__5561 (
            .O(N__23300),
            .I(N__23232));
    SRMux I__5560 (
            .O(N__23299),
            .I(N__23229));
    Span4Mux_h I__5559 (
            .O(N__23296),
            .I(N__23224));
    Span4Mux_v I__5558 (
            .O(N__23289),
            .I(N__23217));
    LocalMux I__5557 (
            .O(N__23286),
            .I(N__23217));
    LocalMux I__5556 (
            .O(N__23283),
            .I(N__23217));
    SRMux I__5555 (
            .O(N__23282),
            .I(N__23214));
    SRMux I__5554 (
            .O(N__23281),
            .I(N__23211));
    LocalMux I__5553 (
            .O(N__23278),
            .I(N__23206));
    LocalMux I__5552 (
            .O(N__23275),
            .I(N__23206));
    Span4Mux_v I__5551 (
            .O(N__23268),
            .I(N__23199));
    LocalMux I__5550 (
            .O(N__23265),
            .I(N__23199));
    LocalMux I__5549 (
            .O(N__23262),
            .I(N__23199));
    SRMux I__5548 (
            .O(N__23261),
            .I(N__23196));
    SRMux I__5547 (
            .O(N__23260),
            .I(N__23193));
    InMux I__5546 (
            .O(N__23257),
            .I(N__23178));
    InMux I__5545 (
            .O(N__23256),
            .I(N__23178));
    InMux I__5544 (
            .O(N__23253),
            .I(N__23178));
    InMux I__5543 (
            .O(N__23252),
            .I(N__23178));
    InMux I__5542 (
            .O(N__23249),
            .I(N__23178));
    InMux I__5541 (
            .O(N__23246),
            .I(N__23175));
    InMux I__5540 (
            .O(N__23245),
            .I(N__23164));
    InMux I__5539 (
            .O(N__23242),
            .I(N__23164));
    InMux I__5538 (
            .O(N__23239),
            .I(N__23164));
    InMux I__5537 (
            .O(N__23238),
            .I(N__23164));
    InMux I__5536 (
            .O(N__23235),
            .I(N__23164));
    Span4Mux_v I__5535 (
            .O(N__23232),
            .I(N__23161));
    LocalMux I__5534 (
            .O(N__23229),
            .I(N__23158));
    SRMux I__5533 (
            .O(N__23228),
            .I(N__23155));
    SRMux I__5532 (
            .O(N__23227),
            .I(N__23152));
    Span4Mux_h I__5531 (
            .O(N__23224),
            .I(N__23143));
    Span4Mux_v I__5530 (
            .O(N__23217),
            .I(N__23143));
    LocalMux I__5529 (
            .O(N__23214),
            .I(N__23143));
    LocalMux I__5528 (
            .O(N__23211),
            .I(N__23143));
    IoSpan4Mux I__5527 (
            .O(N__23206),
            .I(N__23140));
    Span4Mux_v I__5526 (
            .O(N__23199),
            .I(N__23131));
    LocalMux I__5525 (
            .O(N__23196),
            .I(N__23131));
    LocalMux I__5524 (
            .O(N__23193),
            .I(N__23131));
    SRMux I__5523 (
            .O(N__23192),
            .I(N__23128));
    SRMux I__5522 (
            .O(N__23191),
            .I(N__23125));
    SRMux I__5521 (
            .O(N__23190),
            .I(N__23121));
    SRMux I__5520 (
            .O(N__23189),
            .I(N__23118));
    LocalMux I__5519 (
            .O(N__23178),
            .I(N__23112));
    LocalMux I__5518 (
            .O(N__23175),
            .I(N__23112));
    LocalMux I__5517 (
            .O(N__23164),
            .I(N__23109));
    Span4Mux_h I__5516 (
            .O(N__23161),
            .I(N__23098));
    Span4Mux_v I__5515 (
            .O(N__23158),
            .I(N__23098));
    LocalMux I__5514 (
            .O(N__23155),
            .I(N__23098));
    LocalMux I__5513 (
            .O(N__23152),
            .I(N__23098));
    Span4Mux_v I__5512 (
            .O(N__23143),
            .I(N__23098));
    Span4Mux_s0_v I__5511 (
            .O(N__23140),
            .I(N__23095));
    SRMux I__5510 (
            .O(N__23139),
            .I(N__23092));
    SRMux I__5509 (
            .O(N__23138),
            .I(N__23089));
    Span4Mux_v I__5508 (
            .O(N__23131),
            .I(N__23082));
    LocalMux I__5507 (
            .O(N__23128),
            .I(N__23082));
    LocalMux I__5506 (
            .O(N__23125),
            .I(N__23082));
    SRMux I__5505 (
            .O(N__23124),
            .I(N__23079));
    LocalMux I__5504 (
            .O(N__23121),
            .I(N__23074));
    LocalMux I__5503 (
            .O(N__23118),
            .I(N__23074));
    SRMux I__5502 (
            .O(N__23117),
            .I(N__23071));
    Sp12to4 I__5501 (
            .O(N__23112),
            .I(N__23068));
    Span4Mux_v I__5500 (
            .O(N__23109),
            .I(N__23065));
    Span4Mux_v I__5499 (
            .O(N__23098),
            .I(N__23062));
    Span4Mux_h I__5498 (
            .O(N__23095),
            .I(N__23055));
    LocalMux I__5497 (
            .O(N__23092),
            .I(N__23055));
    LocalMux I__5496 (
            .O(N__23089),
            .I(N__23055));
    Span4Mux_v I__5495 (
            .O(N__23082),
            .I(N__23046));
    LocalMux I__5494 (
            .O(N__23079),
            .I(N__23046));
    Span4Mux_v I__5493 (
            .O(N__23074),
            .I(N__23046));
    LocalMux I__5492 (
            .O(N__23071),
            .I(N__23046));
    Span12Mux_v I__5491 (
            .O(N__23068),
            .I(N__23043));
    Sp12to4 I__5490 (
            .O(N__23065),
            .I(N__23040));
    Sp12to4 I__5489 (
            .O(N__23062),
            .I(N__23037));
    Span4Mux_v I__5488 (
            .O(N__23055),
            .I(N__23032));
    Span4Mux_v I__5487 (
            .O(N__23046),
            .I(N__23032));
    Span12Mux_h I__5486 (
            .O(N__23043),
            .I(N__23029));
    Span12Mux_h I__5485 (
            .O(N__23040),
            .I(N__23026));
    Span12Mux_h I__5484 (
            .O(N__23037),
            .I(N__23023));
    Span4Mux_v I__5483 (
            .O(N__23032),
            .I(N__23020));
    Odrv12 I__5482 (
            .O(N__23029),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__5481 (
            .O(N__23026),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__5480 (
            .O(N__23023),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__5479 (
            .O(N__23020),
            .I(CONSTANT_ONE_NET));
    InMux I__5478 (
            .O(N__23011),
            .I(N__23008));
    LocalMux I__5477 (
            .O(N__23008),
            .I(N__23005));
    Span4Mux_v I__5476 (
            .O(N__23005),
            .I(N__23002));
    Sp12to4 I__5475 (
            .O(N__23002),
            .I(N__22999));
    Span12Mux_h I__5474 (
            .O(N__22999),
            .I(N__22996));
    Span12Mux_v I__5473 (
            .O(N__22996),
            .I(N__22993));
    Odrv12 I__5472 (
            .O(N__22993),
            .I(\line_buffer.n673 ));
    CascadeMux I__5471 (
            .O(N__22990),
            .I(N__22987));
    InMux I__5470 (
            .O(N__22987),
            .I(N__22984));
    LocalMux I__5469 (
            .O(N__22984),
            .I(N__22981));
    Span4Mux_v I__5468 (
            .O(N__22981),
            .I(N__22978));
    Sp12to4 I__5467 (
            .O(N__22978),
            .I(N__22975));
    Odrv12 I__5466 (
            .O(N__22975),
            .I(\line_buffer.n681 ));
    InMux I__5465 (
            .O(N__22972),
            .I(N__22969));
    LocalMux I__5464 (
            .O(N__22969),
            .I(\line_buffer.n4146 ));
    InMux I__5463 (
            .O(N__22966),
            .I(N__22963));
    LocalMux I__5462 (
            .O(N__22963),
            .I(\line_buffer.n4149 ));
    InMux I__5461 (
            .O(N__22960),
            .I(N__22957));
    LocalMux I__5460 (
            .O(N__22957),
            .I(N__22954));
    Span4Mux_h I__5459 (
            .O(N__22954),
            .I(N__22951));
    Span4Mux_h I__5458 (
            .O(N__22951),
            .I(N__22948));
    Odrv4 I__5457 (
            .O(N__22948),
            .I(TX_DATA_0));
    InMux I__5456 (
            .O(N__22945),
            .I(N__22942));
    LocalMux I__5455 (
            .O(N__22942),
            .I(N__22939));
    Span12Mux_v I__5454 (
            .O(N__22939),
            .I(N__22936));
    Odrv12 I__5453 (
            .O(N__22936),
            .I(\line_buffer.n621 ));
    InMux I__5452 (
            .O(N__22933),
            .I(N__22930));
    LocalMux I__5451 (
            .O(N__22930),
            .I(N__22927));
    Span4Mux_v I__5450 (
            .O(N__22927),
            .I(N__22924));
    Span4Mux_h I__5449 (
            .O(N__22924),
            .I(N__22921));
    Odrv4 I__5448 (
            .O(N__22921),
            .I(\line_buffer.n613 ));
    InMux I__5447 (
            .O(N__22918),
            .I(N__22915));
    LocalMux I__5446 (
            .O(N__22915),
            .I(N__22912));
    Span12Mux_v I__5445 (
            .O(N__22912),
            .I(N__22909));
    Odrv12 I__5444 (
            .O(N__22909),
            .I(\line_buffer.n653 ));
    InMux I__5443 (
            .O(N__22906),
            .I(N__22903));
    LocalMux I__5442 (
            .O(N__22903),
            .I(N__22900));
    Span4Mux_v I__5441 (
            .O(N__22900),
            .I(N__22897));
    Span4Mux_h I__5440 (
            .O(N__22897),
            .I(N__22894));
    Odrv4 I__5439 (
            .O(N__22894),
            .I(\line_buffer.n645 ));
    InMux I__5438 (
            .O(N__22891),
            .I(N__22888));
    LocalMux I__5437 (
            .O(N__22888),
            .I(N__22885));
    Odrv12 I__5436 (
            .O(N__22885),
            .I(\line_buffer.n4062 ));
    InMux I__5435 (
            .O(N__22882),
            .I(N__22879));
    LocalMux I__5434 (
            .O(N__22879),
            .I(N__22876));
    Odrv4 I__5433 (
            .O(N__22876),
            .I(\line_buffer.n4078 ));
    IoInMux I__5432 (
            .O(N__22873),
            .I(N__22870));
    LocalMux I__5431 (
            .O(N__22870),
            .I(N__22866));
    CascadeMux I__5430 (
            .O(N__22869),
            .I(N__22862));
    IoSpan4Mux I__5429 (
            .O(N__22866),
            .I(N__22859));
    InMux I__5428 (
            .O(N__22865),
            .I(N__22853));
    InMux I__5427 (
            .O(N__22862),
            .I(N__22850));
    IoSpan4Mux I__5426 (
            .O(N__22859),
            .I(N__22847));
    CascadeMux I__5425 (
            .O(N__22858),
            .I(N__22843));
    CascadeMux I__5424 (
            .O(N__22857),
            .I(N__22839));
    InMux I__5423 (
            .O(N__22856),
            .I(N__22836));
    LocalMux I__5422 (
            .O(N__22853),
            .I(N__22830));
    LocalMux I__5421 (
            .O(N__22850),
            .I(N__22830));
    Span4Mux_s2_h I__5420 (
            .O(N__22847),
            .I(N__22826));
    InMux I__5419 (
            .O(N__22846),
            .I(N__22823));
    InMux I__5418 (
            .O(N__22843),
            .I(N__22820));
    InMux I__5417 (
            .O(N__22842),
            .I(N__22815));
    InMux I__5416 (
            .O(N__22839),
            .I(N__22812));
    LocalMux I__5415 (
            .O(N__22836),
            .I(N__22809));
    InMux I__5414 (
            .O(N__22835),
            .I(N__22806));
    Span4Mux_v I__5413 (
            .O(N__22830),
            .I(N__22803));
    InMux I__5412 (
            .O(N__22829),
            .I(N__22799));
    Span4Mux_h I__5411 (
            .O(N__22826),
            .I(N__22794));
    LocalMux I__5410 (
            .O(N__22823),
            .I(N__22794));
    LocalMux I__5409 (
            .O(N__22820),
            .I(N__22790));
    InMux I__5408 (
            .O(N__22819),
            .I(N__22787));
    InMux I__5407 (
            .O(N__22818),
            .I(N__22784));
    LocalMux I__5406 (
            .O(N__22815),
            .I(N__22779));
    LocalMux I__5405 (
            .O(N__22812),
            .I(N__22779));
    Span4Mux_v I__5404 (
            .O(N__22809),
            .I(N__22776));
    LocalMux I__5403 (
            .O(N__22806),
            .I(N__22771));
    Span4Mux_v I__5402 (
            .O(N__22803),
            .I(N__22771));
    InMux I__5401 (
            .O(N__22802),
            .I(N__22768));
    LocalMux I__5400 (
            .O(N__22799),
            .I(N__22765));
    Span4Mux_h I__5399 (
            .O(N__22794),
            .I(N__22761));
    InMux I__5398 (
            .O(N__22793),
            .I(N__22758));
    Span4Mux_v I__5397 (
            .O(N__22790),
            .I(N__22755));
    LocalMux I__5396 (
            .O(N__22787),
            .I(N__22748));
    LocalMux I__5395 (
            .O(N__22784),
            .I(N__22748));
    Span4Mux_v I__5394 (
            .O(N__22779),
            .I(N__22748));
    Span4Mux_v I__5393 (
            .O(N__22776),
            .I(N__22741));
    Span4Mux_h I__5392 (
            .O(N__22771),
            .I(N__22741));
    LocalMux I__5391 (
            .O(N__22768),
            .I(N__22741));
    Span4Mux_h I__5390 (
            .O(N__22765),
            .I(N__22738));
    InMux I__5389 (
            .O(N__22764),
            .I(N__22735));
    Span4Mux_v I__5388 (
            .O(N__22761),
            .I(N__22726));
    LocalMux I__5387 (
            .O(N__22758),
            .I(N__22726));
    Span4Mux_v I__5386 (
            .O(N__22755),
            .I(N__22726));
    Span4Mux_h I__5385 (
            .O(N__22748),
            .I(N__22726));
    Span4Mux_h I__5384 (
            .O(N__22741),
            .I(N__22723));
    Odrv4 I__5383 (
            .O(N__22738),
            .I(DEBUG_c_2));
    LocalMux I__5382 (
            .O(N__22735),
            .I(DEBUG_c_2));
    Odrv4 I__5381 (
            .O(N__22726),
            .I(DEBUG_c_2));
    Odrv4 I__5380 (
            .O(N__22723),
            .I(DEBUG_c_2));
    InMux I__5379 (
            .O(N__22714),
            .I(N__22711));
    LocalMux I__5378 (
            .O(N__22711),
            .I(\line_buffer.n4140 ));
    InMux I__5377 (
            .O(N__22708),
            .I(N__22705));
    LocalMux I__5376 (
            .O(N__22705),
            .I(N__22702));
    Span4Mux_h I__5375 (
            .O(N__22702),
            .I(N__22699));
    Span4Mux_h I__5374 (
            .O(N__22699),
            .I(N__22696));
    Span4Mux_v I__5373 (
            .O(N__22696),
            .I(N__22693));
    Odrv4 I__5372 (
            .O(N__22693),
            .I(TX_DATA_4));
    ClkMux I__5371 (
            .O(N__22690),
            .I(N__22685));
    ClkMux I__5370 (
            .O(N__22689),
            .I(N__22681));
    ClkMux I__5369 (
            .O(N__22688),
            .I(N__22678));
    LocalMux I__5368 (
            .O(N__22685),
            .I(N__22672));
    ClkMux I__5367 (
            .O(N__22684),
            .I(N__22669));
    LocalMux I__5366 (
            .O(N__22681),
            .I(N__22665));
    LocalMux I__5365 (
            .O(N__22678),
            .I(N__22662));
    ClkMux I__5364 (
            .O(N__22677),
            .I(N__22659));
    ClkMux I__5363 (
            .O(N__22676),
            .I(N__22656));
    ClkMux I__5362 (
            .O(N__22675),
            .I(N__22651));
    Span4Mux_s2_v I__5361 (
            .O(N__22672),
            .I(N__22644));
    LocalMux I__5360 (
            .O(N__22669),
            .I(N__22644));
    ClkMux I__5359 (
            .O(N__22668),
            .I(N__22641));
    Span4Mux_s2_v I__5358 (
            .O(N__22665),
            .I(N__22633));
    Span4Mux_h I__5357 (
            .O(N__22662),
            .I(N__22633));
    LocalMux I__5356 (
            .O(N__22659),
            .I(N__22633));
    LocalMux I__5355 (
            .O(N__22656),
            .I(N__22630));
    ClkMux I__5354 (
            .O(N__22655),
            .I(N__22627));
    ClkMux I__5353 (
            .O(N__22654),
            .I(N__22624));
    LocalMux I__5352 (
            .O(N__22651),
            .I(N__22616));
    ClkMux I__5351 (
            .O(N__22650),
            .I(N__22613));
    ClkMux I__5350 (
            .O(N__22649),
            .I(N__22610));
    Span4Mux_v I__5349 (
            .O(N__22644),
            .I(N__22604));
    LocalMux I__5348 (
            .O(N__22641),
            .I(N__22604));
    ClkMux I__5347 (
            .O(N__22640),
            .I(N__22601));
    Span4Mux_v I__5346 (
            .O(N__22633),
            .I(N__22593));
    Span4Mux_h I__5345 (
            .O(N__22630),
            .I(N__22593));
    LocalMux I__5344 (
            .O(N__22627),
            .I(N__22593));
    LocalMux I__5343 (
            .O(N__22624),
            .I(N__22590));
    ClkMux I__5342 (
            .O(N__22623),
            .I(N__22587));
    ClkMux I__5341 (
            .O(N__22622),
            .I(N__22584));
    ClkMux I__5340 (
            .O(N__22621),
            .I(N__22575));
    ClkMux I__5339 (
            .O(N__22620),
            .I(N__22569));
    ClkMux I__5338 (
            .O(N__22619),
            .I(N__22566));
    Span4Mux_v I__5337 (
            .O(N__22616),
            .I(N__22555));
    LocalMux I__5336 (
            .O(N__22613),
            .I(N__22555));
    LocalMux I__5335 (
            .O(N__22610),
            .I(N__22552));
    ClkMux I__5334 (
            .O(N__22609),
            .I(N__22549));
    Span4Mux_h I__5333 (
            .O(N__22604),
            .I(N__22542));
    LocalMux I__5332 (
            .O(N__22601),
            .I(N__22542));
    ClkMux I__5331 (
            .O(N__22600),
            .I(N__22539));
    Span4Mux_v I__5330 (
            .O(N__22593),
            .I(N__22526));
    Span4Mux_h I__5329 (
            .O(N__22590),
            .I(N__22526));
    LocalMux I__5328 (
            .O(N__22587),
            .I(N__22526));
    LocalMux I__5327 (
            .O(N__22584),
            .I(N__22523));
    ClkMux I__5326 (
            .O(N__22583),
            .I(N__22520));
    ClkMux I__5325 (
            .O(N__22582),
            .I(N__22517));
    ClkMux I__5324 (
            .O(N__22581),
            .I(N__22509));
    ClkMux I__5323 (
            .O(N__22580),
            .I(N__22506));
    ClkMux I__5322 (
            .O(N__22579),
            .I(N__22503));
    ClkMux I__5321 (
            .O(N__22578),
            .I(N__22500));
    LocalMux I__5320 (
            .O(N__22575),
            .I(N__22495));
    ClkMux I__5319 (
            .O(N__22574),
            .I(N__22492));
    ClkMux I__5318 (
            .O(N__22573),
            .I(N__22489));
    ClkMux I__5317 (
            .O(N__22572),
            .I(N__22483));
    LocalMux I__5316 (
            .O(N__22569),
            .I(N__22478));
    LocalMux I__5315 (
            .O(N__22566),
            .I(N__22478));
    ClkMux I__5314 (
            .O(N__22565),
            .I(N__22475));
    ClkMux I__5313 (
            .O(N__22564),
            .I(N__22471));
    ClkMux I__5312 (
            .O(N__22563),
            .I(N__22467));
    ClkMux I__5311 (
            .O(N__22562),
            .I(N__22462));
    ClkMux I__5310 (
            .O(N__22561),
            .I(N__22459));
    ClkMux I__5309 (
            .O(N__22560),
            .I(N__22456));
    Span4Mux_h I__5308 (
            .O(N__22555),
            .I(N__22449));
    Span4Mux_h I__5307 (
            .O(N__22552),
            .I(N__22449));
    LocalMux I__5306 (
            .O(N__22549),
            .I(N__22449));
    ClkMux I__5305 (
            .O(N__22548),
            .I(N__22446));
    ClkMux I__5304 (
            .O(N__22547),
            .I(N__22441));
    Span4Mux_v I__5303 (
            .O(N__22542),
            .I(N__22429));
    LocalMux I__5302 (
            .O(N__22539),
            .I(N__22429));
    ClkMux I__5301 (
            .O(N__22538),
            .I(N__22426));
    ClkMux I__5300 (
            .O(N__22537),
            .I(N__22423));
    IoInMux I__5299 (
            .O(N__22536),
            .I(N__22416));
    ClkMux I__5298 (
            .O(N__22535),
            .I(N__22413));
    ClkMux I__5297 (
            .O(N__22534),
            .I(N__22410));
    ClkMux I__5296 (
            .O(N__22533),
            .I(N__22404));
    Span4Mux_v I__5295 (
            .O(N__22526),
            .I(N__22397));
    Span4Mux_h I__5294 (
            .O(N__22523),
            .I(N__22397));
    LocalMux I__5293 (
            .O(N__22520),
            .I(N__22397));
    LocalMux I__5292 (
            .O(N__22517),
            .I(N__22394));
    ClkMux I__5291 (
            .O(N__22516),
            .I(N__22391));
    ClkMux I__5290 (
            .O(N__22515),
            .I(N__22388));
    ClkMux I__5289 (
            .O(N__22514),
            .I(N__22383));
    ClkMux I__5288 (
            .O(N__22513),
            .I(N__22380));
    ClkMux I__5287 (
            .O(N__22512),
            .I(N__22377));
    LocalMux I__5286 (
            .O(N__22509),
            .I(N__22374));
    LocalMux I__5285 (
            .O(N__22506),
            .I(N__22371));
    LocalMux I__5284 (
            .O(N__22503),
            .I(N__22366));
    LocalMux I__5283 (
            .O(N__22500),
            .I(N__22366));
    ClkMux I__5282 (
            .O(N__22499),
            .I(N__22363));
    ClkMux I__5281 (
            .O(N__22498),
            .I(N__22360));
    Span4Mux_v I__5280 (
            .O(N__22495),
            .I(N__22353));
    LocalMux I__5279 (
            .O(N__22492),
            .I(N__22353));
    LocalMux I__5278 (
            .O(N__22489),
            .I(N__22353));
    ClkMux I__5277 (
            .O(N__22488),
            .I(N__22349));
    ClkMux I__5276 (
            .O(N__22487),
            .I(N__22344));
    ClkMux I__5275 (
            .O(N__22486),
            .I(N__22341));
    LocalMux I__5274 (
            .O(N__22483),
            .I(N__22337));
    Span4Mux_h I__5273 (
            .O(N__22478),
            .I(N__22332));
    LocalMux I__5272 (
            .O(N__22475),
            .I(N__22332));
    ClkMux I__5271 (
            .O(N__22474),
            .I(N__22329));
    LocalMux I__5270 (
            .O(N__22471),
            .I(N__22326));
    ClkMux I__5269 (
            .O(N__22470),
            .I(N__22323));
    LocalMux I__5268 (
            .O(N__22467),
            .I(N__22319));
    ClkMux I__5267 (
            .O(N__22466),
            .I(N__22316));
    ClkMux I__5266 (
            .O(N__22465),
            .I(N__22311));
    LocalMux I__5265 (
            .O(N__22462),
            .I(N__22308));
    LocalMux I__5264 (
            .O(N__22459),
            .I(N__22303));
    LocalMux I__5263 (
            .O(N__22456),
            .I(N__22303));
    Span4Mux_h I__5262 (
            .O(N__22449),
            .I(N__22298));
    LocalMux I__5261 (
            .O(N__22446),
            .I(N__22298));
    ClkMux I__5260 (
            .O(N__22445),
            .I(N__22295));
    ClkMux I__5259 (
            .O(N__22444),
            .I(N__22292));
    LocalMux I__5258 (
            .O(N__22441),
            .I(N__22289));
    ClkMux I__5257 (
            .O(N__22440),
            .I(N__22286));
    ClkMux I__5256 (
            .O(N__22439),
            .I(N__22283));
    ClkMux I__5255 (
            .O(N__22438),
            .I(N__22279));
    ClkMux I__5254 (
            .O(N__22437),
            .I(N__22276));
    ClkMux I__5253 (
            .O(N__22436),
            .I(N__22273));
    ClkMux I__5252 (
            .O(N__22435),
            .I(N__22270));
    ClkMux I__5251 (
            .O(N__22434),
            .I(N__22267));
    Span4Mux_h I__5250 (
            .O(N__22429),
            .I(N__22263));
    LocalMux I__5249 (
            .O(N__22426),
            .I(N__22258));
    LocalMux I__5248 (
            .O(N__22423),
            .I(N__22258));
    ClkMux I__5247 (
            .O(N__22422),
            .I(N__22255));
    ClkMux I__5246 (
            .O(N__22421),
            .I(N__22252));
    ClkMux I__5245 (
            .O(N__22420),
            .I(N__22249));
    ClkMux I__5244 (
            .O(N__22419),
            .I(N__22244));
    LocalMux I__5243 (
            .O(N__22416),
            .I(N__22240));
    LocalMux I__5242 (
            .O(N__22413),
            .I(N__22234));
    LocalMux I__5241 (
            .O(N__22410),
            .I(N__22234));
    ClkMux I__5240 (
            .O(N__22409),
            .I(N__22231));
    ClkMux I__5239 (
            .O(N__22408),
            .I(N__22226));
    ClkMux I__5238 (
            .O(N__22407),
            .I(N__22222));
    LocalMux I__5237 (
            .O(N__22404),
            .I(N__22219));
    Span4Mux_v I__5236 (
            .O(N__22397),
            .I(N__22212));
    Span4Mux_h I__5235 (
            .O(N__22394),
            .I(N__22212));
    LocalMux I__5234 (
            .O(N__22391),
            .I(N__22212));
    LocalMux I__5233 (
            .O(N__22388),
            .I(N__22209));
    ClkMux I__5232 (
            .O(N__22387),
            .I(N__22206));
    ClkMux I__5231 (
            .O(N__22386),
            .I(N__22202));
    LocalMux I__5230 (
            .O(N__22383),
            .I(N__22199));
    LocalMux I__5229 (
            .O(N__22380),
            .I(N__22196));
    LocalMux I__5228 (
            .O(N__22377),
            .I(N__22193));
    Span4Mux_h I__5227 (
            .O(N__22374),
            .I(N__22180));
    Span4Mux_v I__5226 (
            .O(N__22371),
            .I(N__22180));
    Span4Mux_h I__5225 (
            .O(N__22366),
            .I(N__22180));
    LocalMux I__5224 (
            .O(N__22363),
            .I(N__22180));
    LocalMux I__5223 (
            .O(N__22360),
            .I(N__22180));
    Span4Mux_h I__5222 (
            .O(N__22353),
            .I(N__22180));
    ClkMux I__5221 (
            .O(N__22352),
            .I(N__22177));
    LocalMux I__5220 (
            .O(N__22349),
            .I(N__22174));
    ClkMux I__5219 (
            .O(N__22348),
            .I(N__22171));
    ClkMux I__5218 (
            .O(N__22347),
            .I(N__22168));
    LocalMux I__5217 (
            .O(N__22344),
            .I(N__22165));
    LocalMux I__5216 (
            .O(N__22341),
            .I(N__22162));
    ClkMux I__5215 (
            .O(N__22340),
            .I(N__22159));
    Span4Mux_h I__5214 (
            .O(N__22337),
            .I(N__22154));
    Span4Mux_h I__5213 (
            .O(N__22332),
            .I(N__22154));
    LocalMux I__5212 (
            .O(N__22329),
            .I(N__22151));
    Span4Mux_h I__5211 (
            .O(N__22326),
            .I(N__22146));
    LocalMux I__5210 (
            .O(N__22323),
            .I(N__22146));
    ClkMux I__5209 (
            .O(N__22322),
            .I(N__22143));
    Span4Mux_h I__5208 (
            .O(N__22319),
            .I(N__22140));
    LocalMux I__5207 (
            .O(N__22316),
            .I(N__22137));
    ClkMux I__5206 (
            .O(N__22315),
            .I(N__22134));
    ClkMux I__5205 (
            .O(N__22314),
            .I(N__22131));
    LocalMux I__5204 (
            .O(N__22311),
            .I(N__22128));
    Span4Mux_h I__5203 (
            .O(N__22308),
            .I(N__22117));
    Span4Mux_h I__5202 (
            .O(N__22303),
            .I(N__22117));
    Span4Mux_h I__5201 (
            .O(N__22298),
            .I(N__22117));
    LocalMux I__5200 (
            .O(N__22295),
            .I(N__22117));
    LocalMux I__5199 (
            .O(N__22292),
            .I(N__22117));
    Span4Mux_h I__5198 (
            .O(N__22289),
            .I(N__22112));
    LocalMux I__5197 (
            .O(N__22286),
            .I(N__22112));
    LocalMux I__5196 (
            .O(N__22283),
            .I(N__22109));
    ClkMux I__5195 (
            .O(N__22282),
            .I(N__22106));
    LocalMux I__5194 (
            .O(N__22279),
            .I(N__22101));
    LocalMux I__5193 (
            .O(N__22276),
            .I(N__22101));
    LocalMux I__5192 (
            .O(N__22273),
            .I(N__22096));
    LocalMux I__5191 (
            .O(N__22270),
            .I(N__22096));
    LocalMux I__5190 (
            .O(N__22267),
            .I(N__22093));
    ClkMux I__5189 (
            .O(N__22266),
            .I(N__22090));
    Span4Mux_v I__5188 (
            .O(N__22263),
            .I(N__22083));
    Span4Mux_h I__5187 (
            .O(N__22258),
            .I(N__22083));
    LocalMux I__5186 (
            .O(N__22255),
            .I(N__22083));
    LocalMux I__5185 (
            .O(N__22252),
            .I(N__22080));
    LocalMux I__5184 (
            .O(N__22249),
            .I(N__22077));
    ClkMux I__5183 (
            .O(N__22248),
            .I(N__22074));
    ClkMux I__5182 (
            .O(N__22247),
            .I(N__22071));
    LocalMux I__5181 (
            .O(N__22244),
            .I(N__22066));
    ClkMux I__5180 (
            .O(N__22243),
            .I(N__22063));
    IoSpan4Mux I__5179 (
            .O(N__22240),
            .I(N__22058));
    ClkMux I__5178 (
            .O(N__22239),
            .I(N__22055));
    Span4Mux_v I__5177 (
            .O(N__22234),
            .I(N__22050));
    LocalMux I__5176 (
            .O(N__22231),
            .I(N__22050));
    ClkMux I__5175 (
            .O(N__22230),
            .I(N__22047));
    ClkMux I__5174 (
            .O(N__22229),
            .I(N__22044));
    LocalMux I__5173 (
            .O(N__22226),
            .I(N__22041));
    ClkMux I__5172 (
            .O(N__22225),
            .I(N__22038));
    LocalMux I__5171 (
            .O(N__22222),
            .I(N__22034));
    Span4Mux_v I__5170 (
            .O(N__22219),
            .I(N__22031));
    Span4Mux_v I__5169 (
            .O(N__22212),
            .I(N__22024));
    Span4Mux_h I__5168 (
            .O(N__22209),
            .I(N__22024));
    LocalMux I__5167 (
            .O(N__22206),
            .I(N__22024));
    ClkMux I__5166 (
            .O(N__22205),
            .I(N__22021));
    LocalMux I__5165 (
            .O(N__22202),
            .I(N__22017));
    Span4Mux_v I__5164 (
            .O(N__22199),
            .I(N__22006));
    Span4Mux_v I__5163 (
            .O(N__22196),
            .I(N__22006));
    Span4Mux_h I__5162 (
            .O(N__22193),
            .I(N__22006));
    Span4Mux_h I__5161 (
            .O(N__22180),
            .I(N__22006));
    LocalMux I__5160 (
            .O(N__22177),
            .I(N__22006));
    Span4Mux_h I__5159 (
            .O(N__22174),
            .I(N__21999));
    LocalMux I__5158 (
            .O(N__22171),
            .I(N__21999));
    LocalMux I__5157 (
            .O(N__22168),
            .I(N__21999));
    Span4Mux_v I__5156 (
            .O(N__22165),
            .I(N__21992));
    Span4Mux_h I__5155 (
            .O(N__22162),
            .I(N__21992));
    LocalMux I__5154 (
            .O(N__22159),
            .I(N__21992));
    Span4Mux_v I__5153 (
            .O(N__22154),
            .I(N__21985));
    Span4Mux_h I__5152 (
            .O(N__22151),
            .I(N__21985));
    Span4Mux_h I__5151 (
            .O(N__22146),
            .I(N__21985));
    LocalMux I__5150 (
            .O(N__22143),
            .I(N__21982));
    Span4Mux_h I__5149 (
            .O(N__22140),
            .I(N__21977));
    Span4Mux_h I__5148 (
            .O(N__22137),
            .I(N__21977));
    LocalMux I__5147 (
            .O(N__22134),
            .I(N__21972));
    LocalMux I__5146 (
            .O(N__22131),
            .I(N__21972));
    Span4Mux_h I__5145 (
            .O(N__22128),
            .I(N__21965));
    Span4Mux_v I__5144 (
            .O(N__22117),
            .I(N__21965));
    Span4Mux_h I__5143 (
            .O(N__22112),
            .I(N__21965));
    Span4Mux_v I__5142 (
            .O(N__22109),
            .I(N__21960));
    LocalMux I__5141 (
            .O(N__22106),
            .I(N__21960));
    Span4Mux_v I__5140 (
            .O(N__22101),
            .I(N__21949));
    Span4Mux_h I__5139 (
            .O(N__22096),
            .I(N__21949));
    Span4Mux_h I__5138 (
            .O(N__22093),
            .I(N__21949));
    LocalMux I__5137 (
            .O(N__22090),
            .I(N__21949));
    Span4Mux_h I__5136 (
            .O(N__22083),
            .I(N__21938));
    Span4Mux_v I__5135 (
            .O(N__22080),
            .I(N__21938));
    Span4Mux_h I__5134 (
            .O(N__22077),
            .I(N__21938));
    LocalMux I__5133 (
            .O(N__22074),
            .I(N__21938));
    LocalMux I__5132 (
            .O(N__22071),
            .I(N__21938));
    ClkMux I__5131 (
            .O(N__22070),
            .I(N__21935));
    ClkMux I__5130 (
            .O(N__22069),
            .I(N__21932));
    Span4Mux_h I__5129 (
            .O(N__22066),
            .I(N__21927));
    LocalMux I__5128 (
            .O(N__22063),
            .I(N__21927));
    ClkMux I__5127 (
            .O(N__22062),
            .I(N__21924));
    ClkMux I__5126 (
            .O(N__22061),
            .I(N__21921));
    Span4Mux_s1_v I__5125 (
            .O(N__22058),
            .I(N__21918));
    LocalMux I__5124 (
            .O(N__22055),
            .I(N__21915));
    Span4Mux_h I__5123 (
            .O(N__22050),
            .I(N__21908));
    LocalMux I__5122 (
            .O(N__22047),
            .I(N__21908));
    LocalMux I__5121 (
            .O(N__22044),
            .I(N__21908));
    Span4Mux_v I__5120 (
            .O(N__22041),
            .I(N__21903));
    LocalMux I__5119 (
            .O(N__22038),
            .I(N__21903));
    ClkMux I__5118 (
            .O(N__22037),
            .I(N__21900));
    Span12Mux_h I__5117 (
            .O(N__22034),
            .I(N__21897));
    Sp12to4 I__5116 (
            .O(N__22031),
            .I(N__21894));
    Span4Mux_v I__5115 (
            .O(N__22024),
            .I(N__21891));
    LocalMux I__5114 (
            .O(N__22021),
            .I(N__21888));
    ClkMux I__5113 (
            .O(N__22020),
            .I(N__21885));
    Span4Mux_h I__5112 (
            .O(N__22017),
            .I(N__21882));
    Span4Mux_v I__5111 (
            .O(N__22006),
            .I(N__21875));
    Span4Mux_h I__5110 (
            .O(N__21999),
            .I(N__21875));
    Span4Mux_h I__5109 (
            .O(N__21992),
            .I(N__21875));
    Span4Mux_v I__5108 (
            .O(N__21985),
            .I(N__21870));
    Span4Mux_h I__5107 (
            .O(N__21982),
            .I(N__21870));
    Span4Mux_v I__5106 (
            .O(N__21977),
            .I(N__21865));
    Span4Mux_h I__5105 (
            .O(N__21972),
            .I(N__21865));
    Span4Mux_v I__5104 (
            .O(N__21965),
            .I(N__21860));
    Span4Mux_h I__5103 (
            .O(N__21960),
            .I(N__21860));
    ClkMux I__5102 (
            .O(N__21959),
            .I(N__21857));
    ClkMux I__5101 (
            .O(N__21958),
            .I(N__21854));
    Span4Mux_h I__5100 (
            .O(N__21949),
            .I(N__21845));
    Span4Mux_v I__5099 (
            .O(N__21938),
            .I(N__21845));
    LocalMux I__5098 (
            .O(N__21935),
            .I(N__21845));
    LocalMux I__5097 (
            .O(N__21932),
            .I(N__21845));
    Span4Mux_v I__5096 (
            .O(N__21927),
            .I(N__21838));
    LocalMux I__5095 (
            .O(N__21924),
            .I(N__21838));
    LocalMux I__5094 (
            .O(N__21921),
            .I(N__21838));
    Span4Mux_h I__5093 (
            .O(N__21918),
            .I(N__21833));
    Span4Mux_h I__5092 (
            .O(N__21915),
            .I(N__21833));
    Span4Mux_v I__5091 (
            .O(N__21908),
            .I(N__21830));
    Span4Mux_v I__5090 (
            .O(N__21903),
            .I(N__21825));
    LocalMux I__5089 (
            .O(N__21900),
            .I(N__21825));
    Span12Mux_v I__5088 (
            .O(N__21897),
            .I(N__21820));
    Span12Mux_h I__5087 (
            .O(N__21894),
            .I(N__21820));
    Sp12to4 I__5086 (
            .O(N__21891),
            .I(N__21815));
    Sp12to4 I__5085 (
            .O(N__21888),
            .I(N__21815));
    LocalMux I__5084 (
            .O(N__21885),
            .I(N__21812));
    Span4Mux_h I__5083 (
            .O(N__21882),
            .I(N__21809));
    Span4Mux_v I__5082 (
            .O(N__21875),
            .I(N__21806));
    Span4Mux_v I__5081 (
            .O(N__21870),
            .I(N__21801));
    Span4Mux_v I__5080 (
            .O(N__21865),
            .I(N__21801));
    Span4Mux_v I__5079 (
            .O(N__21860),
            .I(N__21798));
    LocalMux I__5078 (
            .O(N__21857),
            .I(N__21793));
    LocalMux I__5077 (
            .O(N__21854),
            .I(N__21793));
    Span4Mux_v I__5076 (
            .O(N__21845),
            .I(N__21788));
    Span4Mux_v I__5075 (
            .O(N__21838),
            .I(N__21788));
    Span4Mux_h I__5074 (
            .O(N__21833),
            .I(N__21785));
    Span4Mux_v I__5073 (
            .O(N__21830),
            .I(N__21780));
    Span4Mux_h I__5072 (
            .O(N__21825),
            .I(N__21780));
    Span12Mux_v I__5071 (
            .O(N__21820),
            .I(N__21773));
    Span12Mux_h I__5070 (
            .O(N__21815),
            .I(N__21773));
    Span12Mux_h I__5069 (
            .O(N__21812),
            .I(N__21773));
    Span4Mux_h I__5068 (
            .O(N__21809),
            .I(N__21768));
    Span4Mux_v I__5067 (
            .O(N__21806),
            .I(N__21768));
    Span4Mux_v I__5066 (
            .O(N__21801),
            .I(N__21765));
    Span4Mux_v I__5065 (
            .O(N__21798),
            .I(N__21762));
    Span12Mux_h I__5064 (
            .O(N__21793),
            .I(N__21757));
    Sp12to4 I__5063 (
            .O(N__21788),
            .I(N__21757));
    Span4Mux_h I__5062 (
            .O(N__21785),
            .I(N__21752));
    Span4Mux_h I__5061 (
            .O(N__21780),
            .I(N__21752));
    Odrv12 I__5060 (
            .O(N__21773),
            .I(ADV_CLK_c));
    Odrv4 I__5059 (
            .O(N__21768),
            .I(ADV_CLK_c));
    Odrv4 I__5058 (
            .O(N__21765),
            .I(ADV_CLK_c));
    Odrv4 I__5057 (
            .O(N__21762),
            .I(ADV_CLK_c));
    Odrv12 I__5056 (
            .O(N__21757),
            .I(ADV_CLK_c));
    Odrv4 I__5055 (
            .O(N__21752),
            .I(ADV_CLK_c));
    InMux I__5054 (
            .O(N__21739),
            .I(N__21736));
    LocalMux I__5053 (
            .O(N__21736),
            .I(N__21733));
    Span4Mux_h I__5052 (
            .O(N__21733),
            .I(N__21730));
    Span4Mux_h I__5051 (
            .O(N__21730),
            .I(N__21727));
    Odrv4 I__5050 (
            .O(N__21727),
            .I(\line_buffer.n641 ));
    CascadeMux I__5049 (
            .O(N__21724),
            .I(N__21721));
    InMux I__5048 (
            .O(N__21721),
            .I(N__21718));
    LocalMux I__5047 (
            .O(N__21718),
            .I(N__21715));
    Span12Mux_v I__5046 (
            .O(N__21715),
            .I(N__21712));
    Odrv12 I__5045 (
            .O(N__21712),
            .I(\line_buffer.n649 ));
    InMux I__5044 (
            .O(N__21709),
            .I(N__21706));
    LocalMux I__5043 (
            .O(N__21706),
            .I(N__21703));
    Span4Mux_v I__5042 (
            .O(N__21703),
            .I(N__21700));
    Span4Mux_h I__5041 (
            .O(N__21700),
            .I(N__21697));
    Odrv4 I__5040 (
            .O(N__21697),
            .I(\line_buffer.n552 ));
    InMux I__5039 (
            .O(N__21694),
            .I(N__21691));
    LocalMux I__5038 (
            .O(N__21691),
            .I(\line_buffer.n4116 ));
    CascadeMux I__5037 (
            .O(N__21688),
            .I(N__21685));
    InMux I__5036 (
            .O(N__21685),
            .I(N__21682));
    LocalMux I__5035 (
            .O(N__21682),
            .I(N__21679));
    Span12Mux_h I__5034 (
            .O(N__21679),
            .I(N__21676));
    Span12Mux_v I__5033 (
            .O(N__21676),
            .I(N__21673));
    Odrv12 I__5032 (
            .O(N__21673),
            .I(\line_buffer.n544 ));
    InMux I__5031 (
            .O(N__21670),
            .I(N__21667));
    LocalMux I__5030 (
            .O(N__21667),
            .I(\line_buffer.n4119 ));
    InMux I__5029 (
            .O(N__21664),
            .I(N__21661));
    LocalMux I__5028 (
            .O(N__21661),
            .I(N__21658));
    Span4Mux_h I__5027 (
            .O(N__21658),
            .I(N__21655));
    Span4Mux_h I__5026 (
            .O(N__21655),
            .I(N__21652));
    Span4Mux_h I__5025 (
            .O(N__21652),
            .I(N__21649));
    Odrv4 I__5024 (
            .O(N__21649),
            .I(\line_buffer.n684 ));
    InMux I__5023 (
            .O(N__21646),
            .I(N__21643));
    LocalMux I__5022 (
            .O(N__21643),
            .I(N__21640));
    Span4Mux_v I__5021 (
            .O(N__21640),
            .I(N__21637));
    Sp12to4 I__5020 (
            .O(N__21637),
            .I(N__21634));
    Span12Mux_h I__5019 (
            .O(N__21634),
            .I(N__21631));
    Odrv12 I__5018 (
            .O(N__21631),
            .I(\line_buffer.n676 ));
    InMux I__5017 (
            .O(N__21628),
            .I(N__21625));
    LocalMux I__5016 (
            .O(N__21625),
            .I(\line_buffer.n4066 ));
    InMux I__5015 (
            .O(N__21622),
            .I(N__21619));
    LocalMux I__5014 (
            .O(N__21619),
            .I(N__21616));
    Span4Mux_h I__5013 (
            .O(N__21616),
            .I(N__21613));
    Span4Mux_h I__5012 (
            .O(N__21613),
            .I(N__21610));
    Odrv4 I__5011 (
            .O(N__21610),
            .I(\line_buffer.n555 ));
    InMux I__5010 (
            .O(N__21607),
            .I(N__21604));
    LocalMux I__5009 (
            .O(N__21604),
            .I(N__21601));
    Span4Mux_v I__5008 (
            .O(N__21601),
            .I(N__21598));
    Sp12to4 I__5007 (
            .O(N__21598),
            .I(N__21595));
    Span12Mux_h I__5006 (
            .O(N__21595),
            .I(N__21592));
    Odrv12 I__5005 (
            .O(N__21592),
            .I(\line_buffer.n547 ));
    CascadeMux I__5004 (
            .O(N__21589),
            .I(\line_buffer.n4074_cascade_ ));
    InMux I__5003 (
            .O(N__21586),
            .I(N__21583));
    LocalMux I__5002 (
            .O(N__21583),
            .I(\line_buffer.n4128 ));
    InMux I__5001 (
            .O(N__21580),
            .I(N__21577));
    LocalMux I__5000 (
            .O(N__21577),
            .I(N__21574));
    Odrv12 I__4999 (
            .O(N__21574),
            .I(TX_DATA_3));
    InMux I__4998 (
            .O(N__21571),
            .I(N__21568));
    LocalMux I__4997 (
            .O(N__21568),
            .I(N__21565));
    Span4Mux_h I__4996 (
            .O(N__21565),
            .I(N__21562));
    Span4Mux_h I__4995 (
            .O(N__21562),
            .I(N__21559));
    Span4Mux_h I__4994 (
            .O(N__21559),
            .I(N__21556));
    Span4Mux_v I__4993 (
            .O(N__21556),
            .I(N__21553));
    Span4Mux_v I__4992 (
            .O(N__21553),
            .I(N__21550));
    Odrv4 I__4991 (
            .O(N__21550),
            .I(\line_buffer.n652 ));
    InMux I__4990 (
            .O(N__21547),
            .I(N__21544));
    LocalMux I__4989 (
            .O(N__21544),
            .I(N__21541));
    Span4Mux_v I__4988 (
            .O(N__21541),
            .I(N__21538));
    Span4Mux_h I__4987 (
            .O(N__21538),
            .I(N__21535));
    Span4Mux_h I__4986 (
            .O(N__21535),
            .I(N__21532));
    Odrv4 I__4985 (
            .O(N__21532),
            .I(\line_buffer.n644 ));
    InMux I__4984 (
            .O(N__21529),
            .I(N__21526));
    LocalMux I__4983 (
            .O(N__21526),
            .I(\line_buffer.n4075 ));
    InMux I__4982 (
            .O(N__21523),
            .I(N__21520));
    LocalMux I__4981 (
            .O(N__21520),
            .I(N__21517));
    Span4Mux_v I__4980 (
            .O(N__21517),
            .I(N__21514));
    Odrv4 I__4979 (
            .O(N__21514),
            .I(\transmit_module.Y_DELTA_PATTERN_33 ));
    InMux I__4978 (
            .O(N__21511),
            .I(N__21508));
    LocalMux I__4977 (
            .O(N__21508),
            .I(N__21505));
    Span4Mux_v I__4976 (
            .O(N__21505),
            .I(N__21502));
    Odrv4 I__4975 (
            .O(N__21502),
            .I(\transmit_module.Y_DELTA_PATTERN_35 ));
    InMux I__4974 (
            .O(N__21499),
            .I(N__21496));
    LocalMux I__4973 (
            .O(N__21496),
            .I(\transmit_module.Y_DELTA_PATTERN_34 ));
    CEMux I__4972 (
            .O(N__21493),
            .I(N__21490));
    LocalMux I__4971 (
            .O(N__21490),
            .I(N__21484));
    CEMux I__4970 (
            .O(N__21489),
            .I(N__21481));
    CEMux I__4969 (
            .O(N__21488),
            .I(N__21477));
    CEMux I__4968 (
            .O(N__21487),
            .I(N__21474));
    Span4Mux_h I__4967 (
            .O(N__21484),
            .I(N__21468));
    LocalMux I__4966 (
            .O(N__21481),
            .I(N__21468));
    CEMux I__4965 (
            .O(N__21480),
            .I(N__21465));
    LocalMux I__4964 (
            .O(N__21477),
            .I(N__21460));
    LocalMux I__4963 (
            .O(N__21474),
            .I(N__21453));
    CEMux I__4962 (
            .O(N__21473),
            .I(N__21450));
    Span4Mux_v I__4961 (
            .O(N__21468),
            .I(N__21447));
    LocalMux I__4960 (
            .O(N__21465),
            .I(N__21444));
    CEMux I__4959 (
            .O(N__21464),
            .I(N__21441));
    CEMux I__4958 (
            .O(N__21463),
            .I(N__21438));
    Span4Mux_h I__4957 (
            .O(N__21460),
            .I(N__21433));
    CEMux I__4956 (
            .O(N__21459),
            .I(N__21430));
    CEMux I__4955 (
            .O(N__21458),
            .I(N__21427));
    CEMux I__4954 (
            .O(N__21457),
            .I(N__21424));
    CEMux I__4953 (
            .O(N__21456),
            .I(N__21421));
    Span4Mux_v I__4952 (
            .O(N__21453),
            .I(N__21416));
    LocalMux I__4951 (
            .O(N__21450),
            .I(N__21416));
    Span4Mux_h I__4950 (
            .O(N__21447),
            .I(N__21409));
    Span4Mux_h I__4949 (
            .O(N__21444),
            .I(N__21409));
    LocalMux I__4948 (
            .O(N__21441),
            .I(N__21409));
    LocalMux I__4947 (
            .O(N__21438),
            .I(N__21406));
    CEMux I__4946 (
            .O(N__21437),
            .I(N__21403));
    CEMux I__4945 (
            .O(N__21436),
            .I(N__21400));
    Span4Mux_v I__4944 (
            .O(N__21433),
            .I(N__21395));
    LocalMux I__4943 (
            .O(N__21430),
            .I(N__21395));
    LocalMux I__4942 (
            .O(N__21427),
            .I(N__21392));
    LocalMux I__4941 (
            .O(N__21424),
            .I(N__21389));
    LocalMux I__4940 (
            .O(N__21421),
            .I(N__21386));
    Span4Mux_v I__4939 (
            .O(N__21416),
            .I(N__21379));
    Span4Mux_v I__4938 (
            .O(N__21409),
            .I(N__21379));
    Span4Mux_h I__4937 (
            .O(N__21406),
            .I(N__21379));
    LocalMux I__4936 (
            .O(N__21403),
            .I(N__21374));
    LocalMux I__4935 (
            .O(N__21400),
            .I(N__21374));
    Span4Mux_h I__4934 (
            .O(N__21395),
            .I(N__21371));
    Span12Mux_v I__4933 (
            .O(N__21392),
            .I(N__21368));
    Span4Mux_h I__4932 (
            .O(N__21389),
            .I(N__21365));
    Span4Mux_v I__4931 (
            .O(N__21386),
            .I(N__21360));
    Span4Mux_h I__4930 (
            .O(N__21379),
            .I(N__21360));
    Span4Mux_v I__4929 (
            .O(N__21374),
            .I(N__21357));
    Odrv4 I__4928 (
            .O(N__21371),
            .I(\transmit_module.n4225 ));
    Odrv12 I__4927 (
            .O(N__21368),
            .I(\transmit_module.n4225 ));
    Odrv4 I__4926 (
            .O(N__21365),
            .I(\transmit_module.n4225 ));
    Odrv4 I__4925 (
            .O(N__21360),
            .I(\transmit_module.n4225 ));
    Odrv4 I__4924 (
            .O(N__21357),
            .I(\transmit_module.n4225 ));
    CascadeMux I__4923 (
            .O(N__21346),
            .I(N__21332));
    SRMux I__4922 (
            .O(N__21345),
            .I(N__21329));
    SRMux I__4921 (
            .O(N__21344),
            .I(N__21326));
    SRMux I__4920 (
            .O(N__21343),
            .I(N__21318));
    SRMux I__4919 (
            .O(N__21342),
            .I(N__21314));
    SRMux I__4918 (
            .O(N__21341),
            .I(N__21311));
    SRMux I__4917 (
            .O(N__21340),
            .I(N__21308));
    SRMux I__4916 (
            .O(N__21339),
            .I(N__21303));
    SRMux I__4915 (
            .O(N__21338),
            .I(N__21300));
    SRMux I__4914 (
            .O(N__21337),
            .I(N__21297));
    CascadeMux I__4913 (
            .O(N__21336),
            .I(N__21289));
    CascadeMux I__4912 (
            .O(N__21335),
            .I(N__21285));
    InMux I__4911 (
            .O(N__21332),
            .I(N__21282));
    LocalMux I__4910 (
            .O(N__21329),
            .I(N__21273));
    LocalMux I__4909 (
            .O(N__21326),
            .I(N__21273));
    SRMux I__4908 (
            .O(N__21325),
            .I(N__21270));
    SRMux I__4907 (
            .O(N__21324),
            .I(N__21263));
    SRMux I__4906 (
            .O(N__21323),
            .I(N__21256));
    SRMux I__4905 (
            .O(N__21322),
            .I(N__21253));
    SRMux I__4904 (
            .O(N__21321),
            .I(N__21248));
    LocalMux I__4903 (
            .O(N__21318),
            .I(N__21245));
    SRMux I__4902 (
            .O(N__21317),
            .I(N__21242));
    LocalMux I__4901 (
            .O(N__21314),
            .I(N__21237));
    LocalMux I__4900 (
            .O(N__21311),
            .I(N__21237));
    LocalMux I__4899 (
            .O(N__21308),
            .I(N__21234));
    SRMux I__4898 (
            .O(N__21307),
            .I(N__21231));
    SRMux I__4897 (
            .O(N__21306),
            .I(N__21228));
    LocalMux I__4896 (
            .O(N__21303),
            .I(N__21225));
    LocalMux I__4895 (
            .O(N__21300),
            .I(N__21220));
    LocalMux I__4894 (
            .O(N__21297),
            .I(N__21220));
    SRMux I__4893 (
            .O(N__21296),
            .I(N__21214));
    SRMux I__4892 (
            .O(N__21295),
            .I(N__21211));
    CascadeMux I__4891 (
            .O(N__21294),
            .I(N__21206));
    CascadeMux I__4890 (
            .O(N__21293),
            .I(N__21203));
    CascadeMux I__4889 (
            .O(N__21292),
            .I(N__21200));
    InMux I__4888 (
            .O(N__21289),
            .I(N__21191));
    SRMux I__4887 (
            .O(N__21288),
            .I(N__21188));
    InMux I__4886 (
            .O(N__21285),
            .I(N__21185));
    LocalMux I__4885 (
            .O(N__21282),
            .I(N__21182));
    CascadeMux I__4884 (
            .O(N__21281),
            .I(N__21176));
    CascadeMux I__4883 (
            .O(N__21280),
            .I(N__21173));
    SRMux I__4882 (
            .O(N__21279),
            .I(N__21168));
    SRMux I__4881 (
            .O(N__21278),
            .I(N__21163));
    Span4Mux_v I__4880 (
            .O(N__21273),
            .I(N__21158));
    LocalMux I__4879 (
            .O(N__21270),
            .I(N__21158));
    SRMux I__4878 (
            .O(N__21269),
            .I(N__21155));
    InMux I__4877 (
            .O(N__21268),
            .I(N__21152));
    SRMux I__4876 (
            .O(N__21267),
            .I(N__21148));
    SRMux I__4875 (
            .O(N__21266),
            .I(N__21144));
    LocalMux I__4874 (
            .O(N__21263),
            .I(N__21141));
    SRMux I__4873 (
            .O(N__21262),
            .I(N__21138));
    SRMux I__4872 (
            .O(N__21261),
            .I(N__21135));
    SRMux I__4871 (
            .O(N__21260),
            .I(N__21132));
    CascadeMux I__4870 (
            .O(N__21259),
            .I(N__21129));
    LocalMux I__4869 (
            .O(N__21256),
            .I(N__21124));
    LocalMux I__4868 (
            .O(N__21253),
            .I(N__21124));
    SRMux I__4867 (
            .O(N__21252),
            .I(N__21121));
    SRMux I__4866 (
            .O(N__21251),
            .I(N__21118));
    LocalMux I__4865 (
            .O(N__21248),
            .I(N__21115));
    Span4Mux_h I__4864 (
            .O(N__21245),
            .I(N__21108));
    LocalMux I__4863 (
            .O(N__21242),
            .I(N__21108));
    Span4Mux_h I__4862 (
            .O(N__21237),
            .I(N__21108));
    Span4Mux_v I__4861 (
            .O(N__21234),
            .I(N__21097));
    LocalMux I__4860 (
            .O(N__21231),
            .I(N__21097));
    LocalMux I__4859 (
            .O(N__21228),
            .I(N__21097));
    Span4Mux_h I__4858 (
            .O(N__21225),
            .I(N__21097));
    Span4Mux_h I__4857 (
            .O(N__21220),
            .I(N__21097));
    CascadeMux I__4856 (
            .O(N__21219),
            .I(N__21094));
    InMux I__4855 (
            .O(N__21218),
            .I(N__21087));
    InMux I__4854 (
            .O(N__21217),
            .I(N__21087));
    LocalMux I__4853 (
            .O(N__21214),
            .I(N__21084));
    LocalMux I__4852 (
            .O(N__21211),
            .I(N__21081));
    SRMux I__4851 (
            .O(N__21210),
            .I(N__21078));
    InMux I__4850 (
            .O(N__21209),
            .I(N__21063));
    InMux I__4849 (
            .O(N__21206),
            .I(N__21063));
    InMux I__4848 (
            .O(N__21203),
            .I(N__21063));
    InMux I__4847 (
            .O(N__21200),
            .I(N__21063));
    InMux I__4846 (
            .O(N__21199),
            .I(N__21063));
    InMux I__4845 (
            .O(N__21198),
            .I(N__21063));
    InMux I__4844 (
            .O(N__21197),
            .I(N__21063));
    CascadeMux I__4843 (
            .O(N__21196),
            .I(N__21060));
    CascadeMux I__4842 (
            .O(N__21195),
            .I(N__21057));
    CascadeMux I__4841 (
            .O(N__21194),
            .I(N__21052));
    LocalMux I__4840 (
            .O(N__21191),
            .I(N__21049));
    LocalMux I__4839 (
            .O(N__21188),
            .I(N__21046));
    LocalMux I__4838 (
            .O(N__21185),
            .I(N__21041));
    Span4Mux_h I__4837 (
            .O(N__21182),
            .I(N__21041));
    SRMux I__4836 (
            .O(N__21181),
            .I(N__21038));
    CascadeMux I__4835 (
            .O(N__21180),
            .I(N__21030));
    InMux I__4834 (
            .O(N__21179),
            .I(N__21027));
    InMux I__4833 (
            .O(N__21176),
            .I(N__21024));
    InMux I__4832 (
            .O(N__21173),
            .I(N__21019));
    InMux I__4831 (
            .O(N__21172),
            .I(N__21019));
    IoInMux I__4830 (
            .O(N__21171),
            .I(N__21016));
    LocalMux I__4829 (
            .O(N__21168),
            .I(N__21013));
    SRMux I__4828 (
            .O(N__21167),
            .I(N__21010));
    SRMux I__4827 (
            .O(N__21166),
            .I(N__21007));
    LocalMux I__4826 (
            .O(N__21163),
            .I(N__21000));
    Span4Mux_h I__4825 (
            .O(N__21158),
            .I(N__21000));
    LocalMux I__4824 (
            .O(N__21155),
            .I(N__21000));
    LocalMux I__4823 (
            .O(N__21152),
            .I(N__20997));
    SRMux I__4822 (
            .O(N__21151),
            .I(N__20994));
    LocalMux I__4821 (
            .O(N__21148),
            .I(N__20991));
    SRMux I__4820 (
            .O(N__21147),
            .I(N__20988));
    LocalMux I__4819 (
            .O(N__21144),
            .I(N__20985));
    Span4Mux_h I__4818 (
            .O(N__21141),
            .I(N__20976));
    LocalMux I__4817 (
            .O(N__21138),
            .I(N__20976));
    LocalMux I__4816 (
            .O(N__21135),
            .I(N__20976));
    LocalMux I__4815 (
            .O(N__21132),
            .I(N__20976));
    InMux I__4814 (
            .O(N__21129),
            .I(N__20973));
    Span4Mux_v I__4813 (
            .O(N__21124),
            .I(N__20970));
    LocalMux I__4812 (
            .O(N__21121),
            .I(N__20959));
    LocalMux I__4811 (
            .O(N__21118),
            .I(N__20959));
    Span4Mux_h I__4810 (
            .O(N__21115),
            .I(N__20959));
    Span4Mux_h I__4809 (
            .O(N__21108),
            .I(N__20959));
    Span4Mux_h I__4808 (
            .O(N__21097),
            .I(N__20959));
    InMux I__4807 (
            .O(N__21094),
            .I(N__20956));
    SRMux I__4806 (
            .O(N__21093),
            .I(N__20952));
    SRMux I__4805 (
            .O(N__21092),
            .I(N__20949));
    LocalMux I__4804 (
            .O(N__21087),
            .I(N__20946));
    Span4Mux_h I__4803 (
            .O(N__21084),
            .I(N__20937));
    Span4Mux_h I__4802 (
            .O(N__21081),
            .I(N__20937));
    LocalMux I__4801 (
            .O(N__21078),
            .I(N__20937));
    LocalMux I__4800 (
            .O(N__21063),
            .I(N__20937));
    InMux I__4799 (
            .O(N__21060),
            .I(N__20932));
    InMux I__4798 (
            .O(N__21057),
            .I(N__20932));
    SRMux I__4797 (
            .O(N__21056),
            .I(N__20929));
    SRMux I__4796 (
            .O(N__21055),
            .I(N__20926));
    InMux I__4795 (
            .O(N__21052),
            .I(N__20923));
    Span4Mux_v I__4794 (
            .O(N__21049),
            .I(N__20920));
    Span4Mux_h I__4793 (
            .O(N__21046),
            .I(N__20915));
    Span4Mux_v I__4792 (
            .O(N__21041),
            .I(N__20915));
    LocalMux I__4791 (
            .O(N__21038),
            .I(N__20912));
    InMux I__4790 (
            .O(N__21037),
            .I(N__20909));
    InMux I__4789 (
            .O(N__21036),
            .I(N__20906));
    InMux I__4788 (
            .O(N__21035),
            .I(N__20903));
    InMux I__4787 (
            .O(N__21034),
            .I(N__20896));
    InMux I__4786 (
            .O(N__21033),
            .I(N__20896));
    InMux I__4785 (
            .O(N__21030),
            .I(N__20896));
    LocalMux I__4784 (
            .O(N__21027),
            .I(N__20889));
    LocalMux I__4783 (
            .O(N__21024),
            .I(N__20889));
    LocalMux I__4782 (
            .O(N__21019),
            .I(N__20889));
    LocalMux I__4781 (
            .O(N__21016),
            .I(N__20886));
    Span4Mux_h I__4780 (
            .O(N__21013),
            .I(N__20881));
    LocalMux I__4779 (
            .O(N__21010),
            .I(N__20881));
    LocalMux I__4778 (
            .O(N__21007),
            .I(N__20874));
    Sp12to4 I__4777 (
            .O(N__21000),
            .I(N__20874));
    Sp12to4 I__4776 (
            .O(N__20997),
            .I(N__20874));
    LocalMux I__4775 (
            .O(N__20994),
            .I(N__20871));
    Span4Mux_h I__4774 (
            .O(N__20991),
            .I(N__20862));
    LocalMux I__4773 (
            .O(N__20988),
            .I(N__20862));
    Span4Mux_v I__4772 (
            .O(N__20985),
            .I(N__20862));
    Span4Mux_v I__4771 (
            .O(N__20976),
            .I(N__20862));
    LocalMux I__4770 (
            .O(N__20973),
            .I(N__20853));
    Span4Mux_h I__4769 (
            .O(N__20970),
            .I(N__20853));
    Span4Mux_v I__4768 (
            .O(N__20959),
            .I(N__20853));
    LocalMux I__4767 (
            .O(N__20956),
            .I(N__20853));
    SRMux I__4766 (
            .O(N__20955),
            .I(N__20850));
    LocalMux I__4765 (
            .O(N__20952),
            .I(N__20845));
    LocalMux I__4764 (
            .O(N__20949),
            .I(N__20845));
    Span4Mux_h I__4763 (
            .O(N__20946),
            .I(N__20838));
    Span4Mux_v I__4762 (
            .O(N__20937),
            .I(N__20838));
    LocalMux I__4761 (
            .O(N__20932),
            .I(N__20838));
    LocalMux I__4760 (
            .O(N__20929),
            .I(N__20835));
    LocalMux I__4759 (
            .O(N__20926),
            .I(N__20832));
    LocalMux I__4758 (
            .O(N__20923),
            .I(N__20829));
    Span4Mux_h I__4757 (
            .O(N__20920),
            .I(N__20824));
    Span4Mux_v I__4756 (
            .O(N__20915),
            .I(N__20824));
    Span4Mux_v I__4755 (
            .O(N__20912),
            .I(N__20811));
    LocalMux I__4754 (
            .O(N__20909),
            .I(N__20811));
    LocalMux I__4753 (
            .O(N__20906),
            .I(N__20811));
    LocalMux I__4752 (
            .O(N__20903),
            .I(N__20811));
    LocalMux I__4751 (
            .O(N__20896),
            .I(N__20811));
    Span4Mux_h I__4750 (
            .O(N__20889),
            .I(N__20811));
    Span12Mux_s10_h I__4749 (
            .O(N__20886),
            .I(N__20808));
    Span4Mux_v I__4748 (
            .O(N__20881),
            .I(N__20805));
    Span12Mux_v I__4747 (
            .O(N__20874),
            .I(N__20802));
    Span4Mux_v I__4746 (
            .O(N__20871),
            .I(N__20797));
    Span4Mux_h I__4745 (
            .O(N__20862),
            .I(N__20797));
    Span4Mux_h I__4744 (
            .O(N__20853),
            .I(N__20794));
    LocalMux I__4743 (
            .O(N__20850),
            .I(N__20787));
    Span4Mux_v I__4742 (
            .O(N__20845),
            .I(N__20787));
    Span4Mux_h I__4741 (
            .O(N__20838),
            .I(N__20787));
    Span4Mux_h I__4740 (
            .O(N__20835),
            .I(N__20776));
    Span4Mux_h I__4739 (
            .O(N__20832),
            .I(N__20776));
    Span4Mux_h I__4738 (
            .O(N__20829),
            .I(N__20776));
    Span4Mux_v I__4737 (
            .O(N__20824),
            .I(N__20776));
    Span4Mux_h I__4736 (
            .O(N__20811),
            .I(N__20776));
    Odrv12 I__4735 (
            .O(N__20808),
            .I(ADV_VSYNC_c));
    Odrv4 I__4734 (
            .O(N__20805),
            .I(ADV_VSYNC_c));
    Odrv12 I__4733 (
            .O(N__20802),
            .I(ADV_VSYNC_c));
    Odrv4 I__4732 (
            .O(N__20797),
            .I(ADV_VSYNC_c));
    Odrv4 I__4731 (
            .O(N__20794),
            .I(ADV_VSYNC_c));
    Odrv4 I__4730 (
            .O(N__20787),
            .I(ADV_VSYNC_c));
    Odrv4 I__4729 (
            .O(N__20776),
            .I(ADV_VSYNC_c));
    InMux I__4728 (
            .O(N__20761),
            .I(N__20758));
    LocalMux I__4727 (
            .O(N__20758),
            .I(N__20755));
    Span12Mux_h I__4726 (
            .O(N__20755),
            .I(N__20752));
    Span12Mux_v I__4725 (
            .O(N__20752),
            .I(N__20749));
    Odrv12 I__4724 (
            .O(N__20749),
            .I(\line_buffer.n617 ));
    CascadeMux I__4723 (
            .O(N__20746),
            .I(N__20743));
    InMux I__4722 (
            .O(N__20743),
            .I(N__20740));
    LocalMux I__4721 (
            .O(N__20740),
            .I(N__20737));
    Span4Mux_h I__4720 (
            .O(N__20737),
            .I(N__20734));
    Span4Mux_h I__4719 (
            .O(N__20734),
            .I(N__20731));
    Span4Mux_v I__4718 (
            .O(N__20731),
            .I(N__20728));
    Odrv4 I__4717 (
            .O(N__20728),
            .I(\line_buffer.n609 ));
    InMux I__4716 (
            .O(N__20725),
            .I(N__20722));
    LocalMux I__4715 (
            .O(N__20722),
            .I(N__20719));
    Span4Mux_h I__4714 (
            .O(N__20719),
            .I(N__20716));
    Span4Mux_h I__4713 (
            .O(N__20716),
            .I(N__20713));
    Span4Mux_v I__4712 (
            .O(N__20713),
            .I(N__20710));
    Odrv4 I__4711 (
            .O(N__20710),
            .I(\line_buffer.n610 ));
    CascadeMux I__4710 (
            .O(N__20707),
            .I(N__20704));
    InMux I__4709 (
            .O(N__20704),
            .I(N__20701));
    LocalMux I__4708 (
            .O(N__20701),
            .I(N__20698));
    Span4Mux_v I__4707 (
            .O(N__20698),
            .I(N__20695));
    Sp12to4 I__4706 (
            .O(N__20695),
            .I(N__20692));
    Span12Mux_h I__4705 (
            .O(N__20692),
            .I(N__20689));
    Span12Mux_v I__4704 (
            .O(N__20689),
            .I(N__20686));
    Odrv12 I__4703 (
            .O(N__20686),
            .I(\line_buffer.n618 ));
    InMux I__4702 (
            .O(N__20683),
            .I(N__20680));
    LocalMux I__4701 (
            .O(N__20680),
            .I(\line_buffer.n4161 ));
    InMux I__4700 (
            .O(N__20677),
            .I(N__20674));
    LocalMux I__4699 (
            .O(N__20674),
            .I(N__20671));
    Odrv4 I__4698 (
            .O(N__20671),
            .I(\transmit_module.Y_DELTA_PATTERN_17 ));
    InMux I__4697 (
            .O(N__20668),
            .I(N__20665));
    LocalMux I__4696 (
            .O(N__20665),
            .I(\transmit_module.Y_DELTA_PATTERN_16 ));
    InMux I__4695 (
            .O(N__20662),
            .I(N__20659));
    LocalMux I__4694 (
            .O(N__20659),
            .I(\transmit_module.Y_DELTA_PATTERN_3 ));
    InMux I__4693 (
            .O(N__20656),
            .I(N__20653));
    LocalMux I__4692 (
            .O(N__20653),
            .I(N__20650));
    Odrv4 I__4691 (
            .O(N__20650),
            .I(\transmit_module.Y_DELTA_PATTERN_2 ));
    InMux I__4690 (
            .O(N__20647),
            .I(N__20644));
    LocalMux I__4689 (
            .O(N__20644),
            .I(N__20641));
    Span4Mux_h I__4688 (
            .O(N__20641),
            .I(N__20638));
    Odrv4 I__4687 (
            .O(N__20638),
            .I(\transmit_module.Y_DELTA_PATTERN_22 ));
    InMux I__4686 (
            .O(N__20635),
            .I(N__20632));
    LocalMux I__4685 (
            .O(N__20632),
            .I(\transmit_module.Y_DELTA_PATTERN_24 ));
    InMux I__4684 (
            .O(N__20629),
            .I(N__20626));
    LocalMux I__4683 (
            .O(N__20626),
            .I(\transmit_module.Y_DELTA_PATTERN_23 ));
    CEMux I__4682 (
            .O(N__20623),
            .I(N__20619));
    CEMux I__4681 (
            .O(N__20622),
            .I(N__20615));
    LocalMux I__4680 (
            .O(N__20619),
            .I(N__20611));
    CEMux I__4679 (
            .O(N__20618),
            .I(N__20608));
    LocalMux I__4678 (
            .O(N__20615),
            .I(N__20603));
    CEMux I__4677 (
            .O(N__20614),
            .I(N__20600));
    Span4Mux_v I__4676 (
            .O(N__20611),
            .I(N__20591));
    LocalMux I__4675 (
            .O(N__20608),
            .I(N__20591));
    CEMux I__4674 (
            .O(N__20607),
            .I(N__20588));
    CEMux I__4673 (
            .O(N__20606),
            .I(N__20584));
    Span4Mux_h I__4672 (
            .O(N__20603),
            .I(N__20578));
    LocalMux I__4671 (
            .O(N__20600),
            .I(N__20578));
    CEMux I__4670 (
            .O(N__20599),
            .I(N__20575));
    CEMux I__4669 (
            .O(N__20598),
            .I(N__20572));
    CEMux I__4668 (
            .O(N__20597),
            .I(N__20569));
    CEMux I__4667 (
            .O(N__20596),
            .I(N__20566));
    Span4Mux_h I__4666 (
            .O(N__20591),
            .I(N__20560));
    LocalMux I__4665 (
            .O(N__20588),
            .I(N__20560));
    SRMux I__4664 (
            .O(N__20587),
            .I(N__20557));
    LocalMux I__4663 (
            .O(N__20584),
            .I(N__20554));
    SRMux I__4662 (
            .O(N__20583),
            .I(N__20551));
    Span4Mux_v I__4661 (
            .O(N__20578),
            .I(N__20547));
    LocalMux I__4660 (
            .O(N__20575),
            .I(N__20542));
    LocalMux I__4659 (
            .O(N__20572),
            .I(N__20542));
    LocalMux I__4658 (
            .O(N__20569),
            .I(N__20539));
    LocalMux I__4657 (
            .O(N__20566),
            .I(N__20536));
    SRMux I__4656 (
            .O(N__20565),
            .I(N__20533));
    Span4Mux_v I__4655 (
            .O(N__20560),
            .I(N__20530));
    LocalMux I__4654 (
            .O(N__20557),
            .I(N__20527));
    Span4Mux_v I__4653 (
            .O(N__20554),
            .I(N__20522));
    LocalMux I__4652 (
            .O(N__20551),
            .I(N__20522));
    SRMux I__4651 (
            .O(N__20550),
            .I(N__20519));
    Span4Mux_h I__4650 (
            .O(N__20547),
            .I(N__20514));
    Span4Mux_v I__4649 (
            .O(N__20542),
            .I(N__20514));
    Span4Mux_v I__4648 (
            .O(N__20539),
            .I(N__20511));
    Sp12to4 I__4647 (
            .O(N__20536),
            .I(N__20508));
    LocalMux I__4646 (
            .O(N__20533),
            .I(N__20505));
    Span4Mux_h I__4645 (
            .O(N__20530),
            .I(N__20496));
    Span4Mux_v I__4644 (
            .O(N__20527),
            .I(N__20496));
    Span4Mux_h I__4643 (
            .O(N__20522),
            .I(N__20496));
    LocalMux I__4642 (
            .O(N__20519),
            .I(N__20496));
    Odrv4 I__4641 (
            .O(N__20514),
            .I(\transmit_module.n4224 ));
    Odrv4 I__4640 (
            .O(N__20511),
            .I(\transmit_module.n4224 ));
    Odrv12 I__4639 (
            .O(N__20508),
            .I(\transmit_module.n4224 ));
    Odrv12 I__4638 (
            .O(N__20505),
            .I(\transmit_module.n4224 ));
    Odrv4 I__4637 (
            .O(N__20496),
            .I(\transmit_module.n4224 ));
    InMux I__4636 (
            .O(N__20485),
            .I(N__20482));
    LocalMux I__4635 (
            .O(N__20482),
            .I(N__20479));
    Span4Mux_v I__4634 (
            .O(N__20479),
            .I(N__20476));
    Span4Mux_h I__4633 (
            .O(N__20476),
            .I(N__20473));
    Odrv4 I__4632 (
            .O(N__20473),
            .I(\line_buffer.n642 ));
    CascadeMux I__4631 (
            .O(N__20470),
            .I(N__20467));
    InMux I__4630 (
            .O(N__20467),
            .I(N__20464));
    LocalMux I__4629 (
            .O(N__20464),
            .I(N__20461));
    Span4Mux_v I__4628 (
            .O(N__20461),
            .I(N__20458));
    Span4Mux_v I__4627 (
            .O(N__20458),
            .I(N__20455));
    Sp12to4 I__4626 (
            .O(N__20455),
            .I(N__20452));
    Odrv12 I__4625 (
            .O(N__20452),
            .I(\line_buffer.n650 ));
    InMux I__4624 (
            .O(N__20449),
            .I(N__20446));
    LocalMux I__4623 (
            .O(N__20446),
            .I(N__20443));
    Span4Mux_v I__4622 (
            .O(N__20443),
            .I(N__20440));
    Sp12to4 I__4621 (
            .O(N__20440),
            .I(N__20437));
    Span12Mux_h I__4620 (
            .O(N__20437),
            .I(N__20434));
    Span12Mux_v I__4619 (
            .O(N__20434),
            .I(N__20431));
    Odrv12 I__4618 (
            .O(N__20431),
            .I(\line_buffer.n545 ));
    CascadeMux I__4617 (
            .O(N__20428),
            .I(\line_buffer.n4164_cascade_ ));
    InMux I__4616 (
            .O(N__20425),
            .I(N__20422));
    LocalMux I__4615 (
            .O(N__20422),
            .I(N__20419));
    Span4Mux_h I__4614 (
            .O(N__20419),
            .I(N__20416));
    Span4Mux_v I__4613 (
            .O(N__20416),
            .I(N__20413));
    Span4Mux_h I__4612 (
            .O(N__20413),
            .I(N__20410));
    Odrv4 I__4611 (
            .O(N__20410),
            .I(\line_buffer.n553 ));
    CascadeMux I__4610 (
            .O(N__20407),
            .I(\line_buffer.n4167_cascade_ ));
    InMux I__4609 (
            .O(N__20404),
            .I(N__20401));
    LocalMux I__4608 (
            .O(N__20401),
            .I(N__20398));
    Span4Mux_h I__4607 (
            .O(N__20398),
            .I(N__20395));
    Span4Mux_h I__4606 (
            .O(N__20395),
            .I(N__20392));
    Odrv4 I__4605 (
            .O(N__20392),
            .I(TX_DATA_1));
    InMux I__4604 (
            .O(N__20389),
            .I(N__20386));
    LocalMux I__4603 (
            .O(N__20386),
            .I(N__20383));
    Span12Mux_v I__4602 (
            .O(N__20383),
            .I(N__20380));
    Odrv12 I__4601 (
            .O(N__20380),
            .I(\line_buffer.n4065 ));
    InMux I__4600 (
            .O(N__20377),
            .I(N__20374));
    LocalMux I__4599 (
            .O(N__20374),
            .I(N__20371));
    Span4Mux_v I__4598 (
            .O(N__20371),
            .I(N__20368));
    Span4Mux_v I__4597 (
            .O(N__20368),
            .I(N__20365));
    Sp12to4 I__4596 (
            .O(N__20365),
            .I(N__20362));
    Odrv12 I__4595 (
            .O(N__20362),
            .I(\line_buffer.n620 ));
    InMux I__4594 (
            .O(N__20359),
            .I(N__20356));
    LocalMux I__4593 (
            .O(N__20356),
            .I(N__20353));
    Odrv12 I__4592 (
            .O(N__20353),
            .I(\line_buffer.n612 ));
    InMux I__4591 (
            .O(N__20350),
            .I(N__20347));
    LocalMux I__4590 (
            .O(N__20347),
            .I(\transmit_module.Y_DELTA_PATTERN_6 ));
    InMux I__4589 (
            .O(N__20344),
            .I(N__20341));
    LocalMux I__4588 (
            .O(N__20341),
            .I(\transmit_module.Y_DELTA_PATTERN_5 ));
    InMux I__4587 (
            .O(N__20338),
            .I(N__20335));
    LocalMux I__4586 (
            .O(N__20335),
            .I(\transmit_module.Y_DELTA_PATTERN_7 ));
    InMux I__4585 (
            .O(N__20332),
            .I(N__20329));
    LocalMux I__4584 (
            .O(N__20329),
            .I(\transmit_module.Y_DELTA_PATTERN_11 ));
    InMux I__4583 (
            .O(N__20326),
            .I(N__20323));
    LocalMux I__4582 (
            .O(N__20323),
            .I(\transmit_module.Y_DELTA_PATTERN_10 ));
    InMux I__4581 (
            .O(N__20320),
            .I(N__20317));
    LocalMux I__4580 (
            .O(N__20317),
            .I(\transmit_module.Y_DELTA_PATTERN_9 ));
    InMux I__4579 (
            .O(N__20314),
            .I(N__20311));
    LocalMux I__4578 (
            .O(N__20311),
            .I(\transmit_module.Y_DELTA_PATTERN_8 ));
    InMux I__4577 (
            .O(N__20308),
            .I(N__20305));
    LocalMux I__4576 (
            .O(N__20305),
            .I(\transmit_module.Y_DELTA_PATTERN_15 ));
    InMux I__4575 (
            .O(N__20302),
            .I(N__20299));
    LocalMux I__4574 (
            .O(N__20299),
            .I(N__20296));
    Odrv4 I__4573 (
            .O(N__20296),
            .I(\transmit_module.Y_DELTA_PATTERN_4 ));
    InMux I__4572 (
            .O(N__20293),
            .I(N__20290));
    LocalMux I__4571 (
            .O(N__20290),
            .I(\transmit_module.Y_DELTA_PATTERN_37 ));
    InMux I__4570 (
            .O(N__20287),
            .I(N__20284));
    LocalMux I__4569 (
            .O(N__20284),
            .I(\transmit_module.Y_DELTA_PATTERN_36 ));
    InMux I__4568 (
            .O(N__20281),
            .I(N__20278));
    LocalMux I__4567 (
            .O(N__20278),
            .I(\transmit_module.Y_DELTA_PATTERN_38 ));
    InMux I__4566 (
            .O(N__20275),
            .I(N__20271));
    InMux I__4565 (
            .O(N__20274),
            .I(N__20268));
    LocalMux I__4564 (
            .O(N__20271),
            .I(N__20265));
    LocalMux I__4563 (
            .O(N__20268),
            .I(\transmit_module.n185 ));
    Odrv4 I__4562 (
            .O(N__20265),
            .I(\transmit_module.n185 ));
    InMux I__4561 (
            .O(N__20260),
            .I(N__20256));
    InMux I__4560 (
            .O(N__20259),
            .I(N__20253));
    LocalMux I__4559 (
            .O(N__20256),
            .I(N__20250));
    LocalMux I__4558 (
            .O(N__20253),
            .I(\transmit_module.n216 ));
    Odrv12 I__4557 (
            .O(N__20250),
            .I(\transmit_module.n216 ));
    InMux I__4556 (
            .O(N__20245),
            .I(N__20242));
    LocalMux I__4555 (
            .O(N__20242),
            .I(N__20236));
    InMux I__4554 (
            .O(N__20241),
            .I(N__20233));
    InMux I__4553 (
            .O(N__20240),
            .I(N__20230));
    InMux I__4552 (
            .O(N__20239),
            .I(N__20225));
    Span4Mux_h I__4551 (
            .O(N__20236),
            .I(N__20220));
    LocalMux I__4550 (
            .O(N__20233),
            .I(N__20220));
    LocalMux I__4549 (
            .O(N__20230),
            .I(N__20217));
    InMux I__4548 (
            .O(N__20229),
            .I(N__20210));
    InMux I__4547 (
            .O(N__20228),
            .I(N__20210));
    LocalMux I__4546 (
            .O(N__20225),
            .I(N__20202));
    Span4Mux_v I__4545 (
            .O(N__20220),
            .I(N__20202));
    Span4Mux_h I__4544 (
            .O(N__20217),
            .I(N__20202));
    InMux I__4543 (
            .O(N__20216),
            .I(N__20199));
    InMux I__4542 (
            .O(N__20215),
            .I(N__20188));
    LocalMux I__4541 (
            .O(N__20210),
            .I(N__20185));
    InMux I__4540 (
            .O(N__20209),
            .I(N__20182));
    Span4Mux_v I__4539 (
            .O(N__20202),
            .I(N__20179));
    LocalMux I__4538 (
            .O(N__20199),
            .I(N__20176));
    InMux I__4537 (
            .O(N__20198),
            .I(N__20171));
    InMux I__4536 (
            .O(N__20197),
            .I(N__20171));
    InMux I__4535 (
            .O(N__20196),
            .I(N__20153));
    InMux I__4534 (
            .O(N__20195),
            .I(N__20153));
    InMux I__4533 (
            .O(N__20194),
            .I(N__20153));
    InMux I__4532 (
            .O(N__20193),
            .I(N__20153));
    InMux I__4531 (
            .O(N__20192),
            .I(N__20153));
    InMux I__4530 (
            .O(N__20191),
            .I(N__20153));
    LocalMux I__4529 (
            .O(N__20188),
            .I(N__20150));
    Span4Mux_v I__4528 (
            .O(N__20185),
            .I(N__20139));
    LocalMux I__4527 (
            .O(N__20182),
            .I(N__20139));
    Span4Mux_v I__4526 (
            .O(N__20179),
            .I(N__20139));
    Span4Mux_h I__4525 (
            .O(N__20176),
            .I(N__20139));
    LocalMux I__4524 (
            .O(N__20171),
            .I(N__20139));
    InMux I__4523 (
            .O(N__20170),
            .I(N__20132));
    InMux I__4522 (
            .O(N__20169),
            .I(N__20132));
    InMux I__4521 (
            .O(N__20168),
            .I(N__20132));
    InMux I__4520 (
            .O(N__20167),
            .I(N__20127));
    InMux I__4519 (
            .O(N__20166),
            .I(N__20127));
    LocalMux I__4518 (
            .O(N__20153),
            .I(\transmit_module.n4211 ));
    Odrv4 I__4517 (
            .O(N__20150),
            .I(\transmit_module.n4211 ));
    Odrv4 I__4516 (
            .O(N__20139),
            .I(\transmit_module.n4211 ));
    LocalMux I__4515 (
            .O(N__20132),
            .I(\transmit_module.n4211 ));
    LocalMux I__4514 (
            .O(N__20127),
            .I(\transmit_module.n4211 ));
    CascadeMux I__4513 (
            .O(N__20116),
            .I(N__20112));
    CascadeMux I__4512 (
            .O(N__20115),
            .I(N__20109));
    CascadeBuf I__4511 (
            .O(N__20112),
            .I(N__20106));
    CascadeBuf I__4510 (
            .O(N__20109),
            .I(N__20103));
    CascadeMux I__4509 (
            .O(N__20106),
            .I(N__20100));
    CascadeMux I__4508 (
            .O(N__20103),
            .I(N__20097));
    CascadeBuf I__4507 (
            .O(N__20100),
            .I(N__20094));
    CascadeBuf I__4506 (
            .O(N__20097),
            .I(N__20091));
    CascadeMux I__4505 (
            .O(N__20094),
            .I(N__20088));
    CascadeMux I__4504 (
            .O(N__20091),
            .I(N__20085));
    CascadeBuf I__4503 (
            .O(N__20088),
            .I(N__20082));
    CascadeBuf I__4502 (
            .O(N__20085),
            .I(N__20079));
    CascadeMux I__4501 (
            .O(N__20082),
            .I(N__20076));
    CascadeMux I__4500 (
            .O(N__20079),
            .I(N__20073));
    CascadeBuf I__4499 (
            .O(N__20076),
            .I(N__20070));
    CascadeBuf I__4498 (
            .O(N__20073),
            .I(N__20067));
    CascadeMux I__4497 (
            .O(N__20070),
            .I(N__20064));
    CascadeMux I__4496 (
            .O(N__20067),
            .I(N__20061));
    CascadeBuf I__4495 (
            .O(N__20064),
            .I(N__20058));
    CascadeBuf I__4494 (
            .O(N__20061),
            .I(N__20055));
    CascadeMux I__4493 (
            .O(N__20058),
            .I(N__20052));
    CascadeMux I__4492 (
            .O(N__20055),
            .I(N__20049));
    CascadeBuf I__4491 (
            .O(N__20052),
            .I(N__20046));
    CascadeBuf I__4490 (
            .O(N__20049),
            .I(N__20043));
    CascadeMux I__4489 (
            .O(N__20046),
            .I(N__20040));
    CascadeMux I__4488 (
            .O(N__20043),
            .I(N__20037));
    CascadeBuf I__4487 (
            .O(N__20040),
            .I(N__20034));
    CascadeBuf I__4486 (
            .O(N__20037),
            .I(N__20031));
    CascadeMux I__4485 (
            .O(N__20034),
            .I(N__20028));
    CascadeMux I__4484 (
            .O(N__20031),
            .I(N__20025));
    CascadeBuf I__4483 (
            .O(N__20028),
            .I(N__20022));
    CascadeBuf I__4482 (
            .O(N__20025),
            .I(N__20019));
    CascadeMux I__4481 (
            .O(N__20022),
            .I(N__20016));
    CascadeMux I__4480 (
            .O(N__20019),
            .I(N__20013));
    CascadeBuf I__4479 (
            .O(N__20016),
            .I(N__20010));
    CascadeBuf I__4478 (
            .O(N__20013),
            .I(N__20007));
    CascadeMux I__4477 (
            .O(N__20010),
            .I(N__20004));
    CascadeMux I__4476 (
            .O(N__20007),
            .I(N__20001));
    CascadeBuf I__4475 (
            .O(N__20004),
            .I(N__19998));
    CascadeBuf I__4474 (
            .O(N__20001),
            .I(N__19995));
    CascadeMux I__4473 (
            .O(N__19998),
            .I(N__19992));
    CascadeMux I__4472 (
            .O(N__19995),
            .I(N__19989));
    CascadeBuf I__4471 (
            .O(N__19992),
            .I(N__19986));
    CascadeBuf I__4470 (
            .O(N__19989),
            .I(N__19983));
    CascadeMux I__4469 (
            .O(N__19986),
            .I(N__19980));
    CascadeMux I__4468 (
            .O(N__19983),
            .I(N__19977));
    CascadeBuf I__4467 (
            .O(N__19980),
            .I(N__19974));
    CascadeBuf I__4466 (
            .O(N__19977),
            .I(N__19971));
    CascadeMux I__4465 (
            .O(N__19974),
            .I(N__19968));
    CascadeMux I__4464 (
            .O(N__19971),
            .I(N__19965));
    CascadeBuf I__4463 (
            .O(N__19968),
            .I(N__19962));
    CascadeBuf I__4462 (
            .O(N__19965),
            .I(N__19959));
    CascadeMux I__4461 (
            .O(N__19962),
            .I(N__19956));
    CascadeMux I__4460 (
            .O(N__19959),
            .I(N__19953));
    CascadeBuf I__4459 (
            .O(N__19956),
            .I(N__19950));
    CascadeBuf I__4458 (
            .O(N__19953),
            .I(N__19947));
    CascadeMux I__4457 (
            .O(N__19950),
            .I(N__19944));
    CascadeMux I__4456 (
            .O(N__19947),
            .I(N__19941));
    CascadeBuf I__4455 (
            .O(N__19944),
            .I(N__19938));
    CascadeBuf I__4454 (
            .O(N__19941),
            .I(N__19935));
    CascadeMux I__4453 (
            .O(N__19938),
            .I(N__19932));
    CascadeMux I__4452 (
            .O(N__19935),
            .I(N__19929));
    InMux I__4451 (
            .O(N__19932),
            .I(N__19926));
    InMux I__4450 (
            .O(N__19929),
            .I(N__19923));
    LocalMux I__4449 (
            .O(N__19926),
            .I(N__19920));
    LocalMux I__4448 (
            .O(N__19923),
            .I(N__19917));
    Span12Mux_h I__4447 (
            .O(N__19920),
            .I(N__19912));
    Span12Mux_h I__4446 (
            .O(N__19917),
            .I(N__19912));
    Span12Mux_v I__4445 (
            .O(N__19912),
            .I(N__19909));
    Odrv12 I__4444 (
            .O(N__19909),
            .I(n25));
    CascadeMux I__4443 (
            .O(N__19906),
            .I(N__19903));
    InMux I__4442 (
            .O(N__19903),
            .I(N__19900));
    LocalMux I__4441 (
            .O(N__19900),
            .I(\transmit_module.ADDR_Y_COMPONENT_12 ));
    CascadeMux I__4440 (
            .O(N__19897),
            .I(N__19894));
    InMux I__4439 (
            .O(N__19894),
            .I(N__19891));
    LocalMux I__4438 (
            .O(N__19891),
            .I(N__19888));
    Span4Mux_v I__4437 (
            .O(N__19888),
            .I(N__19885));
    Odrv4 I__4436 (
            .O(N__19885),
            .I(\transmit_module.ADDR_Y_COMPONENT_13 ));
    CEMux I__4435 (
            .O(N__19882),
            .I(N__19878));
    CEMux I__4434 (
            .O(N__19881),
            .I(N__19871));
    LocalMux I__4433 (
            .O(N__19878),
            .I(N__19866));
    CEMux I__4432 (
            .O(N__19877),
            .I(N__19863));
    CEMux I__4431 (
            .O(N__19876),
            .I(N__19860));
    CEMux I__4430 (
            .O(N__19875),
            .I(N__19857));
    CEMux I__4429 (
            .O(N__19874),
            .I(N__19854));
    LocalMux I__4428 (
            .O(N__19871),
            .I(N__19850));
    CEMux I__4427 (
            .O(N__19870),
            .I(N__19847));
    CEMux I__4426 (
            .O(N__19869),
            .I(N__19844));
    Span4Mux_v I__4425 (
            .O(N__19866),
            .I(N__19841));
    LocalMux I__4424 (
            .O(N__19863),
            .I(N__19836));
    LocalMux I__4423 (
            .O(N__19860),
            .I(N__19836));
    LocalMux I__4422 (
            .O(N__19857),
            .I(N__19831));
    LocalMux I__4421 (
            .O(N__19854),
            .I(N__19831));
    CEMux I__4420 (
            .O(N__19853),
            .I(N__19828));
    Span4Mux_h I__4419 (
            .O(N__19850),
            .I(N__19825));
    LocalMux I__4418 (
            .O(N__19847),
            .I(N__19822));
    LocalMux I__4417 (
            .O(N__19844),
            .I(N__19819));
    Span4Mux_v I__4416 (
            .O(N__19841),
            .I(N__19814));
    Span4Mux_h I__4415 (
            .O(N__19836),
            .I(N__19814));
    Span4Mux_v I__4414 (
            .O(N__19831),
            .I(N__19809));
    LocalMux I__4413 (
            .O(N__19828),
            .I(N__19809));
    Span4Mux_v I__4412 (
            .O(N__19825),
            .I(N__19804));
    Span4Mux_h I__4411 (
            .O(N__19822),
            .I(N__19804));
    Span4Mux_h I__4410 (
            .O(N__19819),
            .I(N__19799));
    Span4Mux_h I__4409 (
            .O(N__19814),
            .I(N__19799));
    Span4Mux_h I__4408 (
            .O(N__19809),
            .I(N__19796));
    Odrv4 I__4407 (
            .O(N__19804),
            .I(\transmit_module.n2305 ));
    Odrv4 I__4406 (
            .O(N__19799),
            .I(\transmit_module.n2305 ));
    Odrv4 I__4405 (
            .O(N__19796),
            .I(\transmit_module.n2305 ));
    InMux I__4404 (
            .O(N__19789),
            .I(N__19786));
    LocalMux I__4403 (
            .O(N__19786),
            .I(N__19783));
    Odrv4 I__4402 (
            .O(N__19783),
            .I(\transmit_module.Y_DELTA_PATTERN_39 ));
    InMux I__4401 (
            .O(N__19780),
            .I(N__19777));
    LocalMux I__4400 (
            .O(N__19777),
            .I(\transmit_module.Y_DELTA_PATTERN_41 ));
    InMux I__4399 (
            .O(N__19774),
            .I(N__19771));
    LocalMux I__4398 (
            .O(N__19771),
            .I(\transmit_module.Y_DELTA_PATTERN_40 ));
    InMux I__4397 (
            .O(N__19768),
            .I(N__19765));
    LocalMux I__4396 (
            .O(N__19765),
            .I(\transmit_module.Y_DELTA_PATTERN_12 ));
    InMux I__4395 (
            .O(N__19762),
            .I(N__19759));
    LocalMux I__4394 (
            .O(N__19759),
            .I(\transmit_module.Y_DELTA_PATTERN_32 ));
    InMux I__4393 (
            .O(N__19756),
            .I(N__19753));
    LocalMux I__4392 (
            .O(N__19753),
            .I(\transmit_module.Y_DELTA_PATTERN_13 ));
    InMux I__4391 (
            .O(N__19750),
            .I(N__19747));
    LocalMux I__4390 (
            .O(N__19747),
            .I(\transmit_module.Y_DELTA_PATTERN_14 ));
    InMux I__4389 (
            .O(N__19744),
            .I(N__19741));
    LocalMux I__4388 (
            .O(N__19741),
            .I(\transmit_module.Y_DELTA_PATTERN_26 ));
    InMux I__4387 (
            .O(N__19738),
            .I(N__19735));
    LocalMux I__4386 (
            .O(N__19735),
            .I(\transmit_module.Y_DELTA_PATTERN_25 ));
    InMux I__4385 (
            .O(N__19732),
            .I(N__19729));
    LocalMux I__4384 (
            .O(N__19729),
            .I(N__19726));
    Odrv4 I__4383 (
            .O(N__19726),
            .I(\transmit_module.Y_DELTA_PATTERN_28 ));
    InMux I__4382 (
            .O(N__19723),
            .I(N__19720));
    LocalMux I__4381 (
            .O(N__19720),
            .I(\transmit_module.Y_DELTA_PATTERN_27 ));
    InMux I__4380 (
            .O(N__19717),
            .I(N__19710));
    InMux I__4379 (
            .O(N__19716),
            .I(N__19707));
    InMux I__4378 (
            .O(N__19715),
            .I(N__19702));
    InMux I__4377 (
            .O(N__19714),
            .I(N__19702));
    InMux I__4376 (
            .O(N__19713),
            .I(N__19698));
    LocalMux I__4375 (
            .O(N__19710),
            .I(N__19694));
    LocalMux I__4374 (
            .O(N__19707),
            .I(N__19686));
    LocalMux I__4373 (
            .O(N__19702),
            .I(N__19686));
    InMux I__4372 (
            .O(N__19701),
            .I(N__19683));
    LocalMux I__4371 (
            .O(N__19698),
            .I(N__19680));
    InMux I__4370 (
            .O(N__19697),
            .I(N__19677));
    Span4Mux_v I__4369 (
            .O(N__19694),
            .I(N__19674));
    InMux I__4368 (
            .O(N__19693),
            .I(N__19671));
    InMux I__4367 (
            .O(N__19692),
            .I(N__19667));
    InMux I__4366 (
            .O(N__19691),
            .I(N__19664));
    Span4Mux_v I__4365 (
            .O(N__19686),
            .I(N__19658));
    LocalMux I__4364 (
            .O(N__19683),
            .I(N__19651));
    Span4Mux_v I__4363 (
            .O(N__19680),
            .I(N__19651));
    LocalMux I__4362 (
            .O(N__19677),
            .I(N__19651));
    Span4Mux_h I__4361 (
            .O(N__19674),
            .I(N__19646));
    LocalMux I__4360 (
            .O(N__19671),
            .I(N__19646));
    InMux I__4359 (
            .O(N__19670),
            .I(N__19643));
    LocalMux I__4358 (
            .O(N__19667),
            .I(N__19638));
    LocalMux I__4357 (
            .O(N__19664),
            .I(N__19638));
    InMux I__4356 (
            .O(N__19663),
            .I(N__19635));
    InMux I__4355 (
            .O(N__19662),
            .I(N__19632));
    InMux I__4354 (
            .O(N__19661),
            .I(N__19629));
    Span4Mux_h I__4353 (
            .O(N__19658),
            .I(N__19626));
    Span4Mux_v I__4352 (
            .O(N__19651),
            .I(N__19623));
    Span4Mux_v I__4351 (
            .O(N__19646),
            .I(N__19612));
    LocalMux I__4350 (
            .O(N__19643),
            .I(N__19612));
    Span4Mux_h I__4349 (
            .O(N__19638),
            .I(N__19612));
    LocalMux I__4348 (
            .O(N__19635),
            .I(N__19612));
    LocalMux I__4347 (
            .O(N__19632),
            .I(N__19612));
    LocalMux I__4346 (
            .O(N__19629),
            .I(\transmit_module.Y_DELTA_PATTERN_0 ));
    Odrv4 I__4345 (
            .O(N__19626),
            .I(\transmit_module.Y_DELTA_PATTERN_0 ));
    Odrv4 I__4344 (
            .O(N__19623),
            .I(\transmit_module.Y_DELTA_PATTERN_0 ));
    Odrv4 I__4343 (
            .O(N__19612),
            .I(\transmit_module.Y_DELTA_PATTERN_0 ));
    InMux I__4342 (
            .O(N__19603),
            .I(N__19600));
    LocalMux I__4341 (
            .O(N__19600),
            .I(N__19597));
    Span4Mux_h I__4340 (
            .O(N__19597),
            .I(N__19594));
    Span4Mux_h I__4339 (
            .O(N__19594),
            .I(N__19591));
    Odrv4 I__4338 (
            .O(N__19591),
            .I(\transmit_module.Y_DELTA_PATTERN_99 ));
    InMux I__4337 (
            .O(N__19588),
            .I(N__19584));
    InMux I__4336 (
            .O(N__19587),
            .I(N__19579));
    LocalMux I__4335 (
            .O(N__19584),
            .I(N__19576));
    InMux I__4334 (
            .O(N__19583),
            .I(N__19573));
    InMux I__4333 (
            .O(N__19582),
            .I(N__19569));
    LocalMux I__4332 (
            .O(N__19579),
            .I(N__19566));
    Span4Mux_h I__4331 (
            .O(N__19576),
            .I(N__19563));
    LocalMux I__4330 (
            .O(N__19573),
            .I(N__19560));
    InMux I__4329 (
            .O(N__19572),
            .I(N__19557));
    LocalMux I__4328 (
            .O(N__19569),
            .I(N__19552));
    Span4Mux_h I__4327 (
            .O(N__19566),
            .I(N__19552));
    Odrv4 I__4326 (
            .O(N__19563),
            .I(\transmit_module.n4220 ));
    Odrv12 I__4325 (
            .O(N__19560),
            .I(\transmit_module.n4220 ));
    LocalMux I__4324 (
            .O(N__19557),
            .I(\transmit_module.n4220 ));
    Odrv4 I__4323 (
            .O(N__19552),
            .I(\transmit_module.n4220 ));
    InMux I__4322 (
            .O(N__19543),
            .I(N__19540));
    LocalMux I__4321 (
            .O(N__19540),
            .I(N__19537));
    Odrv4 I__4320 (
            .O(N__19537),
            .I(\transmit_module.n192 ));
    InMux I__4319 (
            .O(N__19534),
            .I(N__19529));
    CascadeMux I__4318 (
            .O(N__19533),
            .I(N__19526));
    InMux I__4317 (
            .O(N__19532),
            .I(N__19522));
    LocalMux I__4316 (
            .O(N__19529),
            .I(N__19517));
    InMux I__4315 (
            .O(N__19526),
            .I(N__19514));
    InMux I__4314 (
            .O(N__19525),
            .I(N__19508));
    LocalMux I__4313 (
            .O(N__19522),
            .I(N__19505));
    InMux I__4312 (
            .O(N__19521),
            .I(N__19502));
    InMux I__4311 (
            .O(N__19520),
            .I(N__19497));
    Span4Mux_v I__4310 (
            .O(N__19517),
            .I(N__19487));
    LocalMux I__4309 (
            .O(N__19514),
            .I(N__19487));
    InMux I__4308 (
            .O(N__19513),
            .I(N__19480));
    InMux I__4307 (
            .O(N__19512),
            .I(N__19480));
    InMux I__4306 (
            .O(N__19511),
            .I(N__19480));
    LocalMux I__4305 (
            .O(N__19508),
            .I(N__19477));
    Span4Mux_v I__4304 (
            .O(N__19505),
            .I(N__19472));
    LocalMux I__4303 (
            .O(N__19502),
            .I(N__19472));
    InMux I__4302 (
            .O(N__19501),
            .I(N__19462));
    InMux I__4301 (
            .O(N__19500),
            .I(N__19462));
    LocalMux I__4300 (
            .O(N__19497),
            .I(N__19459));
    InMux I__4299 (
            .O(N__19496),
            .I(N__19448));
    InMux I__4298 (
            .O(N__19495),
            .I(N__19448));
    InMux I__4297 (
            .O(N__19494),
            .I(N__19448));
    InMux I__4296 (
            .O(N__19493),
            .I(N__19448));
    InMux I__4295 (
            .O(N__19492),
            .I(N__19448));
    Sp12to4 I__4294 (
            .O(N__19487),
            .I(N__19443));
    LocalMux I__4293 (
            .O(N__19480),
            .I(N__19443));
    Span4Mux_h I__4292 (
            .O(N__19477),
            .I(N__19438));
    Span4Mux_h I__4291 (
            .O(N__19472),
            .I(N__19438));
    InMux I__4290 (
            .O(N__19471),
            .I(N__19433));
    InMux I__4289 (
            .O(N__19470),
            .I(N__19433));
    InMux I__4288 (
            .O(N__19469),
            .I(N__19426));
    InMux I__4287 (
            .O(N__19468),
            .I(N__19426));
    InMux I__4286 (
            .O(N__19467),
            .I(N__19426));
    LocalMux I__4285 (
            .O(N__19462),
            .I(\transmit_module.n3926 ));
    Odrv12 I__4284 (
            .O(N__19459),
            .I(\transmit_module.n3926 ));
    LocalMux I__4283 (
            .O(N__19448),
            .I(\transmit_module.n3926 ));
    Odrv12 I__4282 (
            .O(N__19443),
            .I(\transmit_module.n3926 ));
    Odrv4 I__4281 (
            .O(N__19438),
            .I(\transmit_module.n3926 ));
    LocalMux I__4280 (
            .O(N__19433),
            .I(\transmit_module.n3926 ));
    LocalMux I__4279 (
            .O(N__19426),
            .I(\transmit_module.n3926 ));
    CEMux I__4278 (
            .O(N__19411),
            .I(N__19407));
    CEMux I__4277 (
            .O(N__19410),
            .I(N__19404));
    LocalMux I__4276 (
            .O(N__19407),
            .I(N__19401));
    LocalMux I__4275 (
            .O(N__19404),
            .I(N__19398));
    Span4Mux_h I__4274 (
            .O(N__19401),
            .I(N__19394));
    Span4Mux_h I__4273 (
            .O(N__19398),
            .I(N__19391));
    InMux I__4272 (
            .O(N__19397),
            .I(N__19388));
    Odrv4 I__4271 (
            .O(N__19394),
            .I(\transmit_module.n2277 ));
    Odrv4 I__4270 (
            .O(N__19391),
            .I(\transmit_module.n2277 ));
    LocalMux I__4269 (
            .O(N__19388),
            .I(\transmit_module.n2277 ));
    InMux I__4268 (
            .O(N__19381),
            .I(N__19378));
    LocalMux I__4267 (
            .O(N__19378),
            .I(N__19375));
    Odrv4 I__4266 (
            .O(N__19375),
            .I(\transmit_module.Y_DELTA_PATTERN_42 ));
    InMux I__4265 (
            .O(N__19372),
            .I(N__19369));
    LocalMux I__4264 (
            .O(N__19369),
            .I(N__19356));
    ClkMux I__4263 (
            .O(N__19368),
            .I(N__19228));
    ClkMux I__4262 (
            .O(N__19367),
            .I(N__19228));
    ClkMux I__4261 (
            .O(N__19366),
            .I(N__19228));
    ClkMux I__4260 (
            .O(N__19365),
            .I(N__19228));
    ClkMux I__4259 (
            .O(N__19364),
            .I(N__19228));
    ClkMux I__4258 (
            .O(N__19363),
            .I(N__19228));
    ClkMux I__4257 (
            .O(N__19362),
            .I(N__19228));
    ClkMux I__4256 (
            .O(N__19361),
            .I(N__19228));
    ClkMux I__4255 (
            .O(N__19360),
            .I(N__19228));
    ClkMux I__4254 (
            .O(N__19359),
            .I(N__19228));
    Glb2LocalMux I__4253 (
            .O(N__19356),
            .I(N__19228));
    ClkMux I__4252 (
            .O(N__19355),
            .I(N__19228));
    ClkMux I__4251 (
            .O(N__19354),
            .I(N__19228));
    ClkMux I__4250 (
            .O(N__19353),
            .I(N__19228));
    ClkMux I__4249 (
            .O(N__19352),
            .I(N__19228));
    ClkMux I__4248 (
            .O(N__19351),
            .I(N__19228));
    ClkMux I__4247 (
            .O(N__19350),
            .I(N__19228));
    ClkMux I__4246 (
            .O(N__19349),
            .I(N__19228));
    ClkMux I__4245 (
            .O(N__19348),
            .I(N__19228));
    ClkMux I__4244 (
            .O(N__19347),
            .I(N__19228));
    ClkMux I__4243 (
            .O(N__19346),
            .I(N__19228));
    ClkMux I__4242 (
            .O(N__19345),
            .I(N__19228));
    ClkMux I__4241 (
            .O(N__19344),
            .I(N__19228));
    ClkMux I__4240 (
            .O(N__19343),
            .I(N__19228));
    ClkMux I__4239 (
            .O(N__19342),
            .I(N__19228));
    ClkMux I__4238 (
            .O(N__19341),
            .I(N__19228));
    ClkMux I__4237 (
            .O(N__19340),
            .I(N__19228));
    ClkMux I__4236 (
            .O(N__19339),
            .I(N__19228));
    ClkMux I__4235 (
            .O(N__19338),
            .I(N__19228));
    ClkMux I__4234 (
            .O(N__19337),
            .I(N__19228));
    ClkMux I__4233 (
            .O(N__19336),
            .I(N__19228));
    ClkMux I__4232 (
            .O(N__19335),
            .I(N__19228));
    ClkMux I__4231 (
            .O(N__19334),
            .I(N__19228));
    ClkMux I__4230 (
            .O(N__19333),
            .I(N__19228));
    ClkMux I__4229 (
            .O(N__19332),
            .I(N__19228));
    ClkMux I__4228 (
            .O(N__19331),
            .I(N__19228));
    ClkMux I__4227 (
            .O(N__19330),
            .I(N__19228));
    ClkMux I__4226 (
            .O(N__19329),
            .I(N__19228));
    ClkMux I__4225 (
            .O(N__19328),
            .I(N__19228));
    ClkMux I__4224 (
            .O(N__19327),
            .I(N__19228));
    ClkMux I__4223 (
            .O(N__19326),
            .I(N__19228));
    ClkMux I__4222 (
            .O(N__19325),
            .I(N__19228));
    ClkMux I__4221 (
            .O(N__19324),
            .I(N__19228));
    ClkMux I__4220 (
            .O(N__19323),
            .I(N__19228));
    ClkMux I__4219 (
            .O(N__19322),
            .I(N__19228));
    ClkMux I__4218 (
            .O(N__19321),
            .I(N__19228));
    GlobalMux I__4217 (
            .O(N__19228),
            .I(N__19225));
    gio2CtrlBuf I__4216 (
            .O(N__19225),
            .I(DEBUG_c_1_c));
    IoInMux I__4215 (
            .O(N__19222),
            .I(N__19219));
    LocalMux I__4214 (
            .O(N__19219),
            .I(N__19216));
    Span12Mux_s6_h I__4213 (
            .O(N__19216),
            .I(N__19212));
    IoInMux I__4212 (
            .O(N__19215),
            .I(N__19209));
    Span12Mux_v I__4211 (
            .O(N__19212),
            .I(N__19206));
    LocalMux I__4210 (
            .O(N__19209),
            .I(N__19203));
    Span12Mux_v I__4209 (
            .O(N__19206),
            .I(N__19200));
    IoSpan4Mux I__4208 (
            .O(N__19203),
            .I(N__19197));
    Odrv12 I__4207 (
            .O(N__19200),
            .I(GB_BUFFER_DEBUG_c_1_c_THRU_CO));
    Odrv4 I__4206 (
            .O(N__19197),
            .I(GB_BUFFER_DEBUG_c_1_c_THRU_CO));
    InMux I__4205 (
            .O(N__19192),
            .I(N__19189));
    LocalMux I__4204 (
            .O(N__19189),
            .I(\transmit_module.Y_DELTA_PATTERN_29 ));
    InMux I__4203 (
            .O(N__19186),
            .I(N__19183));
    LocalMux I__4202 (
            .O(N__19183),
            .I(\transmit_module.Y_DELTA_PATTERN_31 ));
    InMux I__4201 (
            .O(N__19180),
            .I(N__19177));
    LocalMux I__4200 (
            .O(N__19177),
            .I(\transmit_module.Y_DELTA_PATTERN_30 ));
    CascadeMux I__4199 (
            .O(N__19174),
            .I(N__19171));
    InMux I__4198 (
            .O(N__19171),
            .I(N__19168));
    LocalMux I__4197 (
            .O(N__19168),
            .I(\transmit_module.n200 ));
    CascadeMux I__4196 (
            .O(N__19165),
            .I(\transmit_module.n215_cascade_ ));
    InMux I__4195 (
            .O(N__19162),
            .I(N__19159));
    LocalMux I__4194 (
            .O(N__19159),
            .I(\transmit_module.ADDR_Y_COMPONENT_5 ));
    InMux I__4193 (
            .O(N__19156),
            .I(N__19153));
    LocalMux I__4192 (
            .O(N__19153),
            .I(\transmit_module.n191 ));
    InMux I__4191 (
            .O(N__19150),
            .I(N__19147));
    LocalMux I__4190 (
            .O(N__19147),
            .I(N__19144));
    Span4Mux_v I__4189 (
            .O(N__19144),
            .I(N__19141));
    Odrv4 I__4188 (
            .O(N__19141),
            .I(\transmit_module.BRAM_ADDR_13_N_258_13 ));
    InMux I__4187 (
            .O(N__19138),
            .I(N__19135));
    LocalMux I__4186 (
            .O(N__19135),
            .I(N__19132));
    Odrv4 I__4185 (
            .O(N__19132),
            .I(\transmit_module.n199 ));
    InMux I__4184 (
            .O(N__19129),
            .I(N__19123));
    InMux I__4183 (
            .O(N__19128),
            .I(N__19117));
    InMux I__4182 (
            .O(N__19127),
            .I(N__19114));
    InMux I__4181 (
            .O(N__19126),
            .I(N__19111));
    LocalMux I__4180 (
            .O(N__19123),
            .I(N__19108));
    InMux I__4179 (
            .O(N__19122),
            .I(N__19105));
    CascadeMux I__4178 (
            .O(N__19121),
            .I(N__19096));
    InMux I__4177 (
            .O(N__19120),
            .I(N__19092));
    LocalMux I__4176 (
            .O(N__19117),
            .I(N__19089));
    LocalMux I__4175 (
            .O(N__19114),
            .I(N__19084));
    LocalMux I__4174 (
            .O(N__19111),
            .I(N__19084));
    Span4Mux_v I__4173 (
            .O(N__19108),
            .I(N__19079));
    LocalMux I__4172 (
            .O(N__19105),
            .I(N__19079));
    InMux I__4171 (
            .O(N__19104),
            .I(N__19076));
    InMux I__4170 (
            .O(N__19103),
            .I(N__19071));
    InMux I__4169 (
            .O(N__19102),
            .I(N__19071));
    InMux I__4168 (
            .O(N__19101),
            .I(N__19068));
    InMux I__4167 (
            .O(N__19100),
            .I(N__19065));
    InMux I__4166 (
            .O(N__19099),
            .I(N__19058));
    InMux I__4165 (
            .O(N__19096),
            .I(N__19058));
    InMux I__4164 (
            .O(N__19095),
            .I(N__19058));
    LocalMux I__4163 (
            .O(N__19092),
            .I(N__19053));
    Span4Mux_v I__4162 (
            .O(N__19089),
            .I(N__19053));
    Span4Mux_h I__4161 (
            .O(N__19084),
            .I(N__19042));
    Span4Mux_v I__4160 (
            .O(N__19079),
            .I(N__19042));
    LocalMux I__4159 (
            .O(N__19076),
            .I(N__19042));
    LocalMux I__4158 (
            .O(N__19071),
            .I(N__19042));
    LocalMux I__4157 (
            .O(N__19068),
            .I(N__19042));
    LocalMux I__4156 (
            .O(N__19065),
            .I(N__19037));
    LocalMux I__4155 (
            .O(N__19058),
            .I(N__19037));
    Odrv4 I__4154 (
            .O(N__19053),
            .I(\transmit_module.n3910 ));
    Odrv4 I__4153 (
            .O(N__19042),
            .I(\transmit_module.n3910 ));
    Odrv12 I__4152 (
            .O(N__19037),
            .I(\transmit_module.n3910 ));
    CascadeMux I__4151 (
            .O(N__19030),
            .I(\transmit_module.n214_cascade_ ));
    CascadeMux I__4150 (
            .O(N__19027),
            .I(N__19023));
    InMux I__4149 (
            .O(N__19026),
            .I(N__19018));
    InMux I__4148 (
            .O(N__19023),
            .I(N__19013));
    InMux I__4147 (
            .O(N__19022),
            .I(N__19013));
    InMux I__4146 (
            .O(N__19021),
            .I(N__19010));
    LocalMux I__4145 (
            .O(N__19018),
            .I(\transmit_module.TX_ADDR_5 ));
    LocalMux I__4144 (
            .O(N__19013),
            .I(\transmit_module.TX_ADDR_5 ));
    LocalMux I__4143 (
            .O(N__19010),
            .I(\transmit_module.TX_ADDR_5 ));
    InMux I__4142 (
            .O(N__19003),
            .I(N__19000));
    LocalMux I__4141 (
            .O(N__19000),
            .I(N__18997));
    Span4Mux_h I__4140 (
            .O(N__18997),
            .I(N__18994));
    Odrv4 I__4139 (
            .O(N__18994),
            .I(\transmit_module.ADDR_Y_COMPONENT_4 ));
    InMux I__4138 (
            .O(N__18991),
            .I(N__18988));
    LocalMux I__4137 (
            .O(N__18988),
            .I(N__18984));
    CascadeMux I__4136 (
            .O(N__18987),
            .I(N__18979));
    Span4Mux_v I__4135 (
            .O(N__18984),
            .I(N__18976));
    InMux I__4134 (
            .O(N__18983),
            .I(N__18971));
    InMux I__4133 (
            .O(N__18982),
            .I(N__18971));
    InMux I__4132 (
            .O(N__18979),
            .I(N__18968));
    Odrv4 I__4131 (
            .O(N__18976),
            .I(\transmit_module.TX_ADDR_4 ));
    LocalMux I__4130 (
            .O(N__18971),
            .I(\transmit_module.TX_ADDR_4 ));
    LocalMux I__4129 (
            .O(N__18968),
            .I(\transmit_module.TX_ADDR_4 ));
    InMux I__4128 (
            .O(N__18961),
            .I(N__18957));
    InMux I__4127 (
            .O(N__18960),
            .I(N__18954));
    LocalMux I__4126 (
            .O(N__18957),
            .I(\transmit_module.n184 ));
    LocalMux I__4125 (
            .O(N__18954),
            .I(\transmit_module.n184 ));
    InMux I__4124 (
            .O(N__18949),
            .I(N__18946));
    LocalMux I__4123 (
            .O(N__18946),
            .I(\transmit_module.n215 ));
    CascadeMux I__4122 (
            .O(N__18943),
            .I(N__18939));
    CascadeMux I__4121 (
            .O(N__18942),
            .I(N__18936));
    CascadeBuf I__4120 (
            .O(N__18939),
            .I(N__18933));
    CascadeBuf I__4119 (
            .O(N__18936),
            .I(N__18930));
    CascadeMux I__4118 (
            .O(N__18933),
            .I(N__18927));
    CascadeMux I__4117 (
            .O(N__18930),
            .I(N__18924));
    CascadeBuf I__4116 (
            .O(N__18927),
            .I(N__18921));
    CascadeBuf I__4115 (
            .O(N__18924),
            .I(N__18918));
    CascadeMux I__4114 (
            .O(N__18921),
            .I(N__18915));
    CascadeMux I__4113 (
            .O(N__18918),
            .I(N__18912));
    CascadeBuf I__4112 (
            .O(N__18915),
            .I(N__18909));
    CascadeBuf I__4111 (
            .O(N__18912),
            .I(N__18906));
    CascadeMux I__4110 (
            .O(N__18909),
            .I(N__18903));
    CascadeMux I__4109 (
            .O(N__18906),
            .I(N__18900));
    CascadeBuf I__4108 (
            .O(N__18903),
            .I(N__18897));
    CascadeBuf I__4107 (
            .O(N__18900),
            .I(N__18894));
    CascadeMux I__4106 (
            .O(N__18897),
            .I(N__18891));
    CascadeMux I__4105 (
            .O(N__18894),
            .I(N__18888));
    CascadeBuf I__4104 (
            .O(N__18891),
            .I(N__18885));
    CascadeBuf I__4103 (
            .O(N__18888),
            .I(N__18882));
    CascadeMux I__4102 (
            .O(N__18885),
            .I(N__18879));
    CascadeMux I__4101 (
            .O(N__18882),
            .I(N__18876));
    CascadeBuf I__4100 (
            .O(N__18879),
            .I(N__18873));
    CascadeBuf I__4099 (
            .O(N__18876),
            .I(N__18870));
    CascadeMux I__4098 (
            .O(N__18873),
            .I(N__18867));
    CascadeMux I__4097 (
            .O(N__18870),
            .I(N__18864));
    CascadeBuf I__4096 (
            .O(N__18867),
            .I(N__18861));
    CascadeBuf I__4095 (
            .O(N__18864),
            .I(N__18858));
    CascadeMux I__4094 (
            .O(N__18861),
            .I(N__18855));
    CascadeMux I__4093 (
            .O(N__18858),
            .I(N__18852));
    CascadeBuf I__4092 (
            .O(N__18855),
            .I(N__18849));
    CascadeBuf I__4091 (
            .O(N__18852),
            .I(N__18846));
    CascadeMux I__4090 (
            .O(N__18849),
            .I(N__18843));
    CascadeMux I__4089 (
            .O(N__18846),
            .I(N__18840));
    CascadeBuf I__4088 (
            .O(N__18843),
            .I(N__18837));
    CascadeBuf I__4087 (
            .O(N__18840),
            .I(N__18834));
    CascadeMux I__4086 (
            .O(N__18837),
            .I(N__18831));
    CascadeMux I__4085 (
            .O(N__18834),
            .I(N__18828));
    CascadeBuf I__4084 (
            .O(N__18831),
            .I(N__18825));
    CascadeBuf I__4083 (
            .O(N__18828),
            .I(N__18822));
    CascadeMux I__4082 (
            .O(N__18825),
            .I(N__18819));
    CascadeMux I__4081 (
            .O(N__18822),
            .I(N__18816));
    CascadeBuf I__4080 (
            .O(N__18819),
            .I(N__18813));
    CascadeBuf I__4079 (
            .O(N__18816),
            .I(N__18810));
    CascadeMux I__4078 (
            .O(N__18813),
            .I(N__18807));
    CascadeMux I__4077 (
            .O(N__18810),
            .I(N__18804));
    CascadeBuf I__4076 (
            .O(N__18807),
            .I(N__18801));
    CascadeBuf I__4075 (
            .O(N__18804),
            .I(N__18798));
    CascadeMux I__4074 (
            .O(N__18801),
            .I(N__18795));
    CascadeMux I__4073 (
            .O(N__18798),
            .I(N__18792));
    CascadeBuf I__4072 (
            .O(N__18795),
            .I(N__18789));
    CascadeBuf I__4071 (
            .O(N__18792),
            .I(N__18786));
    CascadeMux I__4070 (
            .O(N__18789),
            .I(N__18783));
    CascadeMux I__4069 (
            .O(N__18786),
            .I(N__18780));
    CascadeBuf I__4068 (
            .O(N__18783),
            .I(N__18777));
    CascadeBuf I__4067 (
            .O(N__18780),
            .I(N__18774));
    CascadeMux I__4066 (
            .O(N__18777),
            .I(N__18771));
    CascadeMux I__4065 (
            .O(N__18774),
            .I(N__18768));
    CascadeBuf I__4064 (
            .O(N__18771),
            .I(N__18765));
    CascadeBuf I__4063 (
            .O(N__18768),
            .I(N__18762));
    CascadeMux I__4062 (
            .O(N__18765),
            .I(N__18759));
    CascadeMux I__4061 (
            .O(N__18762),
            .I(N__18756));
    InMux I__4060 (
            .O(N__18759),
            .I(N__18753));
    InMux I__4059 (
            .O(N__18756),
            .I(N__18750));
    LocalMux I__4058 (
            .O(N__18753),
            .I(N__18747));
    LocalMux I__4057 (
            .O(N__18750),
            .I(N__18744));
    Span12Mux_h I__4056 (
            .O(N__18747),
            .I(N__18739));
    Span12Mux_h I__4055 (
            .O(N__18744),
            .I(N__18739));
    Span12Mux_v I__4054 (
            .O(N__18739),
            .I(N__18736));
    Odrv12 I__4053 (
            .O(N__18736),
            .I(n24));
    CascadeMux I__4052 (
            .O(N__18733),
            .I(N__18729));
    InMux I__4051 (
            .O(N__18732),
            .I(N__18726));
    InMux I__4050 (
            .O(N__18729),
            .I(N__18723));
    LocalMux I__4049 (
            .O(N__18726),
            .I(\transmit_module.n183 ));
    LocalMux I__4048 (
            .O(N__18723),
            .I(\transmit_module.n183 ));
    InMux I__4047 (
            .O(N__18718),
            .I(N__18715));
    LocalMux I__4046 (
            .O(N__18715),
            .I(\transmit_module.n214 ));
    CascadeMux I__4045 (
            .O(N__18712),
            .I(N__18708));
    CascadeMux I__4044 (
            .O(N__18711),
            .I(N__18705));
    CascadeBuf I__4043 (
            .O(N__18708),
            .I(N__18702));
    CascadeBuf I__4042 (
            .O(N__18705),
            .I(N__18699));
    CascadeMux I__4041 (
            .O(N__18702),
            .I(N__18696));
    CascadeMux I__4040 (
            .O(N__18699),
            .I(N__18693));
    CascadeBuf I__4039 (
            .O(N__18696),
            .I(N__18690));
    CascadeBuf I__4038 (
            .O(N__18693),
            .I(N__18687));
    CascadeMux I__4037 (
            .O(N__18690),
            .I(N__18684));
    CascadeMux I__4036 (
            .O(N__18687),
            .I(N__18681));
    CascadeBuf I__4035 (
            .O(N__18684),
            .I(N__18678));
    CascadeBuf I__4034 (
            .O(N__18681),
            .I(N__18675));
    CascadeMux I__4033 (
            .O(N__18678),
            .I(N__18672));
    CascadeMux I__4032 (
            .O(N__18675),
            .I(N__18669));
    CascadeBuf I__4031 (
            .O(N__18672),
            .I(N__18666));
    CascadeBuf I__4030 (
            .O(N__18669),
            .I(N__18663));
    CascadeMux I__4029 (
            .O(N__18666),
            .I(N__18660));
    CascadeMux I__4028 (
            .O(N__18663),
            .I(N__18657));
    CascadeBuf I__4027 (
            .O(N__18660),
            .I(N__18654));
    CascadeBuf I__4026 (
            .O(N__18657),
            .I(N__18651));
    CascadeMux I__4025 (
            .O(N__18654),
            .I(N__18648));
    CascadeMux I__4024 (
            .O(N__18651),
            .I(N__18645));
    CascadeBuf I__4023 (
            .O(N__18648),
            .I(N__18642));
    CascadeBuf I__4022 (
            .O(N__18645),
            .I(N__18639));
    CascadeMux I__4021 (
            .O(N__18642),
            .I(N__18636));
    CascadeMux I__4020 (
            .O(N__18639),
            .I(N__18633));
    CascadeBuf I__4019 (
            .O(N__18636),
            .I(N__18630));
    CascadeBuf I__4018 (
            .O(N__18633),
            .I(N__18627));
    CascadeMux I__4017 (
            .O(N__18630),
            .I(N__18624));
    CascadeMux I__4016 (
            .O(N__18627),
            .I(N__18621));
    CascadeBuf I__4015 (
            .O(N__18624),
            .I(N__18618));
    CascadeBuf I__4014 (
            .O(N__18621),
            .I(N__18615));
    CascadeMux I__4013 (
            .O(N__18618),
            .I(N__18612));
    CascadeMux I__4012 (
            .O(N__18615),
            .I(N__18609));
    CascadeBuf I__4011 (
            .O(N__18612),
            .I(N__18606));
    CascadeBuf I__4010 (
            .O(N__18609),
            .I(N__18603));
    CascadeMux I__4009 (
            .O(N__18606),
            .I(N__18600));
    CascadeMux I__4008 (
            .O(N__18603),
            .I(N__18597));
    CascadeBuf I__4007 (
            .O(N__18600),
            .I(N__18594));
    CascadeBuf I__4006 (
            .O(N__18597),
            .I(N__18591));
    CascadeMux I__4005 (
            .O(N__18594),
            .I(N__18588));
    CascadeMux I__4004 (
            .O(N__18591),
            .I(N__18585));
    CascadeBuf I__4003 (
            .O(N__18588),
            .I(N__18582));
    CascadeBuf I__4002 (
            .O(N__18585),
            .I(N__18579));
    CascadeMux I__4001 (
            .O(N__18582),
            .I(N__18576));
    CascadeMux I__4000 (
            .O(N__18579),
            .I(N__18573));
    CascadeBuf I__3999 (
            .O(N__18576),
            .I(N__18570));
    CascadeBuf I__3998 (
            .O(N__18573),
            .I(N__18567));
    CascadeMux I__3997 (
            .O(N__18570),
            .I(N__18564));
    CascadeMux I__3996 (
            .O(N__18567),
            .I(N__18561));
    CascadeBuf I__3995 (
            .O(N__18564),
            .I(N__18558));
    CascadeBuf I__3994 (
            .O(N__18561),
            .I(N__18555));
    CascadeMux I__3993 (
            .O(N__18558),
            .I(N__18552));
    CascadeMux I__3992 (
            .O(N__18555),
            .I(N__18549));
    CascadeBuf I__3991 (
            .O(N__18552),
            .I(N__18546));
    CascadeBuf I__3990 (
            .O(N__18549),
            .I(N__18543));
    CascadeMux I__3989 (
            .O(N__18546),
            .I(N__18540));
    CascadeMux I__3988 (
            .O(N__18543),
            .I(N__18537));
    CascadeBuf I__3987 (
            .O(N__18540),
            .I(N__18534));
    CascadeBuf I__3986 (
            .O(N__18537),
            .I(N__18531));
    CascadeMux I__3985 (
            .O(N__18534),
            .I(N__18528));
    CascadeMux I__3984 (
            .O(N__18531),
            .I(N__18525));
    InMux I__3983 (
            .O(N__18528),
            .I(N__18522));
    InMux I__3982 (
            .O(N__18525),
            .I(N__18519));
    LocalMux I__3981 (
            .O(N__18522),
            .I(N__18516));
    LocalMux I__3980 (
            .O(N__18519),
            .I(N__18513));
    Span12Mux_h I__3979 (
            .O(N__18516),
            .I(N__18510));
    Span12Mux_v I__3978 (
            .O(N__18513),
            .I(N__18507));
    Span12Mux_v I__3977 (
            .O(N__18510),
            .I(N__18504));
    Odrv12 I__3976 (
            .O(N__18507),
            .I(n23));
    Odrv12 I__3975 (
            .O(N__18504),
            .I(n23));
    InMux I__3974 (
            .O(N__18499),
            .I(N__18496));
    LocalMux I__3973 (
            .O(N__18496),
            .I(\transmit_module.Y_DELTA_PATTERN_18 ));
    InMux I__3972 (
            .O(N__18493),
            .I(N__18490));
    LocalMux I__3971 (
            .O(N__18490),
            .I(\transmit_module.Y_DELTA_PATTERN_21 ));
    InMux I__3970 (
            .O(N__18487),
            .I(N__18484));
    LocalMux I__3969 (
            .O(N__18484),
            .I(\transmit_module.Y_DELTA_PATTERN_20 ));
    InMux I__3968 (
            .O(N__18481),
            .I(N__18478));
    LocalMux I__3967 (
            .O(N__18478),
            .I(\transmit_module.Y_DELTA_PATTERN_19 ));
    InMux I__3966 (
            .O(N__18475),
            .I(N__18472));
    LocalMux I__3965 (
            .O(N__18472),
            .I(\transmit_module.Y_DELTA_PATTERN_1 ));
    InMux I__3964 (
            .O(N__18469),
            .I(N__18466));
    LocalMux I__3963 (
            .O(N__18466),
            .I(N__18461));
    CascadeMux I__3962 (
            .O(N__18465),
            .I(N__18458));
    CascadeMux I__3961 (
            .O(N__18464),
            .I(N__18454));
    Span4Mux_h I__3960 (
            .O(N__18461),
            .I(N__18451));
    InMux I__3959 (
            .O(N__18458),
            .I(N__18448));
    InMux I__3958 (
            .O(N__18457),
            .I(N__18445));
    InMux I__3957 (
            .O(N__18454),
            .I(N__18442));
    Odrv4 I__3956 (
            .O(N__18451),
            .I(\transmit_module.TX_ADDR_9 ));
    LocalMux I__3955 (
            .O(N__18448),
            .I(\transmit_module.TX_ADDR_9 ));
    LocalMux I__3954 (
            .O(N__18445),
            .I(\transmit_module.TX_ADDR_9 ));
    LocalMux I__3953 (
            .O(N__18442),
            .I(\transmit_module.TX_ADDR_9 ));
    InMux I__3952 (
            .O(N__18433),
            .I(N__18430));
    LocalMux I__3951 (
            .O(N__18430),
            .I(N__18427));
    Span4Mux_h I__3950 (
            .O(N__18427),
            .I(N__18424));
    Odrv4 I__3949 (
            .O(N__18424),
            .I(\transmit_module.ADDR_Y_COMPONENT_9 ));
    InMux I__3948 (
            .O(N__18421),
            .I(N__18417));
    InMux I__3947 (
            .O(N__18420),
            .I(N__18414));
    LocalMux I__3946 (
            .O(N__18417),
            .I(N__18411));
    LocalMux I__3945 (
            .O(N__18414),
            .I(N__18408));
    Span4Mux_v I__3944 (
            .O(N__18411),
            .I(N__18403));
    Span4Mux_h I__3943 (
            .O(N__18408),
            .I(N__18400));
    InMux I__3942 (
            .O(N__18407),
            .I(N__18397));
    InMux I__3941 (
            .O(N__18406),
            .I(N__18394));
    Odrv4 I__3940 (
            .O(N__18403),
            .I(\transmit_module.TX_ADDR_0 ));
    Odrv4 I__3939 (
            .O(N__18400),
            .I(\transmit_module.TX_ADDR_0 ));
    LocalMux I__3938 (
            .O(N__18397),
            .I(\transmit_module.TX_ADDR_0 ));
    LocalMux I__3937 (
            .O(N__18394),
            .I(\transmit_module.TX_ADDR_0 ));
    InMux I__3936 (
            .O(N__18385),
            .I(N__18382));
    LocalMux I__3935 (
            .O(N__18382),
            .I(\transmit_module.ADDR_Y_COMPONENT_0 ));
    InMux I__3934 (
            .O(N__18379),
            .I(N__18376));
    LocalMux I__3933 (
            .O(N__18376),
            .I(N__18370));
    InMux I__3932 (
            .O(N__18375),
            .I(N__18367));
    InMux I__3931 (
            .O(N__18374),
            .I(N__18364));
    InMux I__3930 (
            .O(N__18373),
            .I(N__18361));
    Odrv4 I__3929 (
            .O(N__18370),
            .I(\transmit_module.TX_ADDR_3 ));
    LocalMux I__3928 (
            .O(N__18367),
            .I(\transmit_module.TX_ADDR_3 ));
    LocalMux I__3927 (
            .O(N__18364),
            .I(\transmit_module.TX_ADDR_3 ));
    LocalMux I__3926 (
            .O(N__18361),
            .I(\transmit_module.TX_ADDR_3 ));
    InMux I__3925 (
            .O(N__18352),
            .I(N__18349));
    LocalMux I__3924 (
            .O(N__18349),
            .I(\transmit_module.ADDR_Y_COMPONENT_3 ));
    InMux I__3923 (
            .O(N__18346),
            .I(N__18343));
    LocalMux I__3922 (
            .O(N__18343),
            .I(N__18340));
    Odrv4 I__3921 (
            .O(N__18340),
            .I(\transmit_module.n193 ));
    CascadeMux I__3920 (
            .O(N__18337),
            .I(N__18334));
    InMux I__3919 (
            .O(N__18334),
            .I(N__18331));
    LocalMux I__3918 (
            .O(N__18331),
            .I(\transmit_module.ADDR_Y_COMPONENT_11 ));
    InMux I__3917 (
            .O(N__18328),
            .I(N__18325));
    LocalMux I__3916 (
            .O(N__18325),
            .I(\transmit_module.ADDR_Y_COMPONENT_1 ));
    InMux I__3915 (
            .O(N__18322),
            .I(N__18316));
    InMux I__3914 (
            .O(N__18321),
            .I(N__18313));
    InMux I__3913 (
            .O(N__18320),
            .I(N__18310));
    InMux I__3912 (
            .O(N__18319),
            .I(N__18307));
    LocalMux I__3911 (
            .O(N__18316),
            .I(N__18302));
    LocalMux I__3910 (
            .O(N__18313),
            .I(N__18302));
    LocalMux I__3909 (
            .O(N__18310),
            .I(N__18299));
    LocalMux I__3908 (
            .O(N__18307),
            .I(\transmit_module.TX_ADDR_1 ));
    Odrv4 I__3907 (
            .O(N__18302),
            .I(\transmit_module.TX_ADDR_1 ));
    Odrv4 I__3906 (
            .O(N__18299),
            .I(\transmit_module.TX_ADDR_1 ));
    InMux I__3905 (
            .O(N__18292),
            .I(N__18288));
    InMux I__3904 (
            .O(N__18291),
            .I(N__18285));
    LocalMux I__3903 (
            .O(N__18288),
            .I(N__18282));
    LocalMux I__3902 (
            .O(N__18285),
            .I(N__18279));
    Odrv4 I__3901 (
            .O(N__18282),
            .I(\transmit_module.n187 ));
    Odrv12 I__3900 (
            .O(N__18279),
            .I(\transmit_module.n187 ));
    InMux I__3899 (
            .O(N__18274),
            .I(N__18271));
    LocalMux I__3898 (
            .O(N__18271),
            .I(N__18268));
    Odrv12 I__3897 (
            .O(N__18268),
            .I(\transmit_module.n218 ));
    CascadeMux I__3896 (
            .O(N__18265),
            .I(N__18262));
    CascadeBuf I__3895 (
            .O(N__18262),
            .I(N__18258));
    CascadeMux I__3894 (
            .O(N__18261),
            .I(N__18255));
    CascadeMux I__3893 (
            .O(N__18258),
            .I(N__18252));
    CascadeBuf I__3892 (
            .O(N__18255),
            .I(N__18249));
    CascadeBuf I__3891 (
            .O(N__18252),
            .I(N__18246));
    CascadeMux I__3890 (
            .O(N__18249),
            .I(N__18243));
    CascadeMux I__3889 (
            .O(N__18246),
            .I(N__18240));
    CascadeBuf I__3888 (
            .O(N__18243),
            .I(N__18237));
    CascadeBuf I__3887 (
            .O(N__18240),
            .I(N__18234));
    CascadeMux I__3886 (
            .O(N__18237),
            .I(N__18231));
    CascadeMux I__3885 (
            .O(N__18234),
            .I(N__18228));
    CascadeBuf I__3884 (
            .O(N__18231),
            .I(N__18225));
    CascadeBuf I__3883 (
            .O(N__18228),
            .I(N__18222));
    CascadeMux I__3882 (
            .O(N__18225),
            .I(N__18219));
    CascadeMux I__3881 (
            .O(N__18222),
            .I(N__18216));
    CascadeBuf I__3880 (
            .O(N__18219),
            .I(N__18213));
    CascadeBuf I__3879 (
            .O(N__18216),
            .I(N__18210));
    CascadeMux I__3878 (
            .O(N__18213),
            .I(N__18207));
    CascadeMux I__3877 (
            .O(N__18210),
            .I(N__18204));
    CascadeBuf I__3876 (
            .O(N__18207),
            .I(N__18201));
    CascadeBuf I__3875 (
            .O(N__18204),
            .I(N__18198));
    CascadeMux I__3874 (
            .O(N__18201),
            .I(N__18195));
    CascadeMux I__3873 (
            .O(N__18198),
            .I(N__18192));
    CascadeBuf I__3872 (
            .O(N__18195),
            .I(N__18189));
    CascadeBuf I__3871 (
            .O(N__18192),
            .I(N__18186));
    CascadeMux I__3870 (
            .O(N__18189),
            .I(N__18183));
    CascadeMux I__3869 (
            .O(N__18186),
            .I(N__18180));
    CascadeBuf I__3868 (
            .O(N__18183),
            .I(N__18177));
    CascadeBuf I__3867 (
            .O(N__18180),
            .I(N__18174));
    CascadeMux I__3866 (
            .O(N__18177),
            .I(N__18171));
    CascadeMux I__3865 (
            .O(N__18174),
            .I(N__18168));
    CascadeBuf I__3864 (
            .O(N__18171),
            .I(N__18165));
    CascadeBuf I__3863 (
            .O(N__18168),
            .I(N__18162));
    CascadeMux I__3862 (
            .O(N__18165),
            .I(N__18159));
    CascadeMux I__3861 (
            .O(N__18162),
            .I(N__18156));
    CascadeBuf I__3860 (
            .O(N__18159),
            .I(N__18153));
    CascadeBuf I__3859 (
            .O(N__18156),
            .I(N__18150));
    CascadeMux I__3858 (
            .O(N__18153),
            .I(N__18147));
    CascadeMux I__3857 (
            .O(N__18150),
            .I(N__18144));
    CascadeBuf I__3856 (
            .O(N__18147),
            .I(N__18141));
    CascadeBuf I__3855 (
            .O(N__18144),
            .I(N__18138));
    CascadeMux I__3854 (
            .O(N__18141),
            .I(N__18135));
    CascadeMux I__3853 (
            .O(N__18138),
            .I(N__18132));
    CascadeBuf I__3852 (
            .O(N__18135),
            .I(N__18129));
    CascadeBuf I__3851 (
            .O(N__18132),
            .I(N__18126));
    CascadeMux I__3850 (
            .O(N__18129),
            .I(N__18123));
    CascadeMux I__3849 (
            .O(N__18126),
            .I(N__18120));
    CascadeBuf I__3848 (
            .O(N__18123),
            .I(N__18117));
    CascadeBuf I__3847 (
            .O(N__18120),
            .I(N__18114));
    CascadeMux I__3846 (
            .O(N__18117),
            .I(N__18111));
    CascadeMux I__3845 (
            .O(N__18114),
            .I(N__18108));
    CascadeBuf I__3844 (
            .O(N__18111),
            .I(N__18105));
    CascadeBuf I__3843 (
            .O(N__18108),
            .I(N__18102));
    CascadeMux I__3842 (
            .O(N__18105),
            .I(N__18099));
    CascadeMux I__3841 (
            .O(N__18102),
            .I(N__18096));
    CascadeBuf I__3840 (
            .O(N__18099),
            .I(N__18093));
    CascadeBuf I__3839 (
            .O(N__18096),
            .I(N__18090));
    CascadeMux I__3838 (
            .O(N__18093),
            .I(N__18087));
    CascadeMux I__3837 (
            .O(N__18090),
            .I(N__18084));
    CascadeBuf I__3836 (
            .O(N__18087),
            .I(N__18081));
    InMux I__3835 (
            .O(N__18084),
            .I(N__18078));
    CascadeMux I__3834 (
            .O(N__18081),
            .I(N__18075));
    LocalMux I__3833 (
            .O(N__18078),
            .I(N__18072));
    InMux I__3832 (
            .O(N__18075),
            .I(N__18069));
    Span4Mux_v I__3831 (
            .O(N__18072),
            .I(N__18066));
    LocalMux I__3830 (
            .O(N__18069),
            .I(N__18063));
    Span4Mux_h I__3829 (
            .O(N__18066),
            .I(N__18060));
    Span4Mux_v I__3828 (
            .O(N__18063),
            .I(N__18057));
    Span4Mux_h I__3827 (
            .O(N__18060),
            .I(N__18052));
    Span4Mux_h I__3826 (
            .O(N__18057),
            .I(N__18052));
    Odrv4 I__3825 (
            .O(N__18052),
            .I(n27));
    InMux I__3824 (
            .O(N__18049),
            .I(N__18046));
    LocalMux I__3823 (
            .O(N__18046),
            .I(N__18043));
    Span4Mux_h I__3822 (
            .O(N__18043),
            .I(N__18040));
    Sp12to4 I__3821 (
            .O(N__18040),
            .I(N__18037));
    Span12Mux_v I__3820 (
            .O(N__18037),
            .I(N__18034));
    Odrv12 I__3819 (
            .O(N__18034),
            .I(\line_buffer.n678 ));
    CascadeMux I__3818 (
            .O(N__18031),
            .I(N__18028));
    InMux I__3817 (
            .O(N__18028),
            .I(N__18025));
    LocalMux I__3816 (
            .O(N__18025),
            .I(N__18022));
    Odrv12 I__3815 (
            .O(N__18022),
            .I(\line_buffer.n686 ));
    InMux I__3814 (
            .O(N__18019),
            .I(N__18016));
    LocalMux I__3813 (
            .O(N__18016),
            .I(N__18013));
    Span4Mux_v I__3812 (
            .O(N__18013),
            .I(N__18010));
    Span4Mux_h I__3811 (
            .O(N__18010),
            .I(N__18007));
    Span4Mux_h I__3810 (
            .O(N__18007),
            .I(N__18004));
    Odrv4 I__3809 (
            .O(N__18004),
            .I(\line_buffer.n614 ));
    CascadeMux I__3808 (
            .O(N__18001),
            .I(\line_buffer.n4188_cascade_ ));
    InMux I__3807 (
            .O(N__17998),
            .I(N__17995));
    LocalMux I__3806 (
            .O(N__17995),
            .I(N__17992));
    Span4Mux_h I__3805 (
            .O(N__17992),
            .I(N__17989));
    Sp12to4 I__3804 (
            .O(N__17989),
            .I(N__17986));
    Span12Mux_v I__3803 (
            .O(N__17986),
            .I(N__17983));
    Odrv12 I__3802 (
            .O(N__17983),
            .I(\line_buffer.n622 ));
    CascadeMux I__3801 (
            .O(N__17980),
            .I(\line_buffer.n4191_cascade_ ));
    InMux I__3800 (
            .O(N__17977),
            .I(N__17974));
    LocalMux I__3799 (
            .O(N__17974),
            .I(\line_buffer.n4179 ));
    InMux I__3798 (
            .O(N__17971),
            .I(N__17968));
    LocalMux I__3797 (
            .O(N__17968),
            .I(N__17965));
    Span4Mux_h I__3796 (
            .O(N__17965),
            .I(N__17962));
    Span4Mux_v I__3795 (
            .O(N__17962),
            .I(N__17959));
    Odrv4 I__3794 (
            .O(N__17959),
            .I(TX_DATA_5));
    InMux I__3793 (
            .O(N__17956),
            .I(N__17952));
    CascadeMux I__3792 (
            .O(N__17955),
            .I(N__17948));
    LocalMux I__3791 (
            .O(N__17952),
            .I(N__17945));
    InMux I__3790 (
            .O(N__17951),
            .I(N__17941));
    InMux I__3789 (
            .O(N__17948),
            .I(N__17938));
    Span4Mux_h I__3788 (
            .O(N__17945),
            .I(N__17935));
    InMux I__3787 (
            .O(N__17944),
            .I(N__17932));
    LocalMux I__3786 (
            .O(N__17941),
            .I(N__17925));
    LocalMux I__3785 (
            .O(N__17938),
            .I(N__17925));
    Span4Mux_v I__3784 (
            .O(N__17935),
            .I(N__17925));
    LocalMux I__3783 (
            .O(N__17932),
            .I(\transmit_module.TX_ADDR_10 ));
    Odrv4 I__3782 (
            .O(N__17925),
            .I(\transmit_module.TX_ADDR_10 ));
    InMux I__3781 (
            .O(N__17920),
            .I(N__17917));
    LocalMux I__3780 (
            .O(N__17917),
            .I(N__17914));
    Span4Mux_v I__3779 (
            .O(N__17914),
            .I(N__17911));
    Span4Mux_v I__3778 (
            .O(N__17911),
            .I(N__17908));
    Odrv4 I__3777 (
            .O(N__17908),
            .I(\transmit_module.n194 ));
    InMux I__3776 (
            .O(N__17905),
            .I(\transmit_module.n3665 ));
    InMux I__3775 (
            .O(N__17902),
            .I(\transmit_module.n3666 ));
    InMux I__3774 (
            .O(N__17899),
            .I(\transmit_module.n3667 ));
    InMux I__3773 (
            .O(N__17896),
            .I(\transmit_module.n3668 ));
    CascadeMux I__3772 (
            .O(N__17893),
            .I(N__17890));
    InMux I__3771 (
            .O(N__17890),
            .I(N__17887));
    LocalMux I__3770 (
            .O(N__17887),
            .I(N__17881));
    InMux I__3769 (
            .O(N__17886),
            .I(N__17878));
    InMux I__3768 (
            .O(N__17885),
            .I(N__17873));
    InMux I__3767 (
            .O(N__17884),
            .I(N__17873));
    Odrv4 I__3766 (
            .O(N__17881),
            .I(\transmit_module.TX_ADDR_8 ));
    LocalMux I__3765 (
            .O(N__17878),
            .I(\transmit_module.TX_ADDR_8 ));
    LocalMux I__3764 (
            .O(N__17873),
            .I(\transmit_module.TX_ADDR_8 ));
    InMux I__3763 (
            .O(N__17866),
            .I(N__17863));
    LocalMux I__3762 (
            .O(N__17863),
            .I(N__17860));
    Span4Mux_h I__3761 (
            .O(N__17860),
            .I(N__17857));
    Odrv4 I__3760 (
            .O(N__17857),
            .I(\transmit_module.ADDR_Y_COMPONENT_8 ));
    CascadeMux I__3759 (
            .O(N__17854),
            .I(N__17851));
    InMux I__3758 (
            .O(N__17851),
            .I(N__17848));
    LocalMux I__3757 (
            .O(N__17848),
            .I(N__17845));
    Odrv4 I__3756 (
            .O(N__17845),
            .I(\transmit_module.n203 ));
    CascadeMux I__3755 (
            .O(N__17842),
            .I(\transmit_module.n218_cascade_ ));
    InMux I__3754 (
            .O(N__17839),
            .I(N__17835));
    InMux I__3753 (
            .O(N__17838),
            .I(N__17832));
    LocalMux I__3752 (
            .O(N__17835),
            .I(N__17829));
    LocalMux I__3751 (
            .O(N__17832),
            .I(\transmit_module.n188 ));
    Odrv12 I__3750 (
            .O(N__17829),
            .I(\transmit_module.n188 ));
    InMux I__3749 (
            .O(N__17824),
            .I(N__17818));
    InMux I__3748 (
            .O(N__17823),
            .I(N__17815));
    InMux I__3747 (
            .O(N__17822),
            .I(N__17812));
    InMux I__3746 (
            .O(N__17821),
            .I(N__17809));
    LocalMux I__3745 (
            .O(N__17818),
            .I(N__17804));
    LocalMux I__3744 (
            .O(N__17815),
            .I(N__17804));
    LocalMux I__3743 (
            .O(N__17812),
            .I(\transmit_module.TX_ADDR_2 ));
    LocalMux I__3742 (
            .O(N__17809),
            .I(\transmit_module.TX_ADDR_2 ));
    Odrv4 I__3741 (
            .O(N__17804),
            .I(\transmit_module.TX_ADDR_2 ));
    InMux I__3740 (
            .O(N__17797),
            .I(N__17794));
    LocalMux I__3739 (
            .O(N__17794),
            .I(N__17791));
    Span4Mux_h I__3738 (
            .O(N__17791),
            .I(N__17788));
    Odrv4 I__3737 (
            .O(N__17788),
            .I(\transmit_module.n202 ));
    InMux I__3736 (
            .O(N__17785),
            .I(\transmit_module.n3657 ));
    CascadeMux I__3735 (
            .O(N__17782),
            .I(N__17779));
    InMux I__3734 (
            .O(N__17779),
            .I(N__17776));
    LocalMux I__3733 (
            .O(N__17776),
            .I(N__17773));
    Span4Mux_v I__3732 (
            .O(N__17773),
            .I(N__17770));
    Odrv4 I__3731 (
            .O(N__17770),
            .I(\transmit_module.n201 ));
    InMux I__3730 (
            .O(N__17767),
            .I(\transmit_module.n3658 ));
    InMux I__3729 (
            .O(N__17764),
            .I(\transmit_module.n3659 ));
    InMux I__3728 (
            .O(N__17761),
            .I(\transmit_module.n3660 ));
    InMux I__3727 (
            .O(N__17758),
            .I(N__17753));
    InMux I__3726 (
            .O(N__17757),
            .I(N__17750));
    CascadeMux I__3725 (
            .O(N__17756),
            .I(N__17747));
    LocalMux I__3724 (
            .O(N__17753),
            .I(N__17742));
    LocalMux I__3723 (
            .O(N__17750),
            .I(N__17742));
    InMux I__3722 (
            .O(N__17747),
            .I(N__17738));
    Span4Mux_v I__3721 (
            .O(N__17742),
            .I(N__17735));
    InMux I__3720 (
            .O(N__17741),
            .I(N__17732));
    LocalMux I__3719 (
            .O(N__17738),
            .I(\transmit_module.TX_ADDR_6 ));
    Odrv4 I__3718 (
            .O(N__17735),
            .I(\transmit_module.TX_ADDR_6 ));
    LocalMux I__3717 (
            .O(N__17732),
            .I(\transmit_module.TX_ADDR_6 ));
    InMux I__3716 (
            .O(N__17725),
            .I(N__17722));
    LocalMux I__3715 (
            .O(N__17722),
            .I(N__17719));
    Odrv4 I__3714 (
            .O(N__17719),
            .I(\transmit_module.n198 ));
    InMux I__3713 (
            .O(N__17716),
            .I(\transmit_module.n3661 ));
    InMux I__3712 (
            .O(N__17713),
            .I(N__17709));
    CascadeMux I__3711 (
            .O(N__17712),
            .I(N__17705));
    LocalMux I__3710 (
            .O(N__17709),
            .I(N__17701));
    InMux I__3709 (
            .O(N__17708),
            .I(N__17698));
    InMux I__3708 (
            .O(N__17705),
            .I(N__17695));
    InMux I__3707 (
            .O(N__17704),
            .I(N__17692));
    Odrv4 I__3706 (
            .O(N__17701),
            .I(\transmit_module.TX_ADDR_7 ));
    LocalMux I__3705 (
            .O(N__17698),
            .I(\transmit_module.TX_ADDR_7 ));
    LocalMux I__3704 (
            .O(N__17695),
            .I(\transmit_module.TX_ADDR_7 ));
    LocalMux I__3703 (
            .O(N__17692),
            .I(\transmit_module.TX_ADDR_7 ));
    InMux I__3702 (
            .O(N__17683),
            .I(N__17680));
    LocalMux I__3701 (
            .O(N__17680),
            .I(N__17677));
    Span4Mux_h I__3700 (
            .O(N__17677),
            .I(N__17674));
    Odrv4 I__3699 (
            .O(N__17674),
            .I(\transmit_module.n197 ));
    InMux I__3698 (
            .O(N__17671),
            .I(\transmit_module.n3662 ));
    InMux I__3697 (
            .O(N__17668),
            .I(N__17665));
    LocalMux I__3696 (
            .O(N__17665),
            .I(N__17662));
    Span4Mux_h I__3695 (
            .O(N__17662),
            .I(N__17659));
    Odrv4 I__3694 (
            .O(N__17659),
            .I(\transmit_module.n196 ));
    InMux I__3693 (
            .O(N__17656),
            .I(bfn_15_18_0_));
    InMux I__3692 (
            .O(N__17653),
            .I(N__17650));
    LocalMux I__3691 (
            .O(N__17650),
            .I(N__17647));
    Odrv4 I__3690 (
            .O(N__17647),
            .I(\transmit_module.n195 ));
    InMux I__3689 (
            .O(N__17644),
            .I(\transmit_module.n3664 ));
    InMux I__3688 (
            .O(N__17641),
            .I(N__17638));
    LocalMux I__3687 (
            .O(N__17638),
            .I(\transmit_module.X_DELTA_PATTERN_7 ));
    InMux I__3686 (
            .O(N__17635),
            .I(N__17632));
    LocalMux I__3685 (
            .O(N__17632),
            .I(\transmit_module.X_DELTA_PATTERN_6 ));
    InMux I__3684 (
            .O(N__17629),
            .I(N__17626));
    LocalMux I__3683 (
            .O(N__17626),
            .I(N__17623));
    Odrv4 I__3682 (
            .O(N__17623),
            .I(\transmit_module.X_DELTA_PATTERN_14 ));
    InMux I__3681 (
            .O(N__17620),
            .I(N__17617));
    LocalMux I__3680 (
            .O(N__17617),
            .I(\transmit_module.X_DELTA_PATTERN_2 ));
    InMux I__3679 (
            .O(N__17614),
            .I(N__17611));
    LocalMux I__3678 (
            .O(N__17611),
            .I(\transmit_module.X_DELTA_PATTERN_1 ));
    InMux I__3677 (
            .O(N__17608),
            .I(N__17605));
    LocalMux I__3676 (
            .O(N__17605),
            .I(\transmit_module.X_DELTA_PATTERN_3 ));
    InMux I__3675 (
            .O(N__17602),
            .I(N__17599));
    LocalMux I__3674 (
            .O(N__17599),
            .I(\transmit_module.X_DELTA_PATTERN_15 ));
    InMux I__3673 (
            .O(N__17596),
            .I(N__17593));
    LocalMux I__3672 (
            .O(N__17593),
            .I(\transmit_module.X_DELTA_PATTERN_5 ));
    InMux I__3671 (
            .O(N__17590),
            .I(N__17587));
    LocalMux I__3670 (
            .O(N__17587),
            .I(\transmit_module.X_DELTA_PATTERN_4 ));
    CEMux I__3669 (
            .O(N__17584),
            .I(N__17579));
    CEMux I__3668 (
            .O(N__17583),
            .I(N__17575));
    CEMux I__3667 (
            .O(N__17582),
            .I(N__17572));
    LocalMux I__3666 (
            .O(N__17579),
            .I(N__17568));
    CEMux I__3665 (
            .O(N__17578),
            .I(N__17565));
    LocalMux I__3664 (
            .O(N__17575),
            .I(N__17562));
    LocalMux I__3663 (
            .O(N__17572),
            .I(N__17559));
    CEMux I__3662 (
            .O(N__17571),
            .I(N__17556));
    Span4Mux_v I__3661 (
            .O(N__17568),
            .I(N__17551));
    LocalMux I__3660 (
            .O(N__17565),
            .I(N__17551));
    Span4Mux_v I__3659 (
            .O(N__17562),
            .I(N__17548));
    Span4Mux_h I__3658 (
            .O(N__17559),
            .I(N__17541));
    LocalMux I__3657 (
            .O(N__17556),
            .I(N__17541));
    Span4Mux_h I__3656 (
            .O(N__17551),
            .I(N__17541));
    Odrv4 I__3655 (
            .O(N__17548),
            .I(\transmit_module.n2315 ));
    Odrv4 I__3654 (
            .O(N__17541),
            .I(\transmit_module.n2315 ));
    CascadeMux I__3653 (
            .O(N__17536),
            .I(N__17532));
    InMux I__3652 (
            .O(N__17535),
            .I(N__17529));
    InMux I__3651 (
            .O(N__17532),
            .I(N__17526));
    LocalMux I__3650 (
            .O(N__17529),
            .I(\transmit_module.X_DELTA_PATTERN_0 ));
    LocalMux I__3649 (
            .O(N__17526),
            .I(\transmit_module.X_DELTA_PATTERN_0 ));
    CascadeMux I__3648 (
            .O(N__17521),
            .I(N__17518));
    InMux I__3647 (
            .O(N__17518),
            .I(N__17515));
    LocalMux I__3646 (
            .O(N__17515),
            .I(N__17512));
    Span4Mux_h I__3645 (
            .O(N__17512),
            .I(N__17509));
    Odrv4 I__3644 (
            .O(N__17509),
            .I(\transmit_module.n204 ));
    InMux I__3643 (
            .O(N__17506),
            .I(\transmit_module.n3656 ));
    InMux I__3642 (
            .O(N__17503),
            .I(N__17499));
    InMux I__3641 (
            .O(N__17502),
            .I(N__17494));
    LocalMux I__3640 (
            .O(N__17499),
            .I(N__17491));
    InMux I__3639 (
            .O(N__17498),
            .I(N__17488));
    InMux I__3638 (
            .O(N__17497),
            .I(N__17485));
    LocalMux I__3637 (
            .O(N__17494),
            .I(\receive_module.rx_counter.X_8 ));
    Odrv12 I__3636 (
            .O(N__17491),
            .I(\receive_module.rx_counter.X_8 ));
    LocalMux I__3635 (
            .O(N__17488),
            .I(\receive_module.rx_counter.X_8 ));
    LocalMux I__3634 (
            .O(N__17485),
            .I(\receive_module.rx_counter.X_8 ));
    InMux I__3633 (
            .O(N__17476),
            .I(N__17472));
    InMux I__3632 (
            .O(N__17475),
            .I(N__17467));
    LocalMux I__3631 (
            .O(N__17472),
            .I(N__17464));
    InMux I__3630 (
            .O(N__17471),
            .I(N__17461));
    InMux I__3629 (
            .O(N__17470),
            .I(N__17458));
    LocalMux I__3628 (
            .O(N__17467),
            .I(\receive_module.rx_counter.X_9 ));
    Odrv4 I__3627 (
            .O(N__17464),
            .I(\receive_module.rx_counter.X_9 ));
    LocalMux I__3626 (
            .O(N__17461),
            .I(\receive_module.rx_counter.X_9 ));
    LocalMux I__3625 (
            .O(N__17458),
            .I(\receive_module.rx_counter.X_9 ));
    InMux I__3624 (
            .O(N__17449),
            .I(N__17446));
    LocalMux I__3623 (
            .O(N__17446),
            .I(\receive_module.rx_counter.n4219 ));
    CascadeMux I__3622 (
            .O(N__17443),
            .I(N__17438));
    InMux I__3621 (
            .O(N__17442),
            .I(N__17434));
    InMux I__3620 (
            .O(N__17441),
            .I(N__17431));
    InMux I__3619 (
            .O(N__17438),
            .I(N__17426));
    InMux I__3618 (
            .O(N__17437),
            .I(N__17426));
    LocalMux I__3617 (
            .O(N__17434),
            .I(\receive_module.rx_counter.X_7 ));
    LocalMux I__3616 (
            .O(N__17431),
            .I(\receive_module.rx_counter.X_7 ));
    LocalMux I__3615 (
            .O(N__17426),
            .I(\receive_module.rx_counter.X_7 ));
    CascadeMux I__3614 (
            .O(N__17419),
            .I(\receive_module.rx_counter.n4_adj_575_cascade_ ));
    InMux I__3613 (
            .O(N__17416),
            .I(N__17413));
    LocalMux I__3612 (
            .O(N__17413),
            .I(N__17409));
    InMux I__3611 (
            .O(N__17412),
            .I(N__17404));
    Span4Mux_h I__3610 (
            .O(N__17409),
            .I(N__17401));
    InMux I__3609 (
            .O(N__17408),
            .I(N__17398));
    InMux I__3608 (
            .O(N__17407),
            .I(N__17395));
    LocalMux I__3607 (
            .O(N__17404),
            .I(\receive_module.rx_counter.X_6 ));
    Odrv4 I__3606 (
            .O(N__17401),
            .I(\receive_module.rx_counter.X_6 ));
    LocalMux I__3605 (
            .O(N__17398),
            .I(\receive_module.rx_counter.X_6 ));
    LocalMux I__3604 (
            .O(N__17395),
            .I(\receive_module.rx_counter.X_6 ));
    InMux I__3603 (
            .O(N__17386),
            .I(N__17383));
    LocalMux I__3602 (
            .O(N__17383),
            .I(N__17380));
    Span4Mux_h I__3601 (
            .O(N__17380),
            .I(N__17377));
    Odrv4 I__3600 (
            .O(N__17377),
            .I(\receive_module.rx_counter.O_VISIBLE_N_86 ));
    InMux I__3599 (
            .O(N__17374),
            .I(N__17371));
    LocalMux I__3598 (
            .O(N__17371),
            .I(N__17367));
    InMux I__3597 (
            .O(N__17370),
            .I(N__17364));
    Odrv4 I__3596 (
            .O(N__17367),
            .I(\receive_module.rx_counter.n11 ));
    LocalMux I__3595 (
            .O(N__17364),
            .I(\receive_module.rx_counter.n11 ));
    IoInMux I__3594 (
            .O(N__17359),
            .I(N__17356));
    LocalMux I__3593 (
            .O(N__17356),
            .I(N__17353));
    Span4Mux_s1_v I__3592 (
            .O(N__17353),
            .I(N__17350));
    Span4Mux_v I__3591 (
            .O(N__17350),
            .I(N__17347));
    Span4Mux_v I__3590 (
            .O(N__17347),
            .I(N__17344));
    Span4Mux_h I__3589 (
            .O(N__17344),
            .I(N__17340));
    InMux I__3588 (
            .O(N__17343),
            .I(N__17337));
    Odrv4 I__3587 (
            .O(N__17340),
            .I(LED_c));
    LocalMux I__3586 (
            .O(N__17337),
            .I(LED_c));
    CEMux I__3585 (
            .O(N__17332),
            .I(N__17328));
    CEMux I__3584 (
            .O(N__17331),
            .I(N__17325));
    LocalMux I__3583 (
            .O(N__17328),
            .I(\receive_module.rx_counter.n4222 ));
    LocalMux I__3582 (
            .O(N__17325),
            .I(\receive_module.rx_counter.n4222 ));
    InMux I__3581 (
            .O(N__17320),
            .I(N__17317));
    LocalMux I__3580 (
            .O(N__17317),
            .I(N__17314));
    Span4Mux_v I__3579 (
            .O(N__17314),
            .I(N__17311));
    Sp12to4 I__3578 (
            .O(N__17311),
            .I(N__17308));
    Span12Mux_h I__3577 (
            .O(N__17308),
            .I(N__17305));
    Odrv12 I__3576 (
            .O(N__17305),
            .I(\line_buffer.n623 ));
    InMux I__3575 (
            .O(N__17302),
            .I(N__17299));
    LocalMux I__3574 (
            .O(N__17299),
            .I(N__17296));
    Span4Mux_v I__3573 (
            .O(N__17296),
            .I(N__17293));
    Span4Mux_v I__3572 (
            .O(N__17293),
            .I(N__17290));
    Span4Mux_v I__3571 (
            .O(N__17290),
            .I(N__17287));
    Sp12to4 I__3570 (
            .O(N__17287),
            .I(N__17284));
    Odrv12 I__3569 (
            .O(N__17284),
            .I(\line_buffer.n615 ));
    InMux I__3568 (
            .O(N__17281),
            .I(N__17278));
    LocalMux I__3567 (
            .O(N__17278),
            .I(N__17275));
    Odrv4 I__3566 (
            .O(N__17275),
            .I(\line_buffer.n4071 ));
    InMux I__3565 (
            .O(N__17272),
            .I(N__17269));
    LocalMux I__3564 (
            .O(N__17269),
            .I(N__17266));
    Span12Mux_h I__3563 (
            .O(N__17266),
            .I(N__17263));
    Odrv12 I__3562 (
            .O(N__17263),
            .I(\line_buffer.n646 ));
    CascadeMux I__3561 (
            .O(N__17260),
            .I(N__17257));
    InMux I__3560 (
            .O(N__17257),
            .I(N__17254));
    LocalMux I__3559 (
            .O(N__17254),
            .I(N__17251));
    Span4Mux_v I__3558 (
            .O(N__17251),
            .I(N__17248));
    Span4Mux_h I__3557 (
            .O(N__17248),
            .I(N__17245));
    Span4Mux_h I__3556 (
            .O(N__17245),
            .I(N__17242));
    Odrv4 I__3555 (
            .O(N__17242),
            .I(\line_buffer.n654 ));
    InMux I__3554 (
            .O(N__17239),
            .I(N__17236));
    LocalMux I__3553 (
            .O(N__17236),
            .I(N__17233));
    Span4Mux_v I__3552 (
            .O(N__17233),
            .I(N__17230));
    Span4Mux_h I__3551 (
            .O(N__17230),
            .I(N__17227));
    Sp12to4 I__3550 (
            .O(N__17227),
            .I(N__17224));
    Span12Mux_v I__3549 (
            .O(N__17224),
            .I(N__17221));
    Odrv12 I__3548 (
            .O(N__17221),
            .I(\line_buffer.n549 ));
    CascadeMux I__3547 (
            .O(N__17218),
            .I(\line_buffer.n4176_cascade_ ));
    InMux I__3546 (
            .O(N__17215),
            .I(N__17212));
    LocalMux I__3545 (
            .O(N__17212),
            .I(N__17209));
    Span4Mux_v I__3544 (
            .O(N__17209),
            .I(N__17206));
    Span4Mux_v I__3543 (
            .O(N__17206),
            .I(N__17203));
    Sp12to4 I__3542 (
            .O(N__17203),
            .I(N__17200));
    Odrv12 I__3541 (
            .O(N__17200),
            .I(\line_buffer.n557 ));
    InMux I__3540 (
            .O(N__17197),
            .I(N__17194));
    LocalMux I__3539 (
            .O(N__17194),
            .I(\transmit_module.X_DELTA_PATTERN_8 ));
    InMux I__3538 (
            .O(N__17191),
            .I(\receive_module.rx_counter.n3706 ));
    InMux I__3537 (
            .O(N__17188),
            .I(N__17184));
    InMux I__3536 (
            .O(N__17187),
            .I(N__17181));
    LocalMux I__3535 (
            .O(N__17184),
            .I(\receive_module.rx_counter.FRAME_COUNTER_2 ));
    LocalMux I__3534 (
            .O(N__17181),
            .I(\receive_module.rx_counter.FRAME_COUNTER_2 ));
    InMux I__3533 (
            .O(N__17176),
            .I(\receive_module.rx_counter.n3707 ));
    InMux I__3532 (
            .O(N__17173),
            .I(N__17169));
    InMux I__3531 (
            .O(N__17172),
            .I(N__17166));
    LocalMux I__3530 (
            .O(N__17169),
            .I(\receive_module.rx_counter.FRAME_COUNTER_3 ));
    LocalMux I__3529 (
            .O(N__17166),
            .I(\receive_module.rx_counter.FRAME_COUNTER_3 ));
    InMux I__3528 (
            .O(N__17161),
            .I(\receive_module.rx_counter.n3708 ));
    InMux I__3527 (
            .O(N__17158),
            .I(N__17154));
    InMux I__3526 (
            .O(N__17157),
            .I(N__17151));
    LocalMux I__3525 (
            .O(N__17154),
            .I(\receive_module.rx_counter.FRAME_COUNTER_4 ));
    LocalMux I__3524 (
            .O(N__17151),
            .I(\receive_module.rx_counter.FRAME_COUNTER_4 ));
    InMux I__3523 (
            .O(N__17146),
            .I(\receive_module.rx_counter.n3709 ));
    InMux I__3522 (
            .O(N__17143),
            .I(\receive_module.rx_counter.n3710 ));
    InMux I__3521 (
            .O(N__17140),
            .I(N__17136));
    InMux I__3520 (
            .O(N__17139),
            .I(N__17133));
    LocalMux I__3519 (
            .O(N__17136),
            .I(\receive_module.rx_counter.FRAME_COUNTER_5 ));
    LocalMux I__3518 (
            .O(N__17133),
            .I(\receive_module.rx_counter.FRAME_COUNTER_5 ));
    SRMux I__3517 (
            .O(N__17128),
            .I(N__17125));
    LocalMux I__3516 (
            .O(N__17125),
            .I(N__17122));
    Odrv12 I__3515 (
            .O(N__17122),
            .I(\receive_module.rx_counter.n2605 ));
    InMux I__3514 (
            .O(N__17119),
            .I(N__17113));
    InMux I__3513 (
            .O(N__17118),
            .I(N__17113));
    LocalMux I__3512 (
            .O(N__17113),
            .I(\receive_module.rx_counter.old_VS ));
    InMux I__3511 (
            .O(N__17110),
            .I(N__17107));
    LocalMux I__3510 (
            .O(N__17107),
            .I(N__17103));
    InMux I__3509 (
            .O(N__17106),
            .I(N__17100));
    Span4Mux_h I__3508 (
            .O(N__17103),
            .I(N__17094));
    LocalMux I__3507 (
            .O(N__17100),
            .I(N__17091));
    InMux I__3506 (
            .O(N__17099),
            .I(N__17084));
    InMux I__3505 (
            .O(N__17098),
            .I(N__17084));
    InMux I__3504 (
            .O(N__17097),
            .I(N__17084));
    Sp12to4 I__3503 (
            .O(N__17094),
            .I(N__17077));
    Span12Mux_h I__3502 (
            .O(N__17091),
            .I(N__17077));
    LocalMux I__3501 (
            .O(N__17084),
            .I(N__17077));
    Odrv12 I__3500 (
            .O(N__17077),
            .I(TVP_VSYNC_c));
    CascadeMux I__3499 (
            .O(N__17074),
            .I(N__17068));
    InMux I__3498 (
            .O(N__17073),
            .I(N__17065));
    InMux I__3497 (
            .O(N__17072),
            .I(N__17062));
    InMux I__3496 (
            .O(N__17071),
            .I(N__17057));
    InMux I__3495 (
            .O(N__17068),
            .I(N__17057));
    LocalMux I__3494 (
            .O(N__17065),
            .I(\receive_module.rx_counter.X_5 ));
    LocalMux I__3493 (
            .O(N__17062),
            .I(\receive_module.rx_counter.X_5 ));
    LocalMux I__3492 (
            .O(N__17057),
            .I(\receive_module.rx_counter.X_5 ));
    InMux I__3491 (
            .O(N__17050),
            .I(N__17044));
    InMux I__3490 (
            .O(N__17049),
            .I(N__17041));
    InMux I__3489 (
            .O(N__17048),
            .I(N__17036));
    InMux I__3488 (
            .O(N__17047),
            .I(N__17036));
    LocalMux I__3487 (
            .O(N__17044),
            .I(\receive_module.rx_counter.X_4 ));
    LocalMux I__3486 (
            .O(N__17041),
            .I(\receive_module.rx_counter.X_4 ));
    LocalMux I__3485 (
            .O(N__17036),
            .I(\receive_module.rx_counter.X_4 ));
    InMux I__3484 (
            .O(N__17029),
            .I(N__17023));
    InMux I__3483 (
            .O(N__17028),
            .I(N__17020));
    InMux I__3482 (
            .O(N__17027),
            .I(N__17015));
    InMux I__3481 (
            .O(N__17026),
            .I(N__17015));
    LocalMux I__3480 (
            .O(N__17023),
            .I(\receive_module.rx_counter.X_3 ));
    LocalMux I__3479 (
            .O(N__17020),
            .I(\receive_module.rx_counter.X_3 ));
    LocalMux I__3478 (
            .O(N__17015),
            .I(\receive_module.rx_counter.X_3 ));
    CascadeMux I__3477 (
            .O(N__17008),
            .I(N__17005));
    InMux I__3476 (
            .O(N__17005),
            .I(N__17001));
    CascadeMux I__3475 (
            .O(N__17004),
            .I(N__16998));
    LocalMux I__3474 (
            .O(N__17001),
            .I(N__16995));
    InMux I__3473 (
            .O(N__16998),
            .I(N__16992));
    Odrv4 I__3472 (
            .O(N__16995),
            .I(\transmit_module.n180 ));
    LocalMux I__3471 (
            .O(N__16992),
            .I(\transmit_module.n180 ));
    InMux I__3470 (
            .O(N__16987),
            .I(N__16983));
    InMux I__3469 (
            .O(N__16986),
            .I(N__16980));
    LocalMux I__3468 (
            .O(N__16983),
            .I(\transmit_module.n211 ));
    LocalMux I__3467 (
            .O(N__16980),
            .I(\transmit_module.n211 ));
    CascadeMux I__3466 (
            .O(N__16975),
            .I(N__16971));
    CascadeMux I__3465 (
            .O(N__16974),
            .I(N__16968));
    CascadeBuf I__3464 (
            .O(N__16971),
            .I(N__16965));
    CascadeBuf I__3463 (
            .O(N__16968),
            .I(N__16962));
    CascadeMux I__3462 (
            .O(N__16965),
            .I(N__16959));
    CascadeMux I__3461 (
            .O(N__16962),
            .I(N__16956));
    CascadeBuf I__3460 (
            .O(N__16959),
            .I(N__16953));
    CascadeBuf I__3459 (
            .O(N__16956),
            .I(N__16950));
    CascadeMux I__3458 (
            .O(N__16953),
            .I(N__16947));
    CascadeMux I__3457 (
            .O(N__16950),
            .I(N__16944));
    CascadeBuf I__3456 (
            .O(N__16947),
            .I(N__16941));
    CascadeBuf I__3455 (
            .O(N__16944),
            .I(N__16938));
    CascadeMux I__3454 (
            .O(N__16941),
            .I(N__16935));
    CascadeMux I__3453 (
            .O(N__16938),
            .I(N__16932));
    CascadeBuf I__3452 (
            .O(N__16935),
            .I(N__16929));
    CascadeBuf I__3451 (
            .O(N__16932),
            .I(N__16926));
    CascadeMux I__3450 (
            .O(N__16929),
            .I(N__16923));
    CascadeMux I__3449 (
            .O(N__16926),
            .I(N__16920));
    CascadeBuf I__3448 (
            .O(N__16923),
            .I(N__16917));
    CascadeBuf I__3447 (
            .O(N__16920),
            .I(N__16914));
    CascadeMux I__3446 (
            .O(N__16917),
            .I(N__16911));
    CascadeMux I__3445 (
            .O(N__16914),
            .I(N__16908));
    CascadeBuf I__3444 (
            .O(N__16911),
            .I(N__16905));
    CascadeBuf I__3443 (
            .O(N__16908),
            .I(N__16902));
    CascadeMux I__3442 (
            .O(N__16905),
            .I(N__16899));
    CascadeMux I__3441 (
            .O(N__16902),
            .I(N__16896));
    CascadeBuf I__3440 (
            .O(N__16899),
            .I(N__16893));
    CascadeBuf I__3439 (
            .O(N__16896),
            .I(N__16890));
    CascadeMux I__3438 (
            .O(N__16893),
            .I(N__16887));
    CascadeMux I__3437 (
            .O(N__16890),
            .I(N__16884));
    CascadeBuf I__3436 (
            .O(N__16887),
            .I(N__16881));
    CascadeBuf I__3435 (
            .O(N__16884),
            .I(N__16878));
    CascadeMux I__3434 (
            .O(N__16881),
            .I(N__16875));
    CascadeMux I__3433 (
            .O(N__16878),
            .I(N__16872));
    CascadeBuf I__3432 (
            .O(N__16875),
            .I(N__16869));
    CascadeBuf I__3431 (
            .O(N__16872),
            .I(N__16866));
    CascadeMux I__3430 (
            .O(N__16869),
            .I(N__16863));
    CascadeMux I__3429 (
            .O(N__16866),
            .I(N__16860));
    CascadeBuf I__3428 (
            .O(N__16863),
            .I(N__16857));
    CascadeBuf I__3427 (
            .O(N__16860),
            .I(N__16854));
    CascadeMux I__3426 (
            .O(N__16857),
            .I(N__16851));
    CascadeMux I__3425 (
            .O(N__16854),
            .I(N__16848));
    CascadeBuf I__3424 (
            .O(N__16851),
            .I(N__16845));
    CascadeBuf I__3423 (
            .O(N__16848),
            .I(N__16842));
    CascadeMux I__3422 (
            .O(N__16845),
            .I(N__16839));
    CascadeMux I__3421 (
            .O(N__16842),
            .I(N__16836));
    CascadeBuf I__3420 (
            .O(N__16839),
            .I(N__16833));
    CascadeBuf I__3419 (
            .O(N__16836),
            .I(N__16830));
    CascadeMux I__3418 (
            .O(N__16833),
            .I(N__16827));
    CascadeMux I__3417 (
            .O(N__16830),
            .I(N__16824));
    CascadeBuf I__3416 (
            .O(N__16827),
            .I(N__16821));
    CascadeBuf I__3415 (
            .O(N__16824),
            .I(N__16818));
    CascadeMux I__3414 (
            .O(N__16821),
            .I(N__16815));
    CascadeMux I__3413 (
            .O(N__16818),
            .I(N__16812));
    CascadeBuf I__3412 (
            .O(N__16815),
            .I(N__16809));
    CascadeBuf I__3411 (
            .O(N__16812),
            .I(N__16806));
    CascadeMux I__3410 (
            .O(N__16809),
            .I(N__16803));
    CascadeMux I__3409 (
            .O(N__16806),
            .I(N__16800));
    CascadeBuf I__3408 (
            .O(N__16803),
            .I(N__16797));
    CascadeBuf I__3407 (
            .O(N__16800),
            .I(N__16794));
    CascadeMux I__3406 (
            .O(N__16797),
            .I(N__16791));
    CascadeMux I__3405 (
            .O(N__16794),
            .I(N__16788));
    InMux I__3404 (
            .O(N__16791),
            .I(N__16785));
    InMux I__3403 (
            .O(N__16788),
            .I(N__16782));
    LocalMux I__3402 (
            .O(N__16785),
            .I(N__16779));
    LocalMux I__3401 (
            .O(N__16782),
            .I(N__16776));
    Span12Mux_s11_h I__3400 (
            .O(N__16779),
            .I(N__16773));
    Span12Mux_s8_h I__3399 (
            .O(N__16776),
            .I(N__16770));
    Span12Mux_v I__3398 (
            .O(N__16773),
            .I(N__16765));
    Span12Mux_v I__3397 (
            .O(N__16770),
            .I(N__16765));
    Odrv12 I__3396 (
            .O(N__16765),
            .I(n20));
    InMux I__3395 (
            .O(N__16762),
            .I(N__16757));
    InMux I__3394 (
            .O(N__16761),
            .I(N__16752));
    InMux I__3393 (
            .O(N__16760),
            .I(N__16749));
    LocalMux I__3392 (
            .O(N__16757),
            .I(N__16746));
    InMux I__3391 (
            .O(N__16756),
            .I(N__16743));
    InMux I__3390 (
            .O(N__16755),
            .I(N__16740));
    LocalMux I__3389 (
            .O(N__16752),
            .I(\transmit_module.old_VGA_HS ));
    LocalMux I__3388 (
            .O(N__16749),
            .I(\transmit_module.old_VGA_HS ));
    Odrv4 I__3387 (
            .O(N__16746),
            .I(\transmit_module.old_VGA_HS ));
    LocalMux I__3386 (
            .O(N__16743),
            .I(\transmit_module.old_VGA_HS ));
    LocalMux I__3385 (
            .O(N__16740),
            .I(\transmit_module.old_VGA_HS ));
    IoInMux I__3384 (
            .O(N__16729),
            .I(N__16726));
    LocalMux I__3383 (
            .O(N__16726),
            .I(N__16723));
    Span4Mux_s0_h I__3382 (
            .O(N__16723),
            .I(N__16720));
    Span4Mux_h I__3381 (
            .O(N__16720),
            .I(N__16714));
    InMux I__3380 (
            .O(N__16719),
            .I(N__16709));
    InMux I__3379 (
            .O(N__16718),
            .I(N__16706));
    InMux I__3378 (
            .O(N__16717),
            .I(N__16702));
    Span4Mux_h I__3377 (
            .O(N__16714),
            .I(N__16699));
    InMux I__3376 (
            .O(N__16713),
            .I(N__16694));
    InMux I__3375 (
            .O(N__16712),
            .I(N__16694));
    LocalMux I__3374 (
            .O(N__16709),
            .I(N__16689));
    LocalMux I__3373 (
            .O(N__16706),
            .I(N__16689));
    InMux I__3372 (
            .O(N__16705),
            .I(N__16686));
    LocalMux I__3371 (
            .O(N__16702),
            .I(N__16683));
    Span4Mux_h I__3370 (
            .O(N__16699),
            .I(N__16678));
    LocalMux I__3369 (
            .O(N__16694),
            .I(N__16678));
    Span12Mux_v I__3368 (
            .O(N__16689),
            .I(N__16675));
    LocalMux I__3367 (
            .O(N__16686),
            .I(N__16668));
    Span4Mux_v I__3366 (
            .O(N__16683),
            .I(N__16668));
    Span4Mux_v I__3365 (
            .O(N__16678),
            .I(N__16668));
    Odrv12 I__3364 (
            .O(N__16675),
            .I(ADV_HSYNC_c));
    Odrv4 I__3363 (
            .O(N__16668),
            .I(ADV_HSYNC_c));
    CascadeMux I__3362 (
            .O(N__16663),
            .I(N__16660));
    InMux I__3361 (
            .O(N__16660),
            .I(N__16657));
    LocalMux I__3360 (
            .O(N__16657),
            .I(\transmit_module.n181 ));
    InMux I__3359 (
            .O(N__16654),
            .I(N__16650));
    InMux I__3358 (
            .O(N__16653),
            .I(N__16647));
    LocalMux I__3357 (
            .O(N__16650),
            .I(\transmit_module.n212 ));
    LocalMux I__3356 (
            .O(N__16647),
            .I(\transmit_module.n212 ));
    CascadeMux I__3355 (
            .O(N__16642),
            .I(\transmit_module.n181_cascade_ ));
    CascadeMux I__3354 (
            .O(N__16639),
            .I(N__16635));
    CascadeMux I__3353 (
            .O(N__16638),
            .I(N__16632));
    CascadeBuf I__3352 (
            .O(N__16635),
            .I(N__16629));
    CascadeBuf I__3351 (
            .O(N__16632),
            .I(N__16626));
    CascadeMux I__3350 (
            .O(N__16629),
            .I(N__16623));
    CascadeMux I__3349 (
            .O(N__16626),
            .I(N__16620));
    CascadeBuf I__3348 (
            .O(N__16623),
            .I(N__16617));
    CascadeBuf I__3347 (
            .O(N__16620),
            .I(N__16614));
    CascadeMux I__3346 (
            .O(N__16617),
            .I(N__16611));
    CascadeMux I__3345 (
            .O(N__16614),
            .I(N__16608));
    CascadeBuf I__3344 (
            .O(N__16611),
            .I(N__16605));
    CascadeBuf I__3343 (
            .O(N__16608),
            .I(N__16602));
    CascadeMux I__3342 (
            .O(N__16605),
            .I(N__16599));
    CascadeMux I__3341 (
            .O(N__16602),
            .I(N__16596));
    CascadeBuf I__3340 (
            .O(N__16599),
            .I(N__16593));
    CascadeBuf I__3339 (
            .O(N__16596),
            .I(N__16590));
    CascadeMux I__3338 (
            .O(N__16593),
            .I(N__16587));
    CascadeMux I__3337 (
            .O(N__16590),
            .I(N__16584));
    CascadeBuf I__3336 (
            .O(N__16587),
            .I(N__16581));
    CascadeBuf I__3335 (
            .O(N__16584),
            .I(N__16578));
    CascadeMux I__3334 (
            .O(N__16581),
            .I(N__16575));
    CascadeMux I__3333 (
            .O(N__16578),
            .I(N__16572));
    CascadeBuf I__3332 (
            .O(N__16575),
            .I(N__16569));
    CascadeBuf I__3331 (
            .O(N__16572),
            .I(N__16566));
    CascadeMux I__3330 (
            .O(N__16569),
            .I(N__16563));
    CascadeMux I__3329 (
            .O(N__16566),
            .I(N__16560));
    CascadeBuf I__3328 (
            .O(N__16563),
            .I(N__16557));
    CascadeBuf I__3327 (
            .O(N__16560),
            .I(N__16554));
    CascadeMux I__3326 (
            .O(N__16557),
            .I(N__16551));
    CascadeMux I__3325 (
            .O(N__16554),
            .I(N__16548));
    CascadeBuf I__3324 (
            .O(N__16551),
            .I(N__16545));
    CascadeBuf I__3323 (
            .O(N__16548),
            .I(N__16542));
    CascadeMux I__3322 (
            .O(N__16545),
            .I(N__16539));
    CascadeMux I__3321 (
            .O(N__16542),
            .I(N__16536));
    CascadeBuf I__3320 (
            .O(N__16539),
            .I(N__16533));
    CascadeBuf I__3319 (
            .O(N__16536),
            .I(N__16530));
    CascadeMux I__3318 (
            .O(N__16533),
            .I(N__16527));
    CascadeMux I__3317 (
            .O(N__16530),
            .I(N__16524));
    CascadeBuf I__3316 (
            .O(N__16527),
            .I(N__16521));
    CascadeBuf I__3315 (
            .O(N__16524),
            .I(N__16518));
    CascadeMux I__3314 (
            .O(N__16521),
            .I(N__16515));
    CascadeMux I__3313 (
            .O(N__16518),
            .I(N__16512));
    CascadeBuf I__3312 (
            .O(N__16515),
            .I(N__16509));
    CascadeBuf I__3311 (
            .O(N__16512),
            .I(N__16506));
    CascadeMux I__3310 (
            .O(N__16509),
            .I(N__16503));
    CascadeMux I__3309 (
            .O(N__16506),
            .I(N__16500));
    CascadeBuf I__3308 (
            .O(N__16503),
            .I(N__16497));
    CascadeBuf I__3307 (
            .O(N__16500),
            .I(N__16494));
    CascadeMux I__3306 (
            .O(N__16497),
            .I(N__16491));
    CascadeMux I__3305 (
            .O(N__16494),
            .I(N__16488));
    CascadeBuf I__3304 (
            .O(N__16491),
            .I(N__16485));
    CascadeBuf I__3303 (
            .O(N__16488),
            .I(N__16482));
    CascadeMux I__3302 (
            .O(N__16485),
            .I(N__16479));
    CascadeMux I__3301 (
            .O(N__16482),
            .I(N__16476));
    CascadeBuf I__3300 (
            .O(N__16479),
            .I(N__16473));
    CascadeBuf I__3299 (
            .O(N__16476),
            .I(N__16470));
    CascadeMux I__3298 (
            .O(N__16473),
            .I(N__16467));
    CascadeMux I__3297 (
            .O(N__16470),
            .I(N__16464));
    CascadeBuf I__3296 (
            .O(N__16467),
            .I(N__16461));
    CascadeBuf I__3295 (
            .O(N__16464),
            .I(N__16458));
    CascadeMux I__3294 (
            .O(N__16461),
            .I(N__16455));
    CascadeMux I__3293 (
            .O(N__16458),
            .I(N__16452));
    InMux I__3292 (
            .O(N__16455),
            .I(N__16449));
    InMux I__3291 (
            .O(N__16452),
            .I(N__16446));
    LocalMux I__3290 (
            .O(N__16449),
            .I(N__16443));
    LocalMux I__3289 (
            .O(N__16446),
            .I(N__16440));
    Span12Mux_h I__3288 (
            .O(N__16443),
            .I(N__16435));
    Span12Mux_h I__3287 (
            .O(N__16440),
            .I(N__16435));
    Span12Mux_v I__3286 (
            .O(N__16435),
            .I(N__16432));
    Odrv12 I__3285 (
            .O(N__16432),
            .I(n21));
    InMux I__3284 (
            .O(N__16429),
            .I(N__16426));
    LocalMux I__3283 (
            .O(N__16426),
            .I(N__16423));
    Odrv4 I__3282 (
            .O(N__16423),
            .I(\transmit_module.ADDR_Y_COMPONENT_7 ));
    InMux I__3281 (
            .O(N__16420),
            .I(N__16417));
    LocalMux I__3280 (
            .O(N__16417),
            .I(\transmit_module.ADDR_Y_COMPONENT_6 ));
    InMux I__3279 (
            .O(N__16414),
            .I(N__16410));
    InMux I__3278 (
            .O(N__16413),
            .I(N__16407));
    LocalMux I__3277 (
            .O(N__16410),
            .I(N__16404));
    LocalMux I__3276 (
            .O(N__16407),
            .I(N__16401));
    Span4Mux_v I__3275 (
            .O(N__16404),
            .I(N__16398));
    Odrv12 I__3274 (
            .O(N__16401),
            .I(\transmit_module.n182 ));
    Odrv4 I__3273 (
            .O(N__16398),
            .I(\transmit_module.n182 ));
    InMux I__3272 (
            .O(N__16393),
            .I(N__16389));
    InMux I__3271 (
            .O(N__16392),
            .I(N__16386));
    LocalMux I__3270 (
            .O(N__16389),
            .I(\receive_module.rx_counter.FRAME_COUNTER_0 ));
    LocalMux I__3269 (
            .O(N__16386),
            .I(\receive_module.rx_counter.FRAME_COUNTER_0 ));
    InMux I__3268 (
            .O(N__16381),
            .I(bfn_15_8_0_));
    InMux I__3267 (
            .O(N__16378),
            .I(N__16374));
    InMux I__3266 (
            .O(N__16377),
            .I(N__16371));
    LocalMux I__3265 (
            .O(N__16374),
            .I(\receive_module.rx_counter.FRAME_COUNTER_1 ));
    LocalMux I__3264 (
            .O(N__16371),
            .I(\receive_module.rx_counter.FRAME_COUNTER_1 ));
    InMux I__3263 (
            .O(N__16366),
            .I(N__16363));
    LocalMux I__3262 (
            .O(N__16363),
            .I(\transmit_module.ADDR_Y_COMPONENT_2 ));
    InMux I__3261 (
            .O(N__16360),
            .I(N__16357));
    LocalMux I__3260 (
            .O(N__16357),
            .I(N__16354));
    Span4Mux_h I__3259 (
            .O(N__16354),
            .I(N__16351));
    Odrv4 I__3258 (
            .O(N__16351),
            .I(\transmit_module.n219 ));
    CascadeMux I__3257 (
            .O(N__16348),
            .I(\transmit_module.n179_cascade_ ));
    InMux I__3256 (
            .O(N__16345),
            .I(N__16342));
    LocalMux I__3255 (
            .O(N__16342),
            .I(N__16338));
    InMux I__3254 (
            .O(N__16341),
            .I(N__16335));
    Span12Mux_s6_v I__3253 (
            .O(N__16338),
            .I(N__16332));
    LocalMux I__3252 (
            .O(N__16335),
            .I(\transmit_module.n213 ));
    Odrv12 I__3251 (
            .O(N__16332),
            .I(\transmit_module.n213 ));
    InMux I__3250 (
            .O(N__16327),
            .I(N__16324));
    LocalMux I__3249 (
            .O(N__16324),
            .I(\transmit_module.n179 ));
    InMux I__3248 (
            .O(N__16321),
            .I(N__16317));
    InMux I__3247 (
            .O(N__16320),
            .I(N__16314));
    LocalMux I__3246 (
            .O(N__16317),
            .I(\transmit_module.n210 ));
    LocalMux I__3245 (
            .O(N__16314),
            .I(\transmit_module.n210 ));
    CascadeMux I__3244 (
            .O(N__16309),
            .I(N__16305));
    CascadeMux I__3243 (
            .O(N__16308),
            .I(N__16302));
    CascadeBuf I__3242 (
            .O(N__16305),
            .I(N__16299));
    CascadeBuf I__3241 (
            .O(N__16302),
            .I(N__16296));
    CascadeMux I__3240 (
            .O(N__16299),
            .I(N__16293));
    CascadeMux I__3239 (
            .O(N__16296),
            .I(N__16290));
    CascadeBuf I__3238 (
            .O(N__16293),
            .I(N__16287));
    CascadeBuf I__3237 (
            .O(N__16290),
            .I(N__16284));
    CascadeMux I__3236 (
            .O(N__16287),
            .I(N__16281));
    CascadeMux I__3235 (
            .O(N__16284),
            .I(N__16278));
    CascadeBuf I__3234 (
            .O(N__16281),
            .I(N__16275));
    CascadeBuf I__3233 (
            .O(N__16278),
            .I(N__16272));
    CascadeMux I__3232 (
            .O(N__16275),
            .I(N__16269));
    CascadeMux I__3231 (
            .O(N__16272),
            .I(N__16266));
    CascadeBuf I__3230 (
            .O(N__16269),
            .I(N__16263));
    CascadeBuf I__3229 (
            .O(N__16266),
            .I(N__16260));
    CascadeMux I__3228 (
            .O(N__16263),
            .I(N__16257));
    CascadeMux I__3227 (
            .O(N__16260),
            .I(N__16254));
    CascadeBuf I__3226 (
            .O(N__16257),
            .I(N__16251));
    CascadeBuf I__3225 (
            .O(N__16254),
            .I(N__16248));
    CascadeMux I__3224 (
            .O(N__16251),
            .I(N__16245));
    CascadeMux I__3223 (
            .O(N__16248),
            .I(N__16242));
    CascadeBuf I__3222 (
            .O(N__16245),
            .I(N__16239));
    CascadeBuf I__3221 (
            .O(N__16242),
            .I(N__16236));
    CascadeMux I__3220 (
            .O(N__16239),
            .I(N__16233));
    CascadeMux I__3219 (
            .O(N__16236),
            .I(N__16230));
    CascadeBuf I__3218 (
            .O(N__16233),
            .I(N__16227));
    CascadeBuf I__3217 (
            .O(N__16230),
            .I(N__16224));
    CascadeMux I__3216 (
            .O(N__16227),
            .I(N__16221));
    CascadeMux I__3215 (
            .O(N__16224),
            .I(N__16218));
    CascadeBuf I__3214 (
            .O(N__16221),
            .I(N__16215));
    CascadeBuf I__3213 (
            .O(N__16218),
            .I(N__16212));
    CascadeMux I__3212 (
            .O(N__16215),
            .I(N__16209));
    CascadeMux I__3211 (
            .O(N__16212),
            .I(N__16206));
    CascadeBuf I__3210 (
            .O(N__16209),
            .I(N__16203));
    CascadeBuf I__3209 (
            .O(N__16206),
            .I(N__16200));
    CascadeMux I__3208 (
            .O(N__16203),
            .I(N__16197));
    CascadeMux I__3207 (
            .O(N__16200),
            .I(N__16194));
    CascadeBuf I__3206 (
            .O(N__16197),
            .I(N__16191));
    CascadeBuf I__3205 (
            .O(N__16194),
            .I(N__16188));
    CascadeMux I__3204 (
            .O(N__16191),
            .I(N__16185));
    CascadeMux I__3203 (
            .O(N__16188),
            .I(N__16182));
    CascadeBuf I__3202 (
            .O(N__16185),
            .I(N__16179));
    CascadeBuf I__3201 (
            .O(N__16182),
            .I(N__16176));
    CascadeMux I__3200 (
            .O(N__16179),
            .I(N__16173));
    CascadeMux I__3199 (
            .O(N__16176),
            .I(N__16170));
    CascadeBuf I__3198 (
            .O(N__16173),
            .I(N__16167));
    CascadeBuf I__3197 (
            .O(N__16170),
            .I(N__16164));
    CascadeMux I__3196 (
            .O(N__16167),
            .I(N__16161));
    CascadeMux I__3195 (
            .O(N__16164),
            .I(N__16158));
    CascadeBuf I__3194 (
            .O(N__16161),
            .I(N__16155));
    CascadeBuf I__3193 (
            .O(N__16158),
            .I(N__16152));
    CascadeMux I__3192 (
            .O(N__16155),
            .I(N__16149));
    CascadeMux I__3191 (
            .O(N__16152),
            .I(N__16146));
    CascadeBuf I__3190 (
            .O(N__16149),
            .I(N__16143));
    CascadeBuf I__3189 (
            .O(N__16146),
            .I(N__16140));
    CascadeMux I__3188 (
            .O(N__16143),
            .I(N__16137));
    CascadeMux I__3187 (
            .O(N__16140),
            .I(N__16134));
    CascadeBuf I__3186 (
            .O(N__16137),
            .I(N__16131));
    CascadeBuf I__3185 (
            .O(N__16134),
            .I(N__16128));
    CascadeMux I__3184 (
            .O(N__16131),
            .I(N__16125));
    CascadeMux I__3183 (
            .O(N__16128),
            .I(N__16122));
    InMux I__3182 (
            .O(N__16125),
            .I(N__16119));
    InMux I__3181 (
            .O(N__16122),
            .I(N__16116));
    LocalMux I__3180 (
            .O(N__16119),
            .I(N__16113));
    LocalMux I__3179 (
            .O(N__16116),
            .I(N__16110));
    Span4Mux_h I__3178 (
            .O(N__16113),
            .I(N__16107));
    Span4Mux_h I__3177 (
            .O(N__16110),
            .I(N__16104));
    Sp12to4 I__3176 (
            .O(N__16107),
            .I(N__16101));
    Sp12to4 I__3175 (
            .O(N__16104),
            .I(N__16098));
    Span12Mux_v I__3174 (
            .O(N__16101),
            .I(N__16093));
    Span12Mux_v I__3173 (
            .O(N__16098),
            .I(N__16093));
    Odrv12 I__3172 (
            .O(N__16093),
            .I(n19));
    InMux I__3171 (
            .O(N__16090),
            .I(N__16087));
    LocalMux I__3170 (
            .O(N__16087),
            .I(\transmit_module.X_DELTA_PATTERN_13 ));
    InMux I__3169 (
            .O(N__16084),
            .I(N__16081));
    LocalMux I__3168 (
            .O(N__16081),
            .I(\transmit_module.X_DELTA_PATTERN_9 ));
    InMux I__3167 (
            .O(N__16078),
            .I(N__16075));
    LocalMux I__3166 (
            .O(N__16075),
            .I(\transmit_module.X_DELTA_PATTERN_12 ));
    InMux I__3165 (
            .O(N__16072),
            .I(N__16069));
    LocalMux I__3164 (
            .O(N__16069),
            .I(\transmit_module.X_DELTA_PATTERN_11 ));
    InMux I__3163 (
            .O(N__16066),
            .I(N__16063));
    LocalMux I__3162 (
            .O(N__16063),
            .I(\transmit_module.X_DELTA_PATTERN_10 ));
    InMux I__3161 (
            .O(N__16060),
            .I(N__16057));
    LocalMux I__3160 (
            .O(N__16057),
            .I(N__16054));
    Odrv12 I__3159 (
            .O(N__16054),
            .I(\line_buffer.n4072 ));
    InMux I__3158 (
            .O(N__16051),
            .I(N__16048));
    LocalMux I__3157 (
            .O(N__16048),
            .I(N__16045));
    Span4Mux_v I__3156 (
            .O(N__16045),
            .I(N__16042));
    Odrv4 I__3155 (
            .O(N__16042),
            .I(\line_buffer.n4134 ));
    CEMux I__3154 (
            .O(N__16039),
            .I(N__16033));
    CEMux I__3153 (
            .O(N__16038),
            .I(N__16030));
    CEMux I__3152 (
            .O(N__16037),
            .I(N__16026));
    CEMux I__3151 (
            .O(N__16036),
            .I(N__16022));
    LocalMux I__3150 (
            .O(N__16033),
            .I(N__16019));
    LocalMux I__3149 (
            .O(N__16030),
            .I(N__16016));
    CEMux I__3148 (
            .O(N__16029),
            .I(N__16013));
    LocalMux I__3147 (
            .O(N__16026),
            .I(N__16010));
    SRMux I__3146 (
            .O(N__16025),
            .I(N__16007));
    LocalMux I__3145 (
            .O(N__16022),
            .I(N__16004));
    Span4Mux_h I__3144 (
            .O(N__16019),
            .I(N__16001));
    Span4Mux_v I__3143 (
            .O(N__16016),
            .I(N__15996));
    LocalMux I__3142 (
            .O(N__16013),
            .I(N__15996));
    Span4Mux_v I__3141 (
            .O(N__16010),
            .I(N__15993));
    LocalMux I__3140 (
            .O(N__16007),
            .I(N__15990));
    Span4Mux_v I__3139 (
            .O(N__16004),
            .I(N__15983));
    Span4Mux_v I__3138 (
            .O(N__16001),
            .I(N__15983));
    Span4Mux_h I__3137 (
            .O(N__15996),
            .I(N__15983));
    Span4Mux_h I__3136 (
            .O(N__15993),
            .I(N__15978));
    Span4Mux_v I__3135 (
            .O(N__15990),
            .I(N__15978));
    Odrv4 I__3134 (
            .O(N__15983),
            .I(\transmit_module.n2361 ));
    Odrv4 I__3133 (
            .O(N__15978),
            .I(\transmit_module.n2361 ));
    InMux I__3132 (
            .O(N__15973),
            .I(\receive_module.rx_counter.n3722 ));
    InMux I__3131 (
            .O(N__15970),
            .I(\receive_module.rx_counter.n3723 ));
    InMux I__3130 (
            .O(N__15967),
            .I(\receive_module.rx_counter.n3724 ));
    InMux I__3129 (
            .O(N__15964),
            .I(\receive_module.rx_counter.n3725 ));
    InMux I__3128 (
            .O(N__15961),
            .I(\receive_module.rx_counter.n3726 ));
    InMux I__3127 (
            .O(N__15958),
            .I(bfn_14_10_0_));
    InMux I__3126 (
            .O(N__15955),
            .I(\receive_module.rx_counter.n3728 ));
    SRMux I__3125 (
            .O(N__15952),
            .I(N__15949));
    LocalMux I__3124 (
            .O(N__15949),
            .I(N__15945));
    SRMux I__3123 (
            .O(N__15948),
            .I(N__15942));
    Span4Mux_v I__3122 (
            .O(N__15945),
            .I(N__15939));
    LocalMux I__3121 (
            .O(N__15942),
            .I(N__15934));
    Span4Mux_v I__3120 (
            .O(N__15939),
            .I(N__15934));
    Odrv4 I__3119 (
            .O(N__15934),
            .I(n4214));
    CascadeMux I__3118 (
            .O(N__15931),
            .I(N__15924));
    InMux I__3117 (
            .O(N__15930),
            .I(N__15918));
    InMux I__3116 (
            .O(N__15929),
            .I(N__15915));
    InMux I__3115 (
            .O(N__15928),
            .I(N__15908));
    InMux I__3114 (
            .O(N__15927),
            .I(N__15908));
    InMux I__3113 (
            .O(N__15924),
            .I(N__15908));
    InMux I__3112 (
            .O(N__15923),
            .I(N__15901));
    InMux I__3111 (
            .O(N__15922),
            .I(N__15901));
    InMux I__3110 (
            .O(N__15921),
            .I(N__15901));
    LocalMux I__3109 (
            .O(N__15918),
            .I(RX_ADDR_11));
    LocalMux I__3108 (
            .O(N__15915),
            .I(RX_ADDR_11));
    LocalMux I__3107 (
            .O(N__15908),
            .I(RX_ADDR_11));
    LocalMux I__3106 (
            .O(N__15901),
            .I(RX_ADDR_11));
    InMux I__3105 (
            .O(N__15892),
            .I(N__15882));
    InMux I__3104 (
            .O(N__15891),
            .I(N__15879));
    InMux I__3103 (
            .O(N__15890),
            .I(N__15872));
    InMux I__3102 (
            .O(N__15889),
            .I(N__15872));
    InMux I__3101 (
            .O(N__15888),
            .I(N__15872));
    InMux I__3100 (
            .O(N__15887),
            .I(N__15865));
    InMux I__3099 (
            .O(N__15886),
            .I(N__15865));
    InMux I__3098 (
            .O(N__15885),
            .I(N__15865));
    LocalMux I__3097 (
            .O(N__15882),
            .I(RX_ADDR_12));
    LocalMux I__3096 (
            .O(N__15879),
            .I(RX_ADDR_12));
    LocalMux I__3095 (
            .O(N__15872),
            .I(RX_ADDR_12));
    LocalMux I__3094 (
            .O(N__15865),
            .I(RX_ADDR_12));
    IoInMux I__3093 (
            .O(N__15856),
            .I(N__15853));
    LocalMux I__3092 (
            .O(N__15853),
            .I(N__15849));
    CascadeMux I__3091 (
            .O(N__15852),
            .I(N__15845));
    Span4Mux_s2_h I__3090 (
            .O(N__15849),
            .I(N__15839));
    CascadeMux I__3089 (
            .O(N__15848),
            .I(N__15836));
    InMux I__3088 (
            .O(N__15845),
            .I(N__15833));
    CascadeMux I__3087 (
            .O(N__15844),
            .I(N__15830));
    CascadeMux I__3086 (
            .O(N__15843),
            .I(N__15827));
    CascadeMux I__3085 (
            .O(N__15842),
            .I(N__15824));
    Span4Mux_h I__3084 (
            .O(N__15839),
            .I(N__15821));
    InMux I__3083 (
            .O(N__15836),
            .I(N__15818));
    LocalMux I__3082 (
            .O(N__15833),
            .I(N__15815));
    InMux I__3081 (
            .O(N__15830),
            .I(N__15808));
    InMux I__3080 (
            .O(N__15827),
            .I(N__15808));
    InMux I__3079 (
            .O(N__15824),
            .I(N__15808));
    Span4Mux_h I__3078 (
            .O(N__15821),
            .I(N__15803));
    LocalMux I__3077 (
            .O(N__15818),
            .I(N__15796));
    Span4Mux_v I__3076 (
            .O(N__15815),
            .I(N__15796));
    LocalMux I__3075 (
            .O(N__15808),
            .I(N__15796));
    CascadeMux I__3074 (
            .O(N__15807),
            .I(N__15792));
    CascadeMux I__3073 (
            .O(N__15806),
            .I(N__15789));
    Sp12to4 I__3072 (
            .O(N__15803),
            .I(N__15786));
    Span4Mux_h I__3071 (
            .O(N__15796),
            .I(N__15783));
    InMux I__3070 (
            .O(N__15795),
            .I(N__15776));
    InMux I__3069 (
            .O(N__15792),
            .I(N__15776));
    InMux I__3068 (
            .O(N__15789),
            .I(N__15776));
    Odrv12 I__3067 (
            .O(N__15786),
            .I(DEBUG_c_5));
    Odrv4 I__3066 (
            .O(N__15783),
            .I(DEBUG_c_5));
    LocalMux I__3065 (
            .O(N__15776),
            .I(DEBUG_c_5));
    IoInMux I__3064 (
            .O(N__15769),
            .I(N__15766));
    LocalMux I__3063 (
            .O(N__15766),
            .I(N__15763));
    Span12Mux_s9_h I__3062 (
            .O(N__15763),
            .I(N__15752));
    InMux I__3061 (
            .O(N__15762),
            .I(N__15749));
    InMux I__3060 (
            .O(N__15761),
            .I(N__15746));
    InMux I__3059 (
            .O(N__15760),
            .I(N__15739));
    InMux I__3058 (
            .O(N__15759),
            .I(N__15739));
    InMux I__3057 (
            .O(N__15758),
            .I(N__15739));
    InMux I__3056 (
            .O(N__15757),
            .I(N__15732));
    InMux I__3055 (
            .O(N__15756),
            .I(N__15732));
    InMux I__3054 (
            .O(N__15755),
            .I(N__15732));
    Odrv12 I__3053 (
            .O(N__15752),
            .I(DEBUG_c_3));
    LocalMux I__3052 (
            .O(N__15749),
            .I(DEBUG_c_3));
    LocalMux I__3051 (
            .O(N__15746),
            .I(DEBUG_c_3));
    LocalMux I__3050 (
            .O(N__15739),
            .I(DEBUG_c_3));
    LocalMux I__3049 (
            .O(N__15732),
            .I(DEBUG_c_3));
    SRMux I__3048 (
            .O(N__15721),
            .I(N__15716));
    SRMux I__3047 (
            .O(N__15720),
            .I(N__15713));
    SRMux I__3046 (
            .O(N__15719),
            .I(N__15709));
    LocalMux I__3045 (
            .O(N__15716),
            .I(N__15704));
    LocalMux I__3044 (
            .O(N__15713),
            .I(N__15704));
    SRMux I__3043 (
            .O(N__15712),
            .I(N__15701));
    LocalMux I__3042 (
            .O(N__15709),
            .I(N__15698));
    Span4Mux_v I__3041 (
            .O(N__15704),
            .I(N__15693));
    LocalMux I__3040 (
            .O(N__15701),
            .I(N__15693));
    Span4Mux_v I__3039 (
            .O(N__15698),
            .I(N__15690));
    Span4Mux_h I__3038 (
            .O(N__15693),
            .I(N__15687));
    Sp12to4 I__3037 (
            .O(N__15690),
            .I(N__15684));
    Span4Mux_h I__3036 (
            .O(N__15687),
            .I(N__15681));
    Span12Mux_h I__3035 (
            .O(N__15684),
            .I(N__15678));
    Span4Mux_h I__3034 (
            .O(N__15681),
            .I(N__15675));
    Odrv12 I__3033 (
            .O(N__15678),
            .I(n658));
    Odrv4 I__3032 (
            .O(N__15675),
            .I(n658));
    CascadeMux I__3031 (
            .O(N__15670),
            .I(N__15667));
    InMux I__3030 (
            .O(N__15667),
            .I(N__15664));
    LocalMux I__3029 (
            .O(N__15664),
            .I(N__15661));
    Span4Mux_v I__3028 (
            .O(N__15661),
            .I(N__15658));
    Span4Mux_v I__3027 (
            .O(N__15658),
            .I(N__15655));
    Odrv4 I__3026 (
            .O(N__15655),
            .I(\line_buffer.n4101 ));
    CascadeMux I__3025 (
            .O(N__15652),
            .I(N__15649));
    CascadeBuf I__3024 (
            .O(N__15649),
            .I(N__15645));
    CascadeMux I__3023 (
            .O(N__15648),
            .I(N__15642));
    CascadeMux I__3022 (
            .O(N__15645),
            .I(N__15639));
    CascadeBuf I__3021 (
            .O(N__15642),
            .I(N__15636));
    CascadeBuf I__3020 (
            .O(N__15639),
            .I(N__15633));
    CascadeMux I__3019 (
            .O(N__15636),
            .I(N__15630));
    CascadeMux I__3018 (
            .O(N__15633),
            .I(N__15627));
    CascadeBuf I__3017 (
            .O(N__15630),
            .I(N__15624));
    CascadeBuf I__3016 (
            .O(N__15627),
            .I(N__15621));
    CascadeMux I__3015 (
            .O(N__15624),
            .I(N__15618));
    CascadeMux I__3014 (
            .O(N__15621),
            .I(N__15615));
    CascadeBuf I__3013 (
            .O(N__15618),
            .I(N__15612));
    CascadeBuf I__3012 (
            .O(N__15615),
            .I(N__15609));
    CascadeMux I__3011 (
            .O(N__15612),
            .I(N__15606));
    CascadeMux I__3010 (
            .O(N__15609),
            .I(N__15603));
    CascadeBuf I__3009 (
            .O(N__15606),
            .I(N__15600));
    CascadeBuf I__3008 (
            .O(N__15603),
            .I(N__15597));
    CascadeMux I__3007 (
            .O(N__15600),
            .I(N__15594));
    CascadeMux I__3006 (
            .O(N__15597),
            .I(N__15591));
    CascadeBuf I__3005 (
            .O(N__15594),
            .I(N__15588));
    CascadeBuf I__3004 (
            .O(N__15591),
            .I(N__15585));
    CascadeMux I__3003 (
            .O(N__15588),
            .I(N__15582));
    CascadeMux I__3002 (
            .O(N__15585),
            .I(N__15579));
    CascadeBuf I__3001 (
            .O(N__15582),
            .I(N__15576));
    CascadeBuf I__3000 (
            .O(N__15579),
            .I(N__15573));
    CascadeMux I__2999 (
            .O(N__15576),
            .I(N__15570));
    CascadeMux I__2998 (
            .O(N__15573),
            .I(N__15567));
    CascadeBuf I__2997 (
            .O(N__15570),
            .I(N__15564));
    CascadeBuf I__2996 (
            .O(N__15567),
            .I(N__15561));
    CascadeMux I__2995 (
            .O(N__15564),
            .I(N__15558));
    CascadeMux I__2994 (
            .O(N__15561),
            .I(N__15555));
    CascadeBuf I__2993 (
            .O(N__15558),
            .I(N__15552));
    CascadeBuf I__2992 (
            .O(N__15555),
            .I(N__15549));
    CascadeMux I__2991 (
            .O(N__15552),
            .I(N__15546));
    CascadeMux I__2990 (
            .O(N__15549),
            .I(N__15543));
    CascadeBuf I__2989 (
            .O(N__15546),
            .I(N__15540));
    CascadeBuf I__2988 (
            .O(N__15543),
            .I(N__15537));
    CascadeMux I__2987 (
            .O(N__15540),
            .I(N__15534));
    CascadeMux I__2986 (
            .O(N__15537),
            .I(N__15531));
    CascadeBuf I__2985 (
            .O(N__15534),
            .I(N__15528));
    CascadeBuf I__2984 (
            .O(N__15531),
            .I(N__15525));
    CascadeMux I__2983 (
            .O(N__15528),
            .I(N__15522));
    CascadeMux I__2982 (
            .O(N__15525),
            .I(N__15519));
    CascadeBuf I__2981 (
            .O(N__15522),
            .I(N__15516));
    CascadeBuf I__2980 (
            .O(N__15519),
            .I(N__15513));
    CascadeMux I__2979 (
            .O(N__15516),
            .I(N__15510));
    CascadeMux I__2978 (
            .O(N__15513),
            .I(N__15507));
    CascadeBuf I__2977 (
            .O(N__15510),
            .I(N__15504));
    CascadeBuf I__2976 (
            .O(N__15507),
            .I(N__15501));
    CascadeMux I__2975 (
            .O(N__15504),
            .I(N__15498));
    CascadeMux I__2974 (
            .O(N__15501),
            .I(N__15495));
    CascadeBuf I__2973 (
            .O(N__15498),
            .I(N__15492));
    CascadeBuf I__2972 (
            .O(N__15495),
            .I(N__15489));
    CascadeMux I__2971 (
            .O(N__15492),
            .I(N__15486));
    CascadeMux I__2970 (
            .O(N__15489),
            .I(N__15483));
    CascadeBuf I__2969 (
            .O(N__15486),
            .I(N__15480));
    CascadeBuf I__2968 (
            .O(N__15483),
            .I(N__15477));
    CascadeMux I__2967 (
            .O(N__15480),
            .I(N__15474));
    CascadeMux I__2966 (
            .O(N__15477),
            .I(N__15471));
    CascadeBuf I__2965 (
            .O(N__15474),
            .I(N__15468));
    InMux I__2964 (
            .O(N__15471),
            .I(N__15465));
    CascadeMux I__2963 (
            .O(N__15468),
            .I(N__15462));
    LocalMux I__2962 (
            .O(N__15465),
            .I(N__15459));
    InMux I__2961 (
            .O(N__15462),
            .I(N__15456));
    Span12Mux_s10_h I__2960 (
            .O(N__15459),
            .I(N__15453));
    LocalMux I__2959 (
            .O(N__15456),
            .I(N__15450));
    Odrv12 I__2958 (
            .O(N__15453),
            .I(n22));
    Odrv12 I__2957 (
            .O(N__15450),
            .I(n22));
    CascadeMux I__2956 (
            .O(N__15445),
            .I(\receive_module.rx_counter.n5_cascade_ ));
    InMux I__2955 (
            .O(N__15442),
            .I(N__15435));
    InMux I__2954 (
            .O(N__15441),
            .I(N__15435));
    InMux I__2953 (
            .O(N__15440),
            .I(N__15432));
    LocalMux I__2952 (
            .O(N__15435),
            .I(N__15429));
    LocalMux I__2951 (
            .O(N__15432),
            .I(N__15426));
    Span4Mux_h I__2950 (
            .O(N__15429),
            .I(N__15423));
    Span4Mux_h I__2949 (
            .O(N__15426),
            .I(N__15420));
    Span4Mux_h I__2948 (
            .O(N__15423),
            .I(N__15417));
    Span4Mux_h I__2947 (
            .O(N__15420),
            .I(N__15414));
    Sp12to4 I__2946 (
            .O(N__15417),
            .I(N__15411));
    Span4Mux_v I__2945 (
            .O(N__15414),
            .I(N__15408));
    Odrv12 I__2944 (
            .O(N__15411),
            .I(TVP_HSYNC_c));
    Odrv4 I__2943 (
            .O(N__15408),
            .I(TVP_HSYNC_c));
    InMux I__2942 (
            .O(N__15403),
            .I(N__15400));
    LocalMux I__2941 (
            .O(N__15400),
            .I(\receive_module.rx_counter.n4_adj_576 ));
    CascadeMux I__2940 (
            .O(N__15397),
            .I(N__15393));
    CascadeMux I__2939 (
            .O(N__15396),
            .I(N__15390));
    CascadeBuf I__2938 (
            .O(N__15393),
            .I(N__15387));
    CascadeBuf I__2937 (
            .O(N__15390),
            .I(N__15384));
    CascadeMux I__2936 (
            .O(N__15387),
            .I(N__15381));
    CascadeMux I__2935 (
            .O(N__15384),
            .I(N__15378));
    CascadeBuf I__2934 (
            .O(N__15381),
            .I(N__15375));
    CascadeBuf I__2933 (
            .O(N__15378),
            .I(N__15372));
    CascadeMux I__2932 (
            .O(N__15375),
            .I(N__15369));
    CascadeMux I__2931 (
            .O(N__15372),
            .I(N__15366));
    CascadeBuf I__2930 (
            .O(N__15369),
            .I(N__15363));
    CascadeBuf I__2929 (
            .O(N__15366),
            .I(N__15360));
    CascadeMux I__2928 (
            .O(N__15363),
            .I(N__15357));
    CascadeMux I__2927 (
            .O(N__15360),
            .I(N__15354));
    CascadeBuf I__2926 (
            .O(N__15357),
            .I(N__15351));
    CascadeBuf I__2925 (
            .O(N__15354),
            .I(N__15348));
    CascadeMux I__2924 (
            .O(N__15351),
            .I(N__15345));
    CascadeMux I__2923 (
            .O(N__15348),
            .I(N__15342));
    CascadeBuf I__2922 (
            .O(N__15345),
            .I(N__15339));
    CascadeBuf I__2921 (
            .O(N__15342),
            .I(N__15336));
    CascadeMux I__2920 (
            .O(N__15339),
            .I(N__15333));
    CascadeMux I__2919 (
            .O(N__15336),
            .I(N__15330));
    CascadeBuf I__2918 (
            .O(N__15333),
            .I(N__15327));
    CascadeBuf I__2917 (
            .O(N__15330),
            .I(N__15324));
    CascadeMux I__2916 (
            .O(N__15327),
            .I(N__15321));
    CascadeMux I__2915 (
            .O(N__15324),
            .I(N__15318));
    CascadeBuf I__2914 (
            .O(N__15321),
            .I(N__15315));
    CascadeBuf I__2913 (
            .O(N__15318),
            .I(N__15312));
    CascadeMux I__2912 (
            .O(N__15315),
            .I(N__15309));
    CascadeMux I__2911 (
            .O(N__15312),
            .I(N__15306));
    CascadeBuf I__2910 (
            .O(N__15309),
            .I(N__15303));
    CascadeBuf I__2909 (
            .O(N__15306),
            .I(N__15300));
    CascadeMux I__2908 (
            .O(N__15303),
            .I(N__15297));
    CascadeMux I__2907 (
            .O(N__15300),
            .I(N__15294));
    CascadeBuf I__2906 (
            .O(N__15297),
            .I(N__15291));
    CascadeBuf I__2905 (
            .O(N__15294),
            .I(N__15288));
    CascadeMux I__2904 (
            .O(N__15291),
            .I(N__15285));
    CascadeMux I__2903 (
            .O(N__15288),
            .I(N__15282));
    CascadeBuf I__2902 (
            .O(N__15285),
            .I(N__15279));
    CascadeBuf I__2901 (
            .O(N__15282),
            .I(N__15276));
    CascadeMux I__2900 (
            .O(N__15279),
            .I(N__15273));
    CascadeMux I__2899 (
            .O(N__15276),
            .I(N__15270));
    CascadeBuf I__2898 (
            .O(N__15273),
            .I(N__15267));
    CascadeBuf I__2897 (
            .O(N__15270),
            .I(N__15264));
    CascadeMux I__2896 (
            .O(N__15267),
            .I(N__15261));
    CascadeMux I__2895 (
            .O(N__15264),
            .I(N__15258));
    CascadeBuf I__2894 (
            .O(N__15261),
            .I(N__15255));
    CascadeBuf I__2893 (
            .O(N__15258),
            .I(N__15252));
    CascadeMux I__2892 (
            .O(N__15255),
            .I(N__15249));
    CascadeMux I__2891 (
            .O(N__15252),
            .I(N__15246));
    CascadeBuf I__2890 (
            .O(N__15249),
            .I(N__15243));
    CascadeBuf I__2889 (
            .O(N__15246),
            .I(N__15240));
    CascadeMux I__2888 (
            .O(N__15243),
            .I(N__15237));
    CascadeMux I__2887 (
            .O(N__15240),
            .I(N__15234));
    CascadeBuf I__2886 (
            .O(N__15237),
            .I(N__15231));
    CascadeBuf I__2885 (
            .O(N__15234),
            .I(N__15228));
    CascadeMux I__2884 (
            .O(N__15231),
            .I(N__15225));
    CascadeMux I__2883 (
            .O(N__15228),
            .I(N__15222));
    CascadeBuf I__2882 (
            .O(N__15225),
            .I(N__15219));
    CascadeBuf I__2881 (
            .O(N__15222),
            .I(N__15216));
    CascadeMux I__2880 (
            .O(N__15219),
            .I(N__15213));
    CascadeMux I__2879 (
            .O(N__15216),
            .I(N__15210));
    InMux I__2878 (
            .O(N__15213),
            .I(N__15207));
    InMux I__2877 (
            .O(N__15210),
            .I(N__15204));
    LocalMux I__2876 (
            .O(N__15207),
            .I(N__15201));
    LocalMux I__2875 (
            .O(N__15204),
            .I(N__15198));
    Span4Mux_s3_v I__2874 (
            .O(N__15201),
            .I(N__15195));
    Span4Mux_s3_v I__2873 (
            .O(N__15198),
            .I(N__15192));
    Sp12to4 I__2872 (
            .O(N__15195),
            .I(N__15189));
    Sp12to4 I__2871 (
            .O(N__15192),
            .I(N__15186));
    Span12Mux_h I__2870 (
            .O(N__15189),
            .I(N__15182));
    Span12Mux_v I__2869 (
            .O(N__15186),
            .I(N__15179));
    InMux I__2868 (
            .O(N__15185),
            .I(N__15176));
    Span12Mux_v I__2867 (
            .O(N__15182),
            .I(N__15171));
    Span12Mux_h I__2866 (
            .O(N__15179),
            .I(N__15171));
    LocalMux I__2865 (
            .O(N__15176),
            .I(RX_ADDR_0));
    Odrv12 I__2864 (
            .O(N__15171),
            .I(RX_ADDR_0));
    InMux I__2863 (
            .O(N__15166),
            .I(bfn_14_9_0_));
    CascadeMux I__2862 (
            .O(N__15163),
            .I(N__15159));
    CascadeMux I__2861 (
            .O(N__15162),
            .I(N__15156));
    CascadeBuf I__2860 (
            .O(N__15159),
            .I(N__15153));
    CascadeBuf I__2859 (
            .O(N__15156),
            .I(N__15150));
    CascadeMux I__2858 (
            .O(N__15153),
            .I(N__15147));
    CascadeMux I__2857 (
            .O(N__15150),
            .I(N__15144));
    CascadeBuf I__2856 (
            .O(N__15147),
            .I(N__15141));
    CascadeBuf I__2855 (
            .O(N__15144),
            .I(N__15138));
    CascadeMux I__2854 (
            .O(N__15141),
            .I(N__15135));
    CascadeMux I__2853 (
            .O(N__15138),
            .I(N__15132));
    CascadeBuf I__2852 (
            .O(N__15135),
            .I(N__15129));
    CascadeBuf I__2851 (
            .O(N__15132),
            .I(N__15126));
    CascadeMux I__2850 (
            .O(N__15129),
            .I(N__15123));
    CascadeMux I__2849 (
            .O(N__15126),
            .I(N__15120));
    CascadeBuf I__2848 (
            .O(N__15123),
            .I(N__15117));
    CascadeBuf I__2847 (
            .O(N__15120),
            .I(N__15114));
    CascadeMux I__2846 (
            .O(N__15117),
            .I(N__15111));
    CascadeMux I__2845 (
            .O(N__15114),
            .I(N__15108));
    CascadeBuf I__2844 (
            .O(N__15111),
            .I(N__15105));
    CascadeBuf I__2843 (
            .O(N__15108),
            .I(N__15102));
    CascadeMux I__2842 (
            .O(N__15105),
            .I(N__15099));
    CascadeMux I__2841 (
            .O(N__15102),
            .I(N__15096));
    CascadeBuf I__2840 (
            .O(N__15099),
            .I(N__15093));
    CascadeBuf I__2839 (
            .O(N__15096),
            .I(N__15090));
    CascadeMux I__2838 (
            .O(N__15093),
            .I(N__15087));
    CascadeMux I__2837 (
            .O(N__15090),
            .I(N__15084));
    CascadeBuf I__2836 (
            .O(N__15087),
            .I(N__15081));
    CascadeBuf I__2835 (
            .O(N__15084),
            .I(N__15078));
    CascadeMux I__2834 (
            .O(N__15081),
            .I(N__15075));
    CascadeMux I__2833 (
            .O(N__15078),
            .I(N__15072));
    CascadeBuf I__2832 (
            .O(N__15075),
            .I(N__15069));
    CascadeBuf I__2831 (
            .O(N__15072),
            .I(N__15066));
    CascadeMux I__2830 (
            .O(N__15069),
            .I(N__15063));
    CascadeMux I__2829 (
            .O(N__15066),
            .I(N__15060));
    CascadeBuf I__2828 (
            .O(N__15063),
            .I(N__15057));
    CascadeBuf I__2827 (
            .O(N__15060),
            .I(N__15054));
    CascadeMux I__2826 (
            .O(N__15057),
            .I(N__15051));
    CascadeMux I__2825 (
            .O(N__15054),
            .I(N__15048));
    CascadeBuf I__2824 (
            .O(N__15051),
            .I(N__15045));
    CascadeBuf I__2823 (
            .O(N__15048),
            .I(N__15042));
    CascadeMux I__2822 (
            .O(N__15045),
            .I(N__15039));
    CascadeMux I__2821 (
            .O(N__15042),
            .I(N__15036));
    CascadeBuf I__2820 (
            .O(N__15039),
            .I(N__15033));
    CascadeBuf I__2819 (
            .O(N__15036),
            .I(N__15030));
    CascadeMux I__2818 (
            .O(N__15033),
            .I(N__15027));
    CascadeMux I__2817 (
            .O(N__15030),
            .I(N__15024));
    CascadeBuf I__2816 (
            .O(N__15027),
            .I(N__15021));
    CascadeBuf I__2815 (
            .O(N__15024),
            .I(N__15018));
    CascadeMux I__2814 (
            .O(N__15021),
            .I(N__15015));
    CascadeMux I__2813 (
            .O(N__15018),
            .I(N__15012));
    CascadeBuf I__2812 (
            .O(N__15015),
            .I(N__15009));
    CascadeBuf I__2811 (
            .O(N__15012),
            .I(N__15006));
    CascadeMux I__2810 (
            .O(N__15009),
            .I(N__15003));
    CascadeMux I__2809 (
            .O(N__15006),
            .I(N__15000));
    CascadeBuf I__2808 (
            .O(N__15003),
            .I(N__14997));
    CascadeBuf I__2807 (
            .O(N__15000),
            .I(N__14994));
    CascadeMux I__2806 (
            .O(N__14997),
            .I(N__14991));
    CascadeMux I__2805 (
            .O(N__14994),
            .I(N__14988));
    CascadeBuf I__2804 (
            .O(N__14991),
            .I(N__14985));
    CascadeBuf I__2803 (
            .O(N__14988),
            .I(N__14982));
    CascadeMux I__2802 (
            .O(N__14985),
            .I(N__14979));
    CascadeMux I__2801 (
            .O(N__14982),
            .I(N__14976));
    InMux I__2800 (
            .O(N__14979),
            .I(N__14973));
    InMux I__2799 (
            .O(N__14976),
            .I(N__14970));
    LocalMux I__2798 (
            .O(N__14973),
            .I(N__14967));
    LocalMux I__2797 (
            .O(N__14970),
            .I(N__14964));
    Span4Mux_s2_v I__2796 (
            .O(N__14967),
            .I(N__14961));
    Sp12to4 I__2795 (
            .O(N__14964),
            .I(N__14958));
    Sp12to4 I__2794 (
            .O(N__14961),
            .I(N__14955));
    Span12Mux_s11_v I__2793 (
            .O(N__14958),
            .I(N__14951));
    Span12Mux_h I__2792 (
            .O(N__14955),
            .I(N__14948));
    InMux I__2791 (
            .O(N__14954),
            .I(N__14945));
    Span12Mux_v I__2790 (
            .O(N__14951),
            .I(N__14942));
    Span12Mux_v I__2789 (
            .O(N__14948),
            .I(N__14939));
    LocalMux I__2788 (
            .O(N__14945),
            .I(RX_ADDR_1));
    Odrv12 I__2787 (
            .O(N__14942),
            .I(RX_ADDR_1));
    Odrv12 I__2786 (
            .O(N__14939),
            .I(RX_ADDR_1));
    InMux I__2785 (
            .O(N__14932),
            .I(\receive_module.rx_counter.n3720 ));
    CascadeMux I__2784 (
            .O(N__14929),
            .I(N__14926));
    CascadeBuf I__2783 (
            .O(N__14926),
            .I(N__14922));
    CascadeMux I__2782 (
            .O(N__14925),
            .I(N__14919));
    CascadeMux I__2781 (
            .O(N__14922),
            .I(N__14916));
    CascadeBuf I__2780 (
            .O(N__14919),
            .I(N__14913));
    CascadeBuf I__2779 (
            .O(N__14916),
            .I(N__14910));
    CascadeMux I__2778 (
            .O(N__14913),
            .I(N__14907));
    CascadeMux I__2777 (
            .O(N__14910),
            .I(N__14904));
    CascadeBuf I__2776 (
            .O(N__14907),
            .I(N__14901));
    CascadeBuf I__2775 (
            .O(N__14904),
            .I(N__14898));
    CascadeMux I__2774 (
            .O(N__14901),
            .I(N__14895));
    CascadeMux I__2773 (
            .O(N__14898),
            .I(N__14892));
    CascadeBuf I__2772 (
            .O(N__14895),
            .I(N__14889));
    CascadeBuf I__2771 (
            .O(N__14892),
            .I(N__14886));
    CascadeMux I__2770 (
            .O(N__14889),
            .I(N__14883));
    CascadeMux I__2769 (
            .O(N__14886),
            .I(N__14880));
    CascadeBuf I__2768 (
            .O(N__14883),
            .I(N__14877));
    CascadeBuf I__2767 (
            .O(N__14880),
            .I(N__14874));
    CascadeMux I__2766 (
            .O(N__14877),
            .I(N__14871));
    CascadeMux I__2765 (
            .O(N__14874),
            .I(N__14868));
    CascadeBuf I__2764 (
            .O(N__14871),
            .I(N__14865));
    CascadeBuf I__2763 (
            .O(N__14868),
            .I(N__14862));
    CascadeMux I__2762 (
            .O(N__14865),
            .I(N__14859));
    CascadeMux I__2761 (
            .O(N__14862),
            .I(N__14856));
    CascadeBuf I__2760 (
            .O(N__14859),
            .I(N__14853));
    CascadeBuf I__2759 (
            .O(N__14856),
            .I(N__14850));
    CascadeMux I__2758 (
            .O(N__14853),
            .I(N__14847));
    CascadeMux I__2757 (
            .O(N__14850),
            .I(N__14844));
    CascadeBuf I__2756 (
            .O(N__14847),
            .I(N__14841));
    CascadeBuf I__2755 (
            .O(N__14844),
            .I(N__14838));
    CascadeMux I__2754 (
            .O(N__14841),
            .I(N__14835));
    CascadeMux I__2753 (
            .O(N__14838),
            .I(N__14832));
    CascadeBuf I__2752 (
            .O(N__14835),
            .I(N__14829));
    CascadeBuf I__2751 (
            .O(N__14832),
            .I(N__14826));
    CascadeMux I__2750 (
            .O(N__14829),
            .I(N__14823));
    CascadeMux I__2749 (
            .O(N__14826),
            .I(N__14820));
    CascadeBuf I__2748 (
            .O(N__14823),
            .I(N__14817));
    CascadeBuf I__2747 (
            .O(N__14820),
            .I(N__14814));
    CascadeMux I__2746 (
            .O(N__14817),
            .I(N__14811));
    CascadeMux I__2745 (
            .O(N__14814),
            .I(N__14808));
    CascadeBuf I__2744 (
            .O(N__14811),
            .I(N__14805));
    CascadeBuf I__2743 (
            .O(N__14808),
            .I(N__14802));
    CascadeMux I__2742 (
            .O(N__14805),
            .I(N__14799));
    CascadeMux I__2741 (
            .O(N__14802),
            .I(N__14796));
    CascadeBuf I__2740 (
            .O(N__14799),
            .I(N__14793));
    CascadeBuf I__2739 (
            .O(N__14796),
            .I(N__14790));
    CascadeMux I__2738 (
            .O(N__14793),
            .I(N__14787));
    CascadeMux I__2737 (
            .O(N__14790),
            .I(N__14784));
    CascadeBuf I__2736 (
            .O(N__14787),
            .I(N__14781));
    CascadeBuf I__2735 (
            .O(N__14784),
            .I(N__14778));
    CascadeMux I__2734 (
            .O(N__14781),
            .I(N__14775));
    CascadeMux I__2733 (
            .O(N__14778),
            .I(N__14772));
    CascadeBuf I__2732 (
            .O(N__14775),
            .I(N__14769));
    CascadeBuf I__2731 (
            .O(N__14772),
            .I(N__14766));
    CascadeMux I__2730 (
            .O(N__14769),
            .I(N__14763));
    CascadeMux I__2729 (
            .O(N__14766),
            .I(N__14760));
    CascadeBuf I__2728 (
            .O(N__14763),
            .I(N__14757));
    CascadeBuf I__2727 (
            .O(N__14760),
            .I(N__14754));
    CascadeMux I__2726 (
            .O(N__14757),
            .I(N__14751));
    CascadeMux I__2725 (
            .O(N__14754),
            .I(N__14748));
    CascadeBuf I__2724 (
            .O(N__14751),
            .I(N__14745));
    InMux I__2723 (
            .O(N__14748),
            .I(N__14742));
    CascadeMux I__2722 (
            .O(N__14745),
            .I(N__14739));
    LocalMux I__2721 (
            .O(N__14742),
            .I(N__14736));
    InMux I__2720 (
            .O(N__14739),
            .I(N__14733));
    Span4Mux_s3_v I__2719 (
            .O(N__14736),
            .I(N__14730));
    LocalMux I__2718 (
            .O(N__14733),
            .I(N__14727));
    Sp12to4 I__2717 (
            .O(N__14730),
            .I(N__14724));
    Span12Mux_s11_v I__2716 (
            .O(N__14727),
            .I(N__14720));
    Span12Mux_v I__2715 (
            .O(N__14724),
            .I(N__14717));
    InMux I__2714 (
            .O(N__14723),
            .I(N__14714));
    Span12Mux_v I__2713 (
            .O(N__14720),
            .I(N__14711));
    Span12Mux_h I__2712 (
            .O(N__14717),
            .I(N__14708));
    LocalMux I__2711 (
            .O(N__14714),
            .I(RX_ADDR_2));
    Odrv12 I__2710 (
            .O(N__14711),
            .I(RX_ADDR_2));
    Odrv12 I__2709 (
            .O(N__14708),
            .I(RX_ADDR_2));
    InMux I__2708 (
            .O(N__14701),
            .I(\receive_module.rx_counter.n3721 ));
    InMux I__2707 (
            .O(N__14698),
            .I(N__14695));
    LocalMux I__2706 (
            .O(N__14695),
            .I(\transmit_module.Y_DELTA_PATTERN_49 ));
    InMux I__2705 (
            .O(N__14692),
            .I(N__14689));
    LocalMux I__2704 (
            .O(N__14689),
            .I(\transmit_module.Y_DELTA_PATTERN_54 ));
    InMux I__2703 (
            .O(N__14686),
            .I(N__14683));
    LocalMux I__2702 (
            .O(N__14683),
            .I(\transmit_module.Y_DELTA_PATTERN_51 ));
    InMux I__2701 (
            .O(N__14680),
            .I(N__14677));
    LocalMux I__2700 (
            .O(N__14677),
            .I(\transmit_module.Y_DELTA_PATTERN_50 ));
    InMux I__2699 (
            .O(N__14674),
            .I(N__14671));
    LocalMux I__2698 (
            .O(N__14671),
            .I(\transmit_module.Y_DELTA_PATTERN_56 ));
    InMux I__2697 (
            .O(N__14668),
            .I(N__14665));
    LocalMux I__2696 (
            .O(N__14665),
            .I(\transmit_module.Y_DELTA_PATTERN_55 ));
    InMux I__2695 (
            .O(N__14662),
            .I(N__14659));
    LocalMux I__2694 (
            .O(N__14659),
            .I(\transmit_module.Y_DELTA_PATTERN_59 ));
    InMux I__2693 (
            .O(N__14656),
            .I(N__14653));
    LocalMux I__2692 (
            .O(N__14653),
            .I(\transmit_module.Y_DELTA_PATTERN_58 ));
    InMux I__2691 (
            .O(N__14650),
            .I(N__14647));
    LocalMux I__2690 (
            .O(N__14647),
            .I(\transmit_module.Y_DELTA_PATTERN_61 ));
    InMux I__2689 (
            .O(N__14644),
            .I(N__14641));
    LocalMux I__2688 (
            .O(N__14641),
            .I(\transmit_module.Y_DELTA_PATTERN_60 ));
    InMux I__2687 (
            .O(N__14638),
            .I(N__14635));
    LocalMux I__2686 (
            .O(N__14635),
            .I(N__14632));
    Span4Mux_h I__2685 (
            .O(N__14632),
            .I(N__14629));
    Span4Mux_h I__2684 (
            .O(N__14629),
            .I(N__14626));
    Span4Mux_h I__2683 (
            .O(N__14626),
            .I(N__14623));
    Odrv4 I__2682 (
            .O(N__14623),
            .I(\line_buffer.n558 ));
    InMux I__2681 (
            .O(N__14620),
            .I(N__14617));
    LocalMux I__2680 (
            .O(N__14617),
            .I(N__14614));
    Span4Mux_v I__2679 (
            .O(N__14614),
            .I(N__14611));
    Span4Mux_h I__2678 (
            .O(N__14611),
            .I(N__14608));
    Odrv4 I__2677 (
            .O(N__14608),
            .I(\line_buffer.n550 ));
    SRMux I__2676 (
            .O(N__14605),
            .I(N__14601));
    SRMux I__2675 (
            .O(N__14604),
            .I(N__14598));
    LocalMux I__2674 (
            .O(N__14601),
            .I(N__14595));
    LocalMux I__2673 (
            .O(N__14598),
            .I(N__14592));
    Odrv4 I__2672 (
            .O(N__14595),
            .I(n2587));
    Odrv4 I__2671 (
            .O(N__14592),
            .I(n2587));
    InMux I__2670 (
            .O(N__14587),
            .I(N__14584));
    LocalMux I__2669 (
            .O(N__14584),
            .I(\transmit_module.Y_DELTA_PATTERN_43 ));
    InMux I__2668 (
            .O(N__14581),
            .I(N__14578));
    LocalMux I__2667 (
            .O(N__14578),
            .I(\transmit_module.Y_DELTA_PATTERN_44 ));
    InMux I__2666 (
            .O(N__14575),
            .I(N__14572));
    LocalMux I__2665 (
            .O(N__14572),
            .I(\transmit_module.Y_DELTA_PATTERN_46 ));
    InMux I__2664 (
            .O(N__14569),
            .I(N__14566));
    LocalMux I__2663 (
            .O(N__14566),
            .I(\transmit_module.Y_DELTA_PATTERN_45 ));
    InMux I__2662 (
            .O(N__14563),
            .I(N__14560));
    LocalMux I__2661 (
            .O(N__14560),
            .I(\transmit_module.Y_DELTA_PATTERN_47 ));
    InMux I__2660 (
            .O(N__14557),
            .I(N__14554));
    LocalMux I__2659 (
            .O(N__14554),
            .I(\transmit_module.Y_DELTA_PATTERN_48 ));
    InMux I__2658 (
            .O(N__14551),
            .I(N__14548));
    LocalMux I__2657 (
            .O(N__14548),
            .I(\transmit_module.Y_DELTA_PATTERN_53 ));
    InMux I__2656 (
            .O(N__14545),
            .I(N__14542));
    LocalMux I__2655 (
            .O(N__14542),
            .I(\transmit_module.Y_DELTA_PATTERN_52 ));
    CascadeMux I__2654 (
            .O(N__14539),
            .I(\line_buffer.n4185_cascade_ ));
    InMux I__2653 (
            .O(N__14536),
            .I(N__14533));
    LocalMux I__2652 (
            .O(N__14533),
            .I(N__14530));
    Span4Mux_v I__2651 (
            .O(N__14530),
            .I(N__14527));
    Odrv4 I__2650 (
            .O(N__14527),
            .I(\line_buffer.n4125 ));
    IoInMux I__2649 (
            .O(N__14524),
            .I(N__14521));
    LocalMux I__2648 (
            .O(N__14521),
            .I(N__14517));
    IoInMux I__2647 (
            .O(N__14520),
            .I(N__14514));
    IoSpan4Mux I__2646 (
            .O(N__14517),
            .I(N__14508));
    LocalMux I__2645 (
            .O(N__14514),
            .I(N__14508));
    IoInMux I__2644 (
            .O(N__14513),
            .I(N__14505));
    IoSpan4Mux I__2643 (
            .O(N__14508),
            .I(N__14502));
    LocalMux I__2642 (
            .O(N__14505),
            .I(N__14499));
    Span4Mux_s0_h I__2641 (
            .O(N__14502),
            .I(N__14496));
    Span4Mux_s3_v I__2640 (
            .O(N__14499),
            .I(N__14493));
    Sp12to4 I__2639 (
            .O(N__14496),
            .I(N__14490));
    Sp12to4 I__2638 (
            .O(N__14493),
            .I(N__14487));
    Span12Mux_h I__2637 (
            .O(N__14490),
            .I(N__14482));
    Span12Mux_h I__2636 (
            .O(N__14487),
            .I(N__14482));
    Odrv12 I__2635 (
            .O(N__14482),
            .I(n1995));
    InMux I__2634 (
            .O(N__14479),
            .I(N__14476));
    LocalMux I__2633 (
            .O(N__14476),
            .I(N__14473));
    Span4Mux_h I__2632 (
            .O(N__14473),
            .I(N__14470));
    Span4Mux_v I__2631 (
            .O(N__14470),
            .I(N__14467));
    Odrv4 I__2630 (
            .O(N__14467),
            .I(TX_DATA_2));
    IoInMux I__2629 (
            .O(N__14464),
            .I(N__14459));
    IoInMux I__2628 (
            .O(N__14463),
            .I(N__14456));
    IoInMux I__2627 (
            .O(N__14462),
            .I(N__14453));
    LocalMux I__2626 (
            .O(N__14459),
            .I(N__14450));
    LocalMux I__2625 (
            .O(N__14456),
            .I(N__14447));
    LocalMux I__2624 (
            .O(N__14453),
            .I(N__14444));
    Span4Mux_s2_v I__2623 (
            .O(N__14450),
            .I(N__14441));
    Span4Mux_s2_v I__2622 (
            .O(N__14447),
            .I(N__14438));
    IoSpan4Mux I__2621 (
            .O(N__14444),
            .I(N__14435));
    Sp12to4 I__2620 (
            .O(N__14441),
            .I(N__14432));
    Sp12to4 I__2619 (
            .O(N__14438),
            .I(N__14429));
    Sp12to4 I__2618 (
            .O(N__14435),
            .I(N__14426));
    Span12Mux_h I__2617 (
            .O(N__14432),
            .I(N__14419));
    Span12Mux_h I__2616 (
            .O(N__14429),
            .I(N__14419));
    Span12Mux_h I__2615 (
            .O(N__14426),
            .I(N__14419));
    Odrv12 I__2614 (
            .O(N__14419),
            .I(n1994));
    IoInMux I__2613 (
            .O(N__14416),
            .I(N__14412));
    IoInMux I__2612 (
            .O(N__14415),
            .I(N__14408));
    LocalMux I__2611 (
            .O(N__14412),
            .I(N__14405));
    IoInMux I__2610 (
            .O(N__14411),
            .I(N__14402));
    LocalMux I__2609 (
            .O(N__14408),
            .I(N__14399));
    IoSpan4Mux I__2608 (
            .O(N__14405),
            .I(N__14396));
    LocalMux I__2607 (
            .O(N__14402),
            .I(N__14393));
    IoSpan4Mux I__2606 (
            .O(N__14399),
            .I(N__14390));
    Sp12to4 I__2605 (
            .O(N__14396),
            .I(N__14387));
    IoSpan4Mux I__2604 (
            .O(N__14393),
            .I(N__14384));
    Span4Mux_s3_h I__2603 (
            .O(N__14390),
            .I(N__14381));
    Span12Mux_v I__2602 (
            .O(N__14387),
            .I(N__14378));
    Sp12to4 I__2601 (
            .O(N__14384),
            .I(N__14375));
    Span4Mux_h I__2600 (
            .O(N__14381),
            .I(N__14372));
    Span12Mux_h I__2599 (
            .O(N__14378),
            .I(N__14367));
    Span12Mux_v I__2598 (
            .O(N__14375),
            .I(N__14367));
    Span4Mux_h I__2597 (
            .O(N__14372),
            .I(N__14364));
    Odrv12 I__2596 (
            .O(N__14367),
            .I(n1993));
    Odrv4 I__2595 (
            .O(N__14364),
            .I(n1993));
    IoInMux I__2594 (
            .O(N__14359),
            .I(N__14356));
    LocalMux I__2593 (
            .O(N__14356),
            .I(N__14353));
    Span4Mux_s0_v I__2592 (
            .O(N__14353),
            .I(N__14348));
    IoInMux I__2591 (
            .O(N__14352),
            .I(N__14345));
    IoInMux I__2590 (
            .O(N__14351),
            .I(N__14342));
    Span4Mux_v I__2589 (
            .O(N__14348),
            .I(N__14339));
    LocalMux I__2588 (
            .O(N__14345),
            .I(N__14336));
    LocalMux I__2587 (
            .O(N__14342),
            .I(N__14333));
    Span4Mux_v I__2586 (
            .O(N__14339),
            .I(N__14330));
    IoSpan4Mux I__2585 (
            .O(N__14336),
            .I(N__14327));
    Span12Mux_s0_v I__2584 (
            .O(N__14333),
            .I(N__14324));
    Sp12to4 I__2583 (
            .O(N__14330),
            .I(N__14321));
    Sp12to4 I__2582 (
            .O(N__14327),
            .I(N__14318));
    Span12Mux_v I__2581 (
            .O(N__14324),
            .I(N__14315));
    Span12Mux_h I__2580 (
            .O(N__14321),
            .I(N__14310));
    Span12Mux_h I__2579 (
            .O(N__14318),
            .I(N__14310));
    Odrv12 I__2578 (
            .O(N__14315),
            .I(n1992));
    Odrv12 I__2577 (
            .O(N__14310),
            .I(n1992));
    IoInMux I__2576 (
            .O(N__14305),
            .I(N__14301));
    IoInMux I__2575 (
            .O(N__14304),
            .I(N__14297));
    LocalMux I__2574 (
            .O(N__14301),
            .I(N__14294));
    IoInMux I__2573 (
            .O(N__14300),
            .I(N__14291));
    LocalMux I__2572 (
            .O(N__14297),
            .I(N__14288));
    Sp12to4 I__2571 (
            .O(N__14294),
            .I(N__14285));
    LocalMux I__2570 (
            .O(N__14291),
            .I(N__14282));
    IoSpan4Mux I__2569 (
            .O(N__14288),
            .I(N__14279));
    Span12Mux_v I__2568 (
            .O(N__14285),
            .I(N__14276));
    Span12Mux_s0_h I__2567 (
            .O(N__14282),
            .I(N__14273));
    Sp12to4 I__2566 (
            .O(N__14279),
            .I(N__14270));
    Span12Mux_h I__2565 (
            .O(N__14276),
            .I(N__14267));
    Span12Mux_h I__2564 (
            .O(N__14273),
            .I(N__14264));
    Span12Mux_v I__2563 (
            .O(N__14270),
            .I(N__14261));
    Odrv12 I__2562 (
            .O(N__14267),
            .I(n1991));
    Odrv12 I__2561 (
            .O(N__14264),
            .I(n1991));
    Odrv12 I__2560 (
            .O(N__14261),
            .I(n1991));
    InMux I__2559 (
            .O(N__14254),
            .I(N__14251));
    LocalMux I__2558 (
            .O(N__14251),
            .I(N__14248));
    Odrv4 I__2557 (
            .O(N__14248),
            .I(TX_DATA_6));
    IoInMux I__2556 (
            .O(N__14245),
            .I(N__14240));
    IoInMux I__2555 (
            .O(N__14244),
            .I(N__14237));
    IoInMux I__2554 (
            .O(N__14243),
            .I(N__14234));
    LocalMux I__2553 (
            .O(N__14240),
            .I(N__14231));
    LocalMux I__2552 (
            .O(N__14237),
            .I(N__14228));
    LocalMux I__2551 (
            .O(N__14234),
            .I(N__14225));
    Span4Mux_s0_v I__2550 (
            .O(N__14231),
            .I(N__14222));
    IoSpan4Mux I__2549 (
            .O(N__14228),
            .I(N__14219));
    Span4Mux_s2_h I__2548 (
            .O(N__14225),
            .I(N__14216));
    Sp12to4 I__2547 (
            .O(N__14222),
            .I(N__14213));
    Span4Mux_s0_v I__2546 (
            .O(N__14219),
            .I(N__14210));
    Sp12to4 I__2545 (
            .O(N__14216),
            .I(N__14207));
    Span12Mux_s9_h I__2544 (
            .O(N__14213),
            .I(N__14204));
    Sp12to4 I__2543 (
            .O(N__14210),
            .I(N__14201));
    Span12Mux_v I__2542 (
            .O(N__14207),
            .I(N__14198));
    Span12Mux_v I__2541 (
            .O(N__14204),
            .I(N__14193));
    Span12Mux_v I__2540 (
            .O(N__14201),
            .I(N__14193));
    Odrv12 I__2539 (
            .O(N__14198),
            .I(n1990));
    Odrv12 I__2538 (
            .O(N__14193),
            .I(n1990));
    InMux I__2537 (
            .O(N__14188),
            .I(N__14185));
    LocalMux I__2536 (
            .O(N__14185),
            .I(TX_DATA_7));
    IoInMux I__2535 (
            .O(N__14182),
            .I(N__14178));
    IoInMux I__2534 (
            .O(N__14181),
            .I(N__14175));
    LocalMux I__2533 (
            .O(N__14178),
            .I(N__14172));
    LocalMux I__2532 (
            .O(N__14175),
            .I(N__14168));
    IoSpan4Mux I__2531 (
            .O(N__14172),
            .I(N__14165));
    IoInMux I__2530 (
            .O(N__14171),
            .I(N__14162));
    IoSpan4Mux I__2529 (
            .O(N__14168),
            .I(N__14159));
    Span4Mux_s2_h I__2528 (
            .O(N__14165),
            .I(N__14156));
    LocalMux I__2527 (
            .O(N__14162),
            .I(N__14153));
    Span4Mux_s0_h I__2526 (
            .O(N__14159),
            .I(N__14150));
    Sp12to4 I__2525 (
            .O(N__14156),
            .I(N__14147));
    IoSpan4Mux I__2524 (
            .O(N__14153),
            .I(N__14144));
    Sp12to4 I__2523 (
            .O(N__14150),
            .I(N__14141));
    Span12Mux_s10_h I__2522 (
            .O(N__14147),
            .I(N__14138));
    Sp12to4 I__2521 (
            .O(N__14144),
            .I(N__14135));
    Span12Mux_h I__2520 (
            .O(N__14141),
            .I(N__14132));
    Span12Mux_v I__2519 (
            .O(N__14138),
            .I(N__14127));
    Span12Mux_v I__2518 (
            .O(N__14135),
            .I(N__14127));
    Odrv12 I__2517 (
            .O(N__14132),
            .I(ADV_B_c));
    Odrv12 I__2516 (
            .O(N__14127),
            .I(ADV_B_c));
    InMux I__2515 (
            .O(N__14122),
            .I(N__14118));
    InMux I__2514 (
            .O(N__14121),
            .I(N__14115));
    LocalMux I__2513 (
            .O(N__14118),
            .I(\transmit_module.n186 ));
    LocalMux I__2512 (
            .O(N__14115),
            .I(\transmit_module.n186 ));
    CascadeMux I__2511 (
            .O(N__14110),
            .I(\transmit_module.n4211_cascade_ ));
    InMux I__2510 (
            .O(N__14107),
            .I(N__14103));
    InMux I__2509 (
            .O(N__14106),
            .I(N__14100));
    LocalMux I__2508 (
            .O(N__14103),
            .I(\transmit_module.n217 ));
    LocalMux I__2507 (
            .O(N__14100),
            .I(\transmit_module.n217 ));
    CascadeMux I__2506 (
            .O(N__14095),
            .I(N__14091));
    CascadeMux I__2505 (
            .O(N__14094),
            .I(N__14088));
    CascadeBuf I__2504 (
            .O(N__14091),
            .I(N__14085));
    CascadeBuf I__2503 (
            .O(N__14088),
            .I(N__14082));
    CascadeMux I__2502 (
            .O(N__14085),
            .I(N__14079));
    CascadeMux I__2501 (
            .O(N__14082),
            .I(N__14076));
    CascadeBuf I__2500 (
            .O(N__14079),
            .I(N__14073));
    CascadeBuf I__2499 (
            .O(N__14076),
            .I(N__14070));
    CascadeMux I__2498 (
            .O(N__14073),
            .I(N__14067));
    CascadeMux I__2497 (
            .O(N__14070),
            .I(N__14064));
    CascadeBuf I__2496 (
            .O(N__14067),
            .I(N__14061));
    CascadeBuf I__2495 (
            .O(N__14064),
            .I(N__14058));
    CascadeMux I__2494 (
            .O(N__14061),
            .I(N__14055));
    CascadeMux I__2493 (
            .O(N__14058),
            .I(N__14052));
    CascadeBuf I__2492 (
            .O(N__14055),
            .I(N__14049));
    CascadeBuf I__2491 (
            .O(N__14052),
            .I(N__14046));
    CascadeMux I__2490 (
            .O(N__14049),
            .I(N__14043));
    CascadeMux I__2489 (
            .O(N__14046),
            .I(N__14040));
    CascadeBuf I__2488 (
            .O(N__14043),
            .I(N__14037));
    CascadeBuf I__2487 (
            .O(N__14040),
            .I(N__14034));
    CascadeMux I__2486 (
            .O(N__14037),
            .I(N__14031));
    CascadeMux I__2485 (
            .O(N__14034),
            .I(N__14028));
    CascadeBuf I__2484 (
            .O(N__14031),
            .I(N__14025));
    CascadeBuf I__2483 (
            .O(N__14028),
            .I(N__14022));
    CascadeMux I__2482 (
            .O(N__14025),
            .I(N__14019));
    CascadeMux I__2481 (
            .O(N__14022),
            .I(N__14016));
    CascadeBuf I__2480 (
            .O(N__14019),
            .I(N__14013));
    CascadeBuf I__2479 (
            .O(N__14016),
            .I(N__14010));
    CascadeMux I__2478 (
            .O(N__14013),
            .I(N__14007));
    CascadeMux I__2477 (
            .O(N__14010),
            .I(N__14004));
    CascadeBuf I__2476 (
            .O(N__14007),
            .I(N__14001));
    CascadeBuf I__2475 (
            .O(N__14004),
            .I(N__13998));
    CascadeMux I__2474 (
            .O(N__14001),
            .I(N__13995));
    CascadeMux I__2473 (
            .O(N__13998),
            .I(N__13992));
    CascadeBuf I__2472 (
            .O(N__13995),
            .I(N__13989));
    CascadeBuf I__2471 (
            .O(N__13992),
            .I(N__13986));
    CascadeMux I__2470 (
            .O(N__13989),
            .I(N__13983));
    CascadeMux I__2469 (
            .O(N__13986),
            .I(N__13980));
    CascadeBuf I__2468 (
            .O(N__13983),
            .I(N__13977));
    CascadeBuf I__2467 (
            .O(N__13980),
            .I(N__13974));
    CascadeMux I__2466 (
            .O(N__13977),
            .I(N__13971));
    CascadeMux I__2465 (
            .O(N__13974),
            .I(N__13968));
    CascadeBuf I__2464 (
            .O(N__13971),
            .I(N__13965));
    CascadeBuf I__2463 (
            .O(N__13968),
            .I(N__13962));
    CascadeMux I__2462 (
            .O(N__13965),
            .I(N__13959));
    CascadeMux I__2461 (
            .O(N__13962),
            .I(N__13956));
    CascadeBuf I__2460 (
            .O(N__13959),
            .I(N__13953));
    CascadeBuf I__2459 (
            .O(N__13956),
            .I(N__13950));
    CascadeMux I__2458 (
            .O(N__13953),
            .I(N__13947));
    CascadeMux I__2457 (
            .O(N__13950),
            .I(N__13944));
    CascadeBuf I__2456 (
            .O(N__13947),
            .I(N__13941));
    CascadeBuf I__2455 (
            .O(N__13944),
            .I(N__13938));
    CascadeMux I__2454 (
            .O(N__13941),
            .I(N__13935));
    CascadeMux I__2453 (
            .O(N__13938),
            .I(N__13932));
    CascadeBuf I__2452 (
            .O(N__13935),
            .I(N__13929));
    CascadeBuf I__2451 (
            .O(N__13932),
            .I(N__13926));
    CascadeMux I__2450 (
            .O(N__13929),
            .I(N__13923));
    CascadeMux I__2449 (
            .O(N__13926),
            .I(N__13920));
    CascadeBuf I__2448 (
            .O(N__13923),
            .I(N__13917));
    CascadeBuf I__2447 (
            .O(N__13920),
            .I(N__13914));
    CascadeMux I__2446 (
            .O(N__13917),
            .I(N__13911));
    CascadeMux I__2445 (
            .O(N__13914),
            .I(N__13908));
    InMux I__2444 (
            .O(N__13911),
            .I(N__13905));
    InMux I__2443 (
            .O(N__13908),
            .I(N__13902));
    LocalMux I__2442 (
            .O(N__13905),
            .I(N__13899));
    LocalMux I__2441 (
            .O(N__13902),
            .I(N__13896));
    Span4Mux_h I__2440 (
            .O(N__13899),
            .I(N__13893));
    Span12Mux_s10_v I__2439 (
            .O(N__13896),
            .I(N__13890));
    Span4Mux_h I__2438 (
            .O(N__13893),
            .I(N__13887));
    Span12Mux_h I__2437 (
            .O(N__13890),
            .I(N__13884));
    Sp12to4 I__2436 (
            .O(N__13887),
            .I(N__13881));
    Odrv12 I__2435 (
            .O(N__13884),
            .I(n26));
    Odrv12 I__2434 (
            .O(N__13881),
            .I(n26));
    InMux I__2433 (
            .O(N__13876),
            .I(N__13873));
    LocalMux I__2432 (
            .O(N__13873),
            .I(N__13870));
    Span12Mux_v I__2431 (
            .O(N__13870),
            .I(N__13867));
    Span12Mux_h I__2430 (
            .O(N__13867),
            .I(N__13864));
    Odrv12 I__2429 (
            .O(N__13864),
            .I(\line_buffer.n559 ));
    InMux I__2428 (
            .O(N__13861),
            .I(N__13858));
    LocalMux I__2427 (
            .O(N__13858),
            .I(N__13855));
    Odrv4 I__2426 (
            .O(N__13855),
            .I(\line_buffer.n4182 ));
    CascadeMux I__2425 (
            .O(N__13852),
            .I(N__13849));
    InMux I__2424 (
            .O(N__13849),
            .I(N__13846));
    LocalMux I__2423 (
            .O(N__13846),
            .I(N__13843));
    Span12Mux_h I__2422 (
            .O(N__13843),
            .I(N__13840));
    Odrv12 I__2421 (
            .O(N__13840),
            .I(\line_buffer.n551 ));
    InMux I__2420 (
            .O(N__13837),
            .I(N__13827));
    InMux I__2419 (
            .O(N__13836),
            .I(N__13827));
    InMux I__2418 (
            .O(N__13835),
            .I(N__13827));
    InMux I__2417 (
            .O(N__13834),
            .I(N__13824));
    LocalMux I__2416 (
            .O(N__13827),
            .I(N__13821));
    LocalMux I__2415 (
            .O(N__13824),
            .I(\transmit_module.video_signal_controller.VGA_X_9 ));
    Odrv4 I__2414 (
            .O(N__13821),
            .I(\transmit_module.video_signal_controller.VGA_X_9 ));
    InMux I__2413 (
            .O(N__13816),
            .I(\transmit_module.video_signal_controller.n3696 ));
    CascadeMux I__2412 (
            .O(N__13813),
            .I(N__13808));
    InMux I__2411 (
            .O(N__13812),
            .I(N__13804));
    InMux I__2410 (
            .O(N__13811),
            .I(N__13797));
    InMux I__2409 (
            .O(N__13808),
            .I(N__13797));
    InMux I__2408 (
            .O(N__13807),
            .I(N__13797));
    LocalMux I__2407 (
            .O(N__13804),
            .I(\transmit_module.video_signal_controller.VGA_X_10 ));
    LocalMux I__2406 (
            .O(N__13797),
            .I(\transmit_module.video_signal_controller.VGA_X_10 ));
    InMux I__2405 (
            .O(N__13792),
            .I(\transmit_module.video_signal_controller.n3697 ));
    InMux I__2404 (
            .O(N__13789),
            .I(\transmit_module.video_signal_controller.n3698 ));
    InMux I__2403 (
            .O(N__13786),
            .I(N__13780));
    InMux I__2402 (
            .O(N__13785),
            .I(N__13773));
    InMux I__2401 (
            .O(N__13784),
            .I(N__13773));
    InMux I__2400 (
            .O(N__13783),
            .I(N__13773));
    LocalMux I__2399 (
            .O(N__13780),
            .I(\transmit_module.video_signal_controller.VGA_X_11 ));
    LocalMux I__2398 (
            .O(N__13773),
            .I(\transmit_module.video_signal_controller.VGA_X_11 ));
    CEMux I__2397 (
            .O(N__13768),
            .I(N__13765));
    LocalMux I__2396 (
            .O(N__13765),
            .I(N__13762));
    Span4Mux_v I__2395 (
            .O(N__13762),
            .I(N__13758));
    CEMux I__2394 (
            .O(N__13761),
            .I(N__13755));
    Span4Mux_h I__2393 (
            .O(N__13758),
            .I(N__13748));
    LocalMux I__2392 (
            .O(N__13755),
            .I(N__13748));
    SRMux I__2391 (
            .O(N__13754),
            .I(N__13745));
    SRMux I__2390 (
            .O(N__13753),
            .I(N__13742));
    Span4Mux_v I__2389 (
            .O(N__13748),
            .I(N__13739));
    LocalMux I__2388 (
            .O(N__13745),
            .I(N__13736));
    LocalMux I__2387 (
            .O(N__13742),
            .I(N__13733));
    Odrv4 I__2386 (
            .O(N__13739),
            .I(\transmit_module.video_signal_controller.n2274 ));
    Odrv4 I__2385 (
            .O(N__13736),
            .I(\transmit_module.video_signal_controller.n2274 ));
    Odrv4 I__2384 (
            .O(N__13733),
            .I(\transmit_module.video_signal_controller.n2274 ));
    InMux I__2383 (
            .O(N__13726),
            .I(N__13723));
    LocalMux I__2382 (
            .O(N__13723),
            .I(N__13720));
    Odrv4 I__2381 (
            .O(N__13720),
            .I(\line_buffer.n4102 ));
    InMux I__2380 (
            .O(N__13717),
            .I(N__13714));
    LocalMux I__2379 (
            .O(N__13714),
            .I(N__13711));
    Span12Mux_v I__2378 (
            .O(N__13711),
            .I(N__13708));
    Span12Mux_h I__2377 (
            .O(N__13708),
            .I(N__13705));
    Odrv12 I__2376 (
            .O(N__13705),
            .I(\line_buffer.n648 ));
    CascadeMux I__2375 (
            .O(N__13702),
            .I(N__13699));
    InMux I__2374 (
            .O(N__13699),
            .I(N__13696));
    LocalMux I__2373 (
            .O(N__13696),
            .I(N__13693));
    Span4Mux_v I__2372 (
            .O(N__13693),
            .I(N__13690));
    Span4Mux_h I__2371 (
            .O(N__13690),
            .I(N__13687));
    Odrv4 I__2370 (
            .O(N__13687),
            .I(\line_buffer.n656 ));
    InMux I__2369 (
            .O(N__13684),
            .I(N__13678));
    InMux I__2368 (
            .O(N__13683),
            .I(N__13673));
    InMux I__2367 (
            .O(N__13682),
            .I(N__13673));
    InMux I__2366 (
            .O(N__13681),
            .I(N__13670));
    LocalMux I__2365 (
            .O(N__13678),
            .I(\transmit_module.video_signal_controller.VGA_X_1 ));
    LocalMux I__2364 (
            .O(N__13673),
            .I(\transmit_module.video_signal_controller.VGA_X_1 ));
    LocalMux I__2363 (
            .O(N__13670),
            .I(\transmit_module.video_signal_controller.VGA_X_1 ));
    InMux I__2362 (
            .O(N__13663),
            .I(\transmit_module.video_signal_controller.n3688 ));
    CascadeMux I__2361 (
            .O(N__13660),
            .I(N__13656));
    InMux I__2360 (
            .O(N__13659),
            .I(N__13651));
    InMux I__2359 (
            .O(N__13656),
            .I(N__13646));
    InMux I__2358 (
            .O(N__13655),
            .I(N__13646));
    InMux I__2357 (
            .O(N__13654),
            .I(N__13643));
    LocalMux I__2356 (
            .O(N__13651),
            .I(\transmit_module.video_signal_controller.VGA_X_2 ));
    LocalMux I__2355 (
            .O(N__13646),
            .I(\transmit_module.video_signal_controller.VGA_X_2 ));
    LocalMux I__2354 (
            .O(N__13643),
            .I(\transmit_module.video_signal_controller.VGA_X_2 ));
    InMux I__2353 (
            .O(N__13636),
            .I(\transmit_module.video_signal_controller.n3689 ));
    InMux I__2352 (
            .O(N__13633),
            .I(N__13627));
    InMux I__2351 (
            .O(N__13632),
            .I(N__13624));
    InMux I__2350 (
            .O(N__13631),
            .I(N__13621));
    InMux I__2349 (
            .O(N__13630),
            .I(N__13618));
    LocalMux I__2348 (
            .O(N__13627),
            .I(\transmit_module.video_signal_controller.VGA_X_3 ));
    LocalMux I__2347 (
            .O(N__13624),
            .I(\transmit_module.video_signal_controller.VGA_X_3 ));
    LocalMux I__2346 (
            .O(N__13621),
            .I(\transmit_module.video_signal_controller.VGA_X_3 ));
    LocalMux I__2345 (
            .O(N__13618),
            .I(\transmit_module.video_signal_controller.VGA_X_3 ));
    InMux I__2344 (
            .O(N__13609),
            .I(\transmit_module.video_signal_controller.n3690 ));
    InMux I__2343 (
            .O(N__13606),
            .I(N__13600));
    InMux I__2342 (
            .O(N__13605),
            .I(N__13593));
    InMux I__2341 (
            .O(N__13604),
            .I(N__13593));
    InMux I__2340 (
            .O(N__13603),
            .I(N__13593));
    LocalMux I__2339 (
            .O(N__13600),
            .I(\transmit_module.video_signal_controller.VGA_X_4 ));
    LocalMux I__2338 (
            .O(N__13593),
            .I(\transmit_module.video_signal_controller.VGA_X_4 ));
    InMux I__2337 (
            .O(N__13588),
            .I(\transmit_module.video_signal_controller.n3691 ));
    InMux I__2336 (
            .O(N__13585),
            .I(N__13579));
    InMux I__2335 (
            .O(N__13584),
            .I(N__13574));
    InMux I__2334 (
            .O(N__13583),
            .I(N__13574));
    InMux I__2333 (
            .O(N__13582),
            .I(N__13571));
    LocalMux I__2332 (
            .O(N__13579),
            .I(\transmit_module.video_signal_controller.VGA_X_5 ));
    LocalMux I__2331 (
            .O(N__13574),
            .I(\transmit_module.video_signal_controller.VGA_X_5 ));
    LocalMux I__2330 (
            .O(N__13571),
            .I(\transmit_module.video_signal_controller.VGA_X_5 ));
    InMux I__2329 (
            .O(N__13564),
            .I(\transmit_module.video_signal_controller.n3692 ));
    InMux I__2328 (
            .O(N__13561),
            .I(N__13555));
    InMux I__2327 (
            .O(N__13560),
            .I(N__13550));
    InMux I__2326 (
            .O(N__13559),
            .I(N__13550));
    InMux I__2325 (
            .O(N__13558),
            .I(N__13547));
    LocalMux I__2324 (
            .O(N__13555),
            .I(\transmit_module.video_signal_controller.VGA_X_6 ));
    LocalMux I__2323 (
            .O(N__13550),
            .I(\transmit_module.video_signal_controller.VGA_X_6 ));
    LocalMux I__2322 (
            .O(N__13547),
            .I(\transmit_module.video_signal_controller.VGA_X_6 ));
    InMux I__2321 (
            .O(N__13540),
            .I(\transmit_module.video_signal_controller.n3693 ));
    InMux I__2320 (
            .O(N__13537),
            .I(N__13529));
    InMux I__2319 (
            .O(N__13536),
            .I(N__13529));
    InMux I__2318 (
            .O(N__13535),
            .I(N__13526));
    InMux I__2317 (
            .O(N__13534),
            .I(N__13523));
    LocalMux I__2316 (
            .O(N__13529),
            .I(\transmit_module.video_signal_controller.VGA_X_7 ));
    LocalMux I__2315 (
            .O(N__13526),
            .I(\transmit_module.video_signal_controller.VGA_X_7 ));
    LocalMux I__2314 (
            .O(N__13523),
            .I(\transmit_module.video_signal_controller.VGA_X_7 ));
    InMux I__2313 (
            .O(N__13516),
            .I(\transmit_module.video_signal_controller.n3694 ));
    InMux I__2312 (
            .O(N__13513),
            .I(N__13510));
    LocalMux I__2311 (
            .O(N__13510),
            .I(N__13504));
    InMux I__2310 (
            .O(N__13509),
            .I(N__13501));
    InMux I__2309 (
            .O(N__13508),
            .I(N__13496));
    InMux I__2308 (
            .O(N__13507),
            .I(N__13496));
    Odrv4 I__2307 (
            .O(N__13504),
            .I(\transmit_module.video_signal_controller.VGA_X_8 ));
    LocalMux I__2306 (
            .O(N__13501),
            .I(\transmit_module.video_signal_controller.VGA_X_8 ));
    LocalMux I__2305 (
            .O(N__13496),
            .I(\transmit_module.video_signal_controller.VGA_X_8 ));
    InMux I__2304 (
            .O(N__13489),
            .I(bfn_13_16_0_));
    SRMux I__2303 (
            .O(N__13486),
            .I(N__13482));
    SRMux I__2302 (
            .O(N__13485),
            .I(N__13479));
    LocalMux I__2301 (
            .O(N__13482),
            .I(N__13476));
    LocalMux I__2300 (
            .O(N__13479),
            .I(N__13471));
    Span4Mux_v I__2299 (
            .O(N__13476),
            .I(N__13468));
    SRMux I__2298 (
            .O(N__13475),
            .I(N__13465));
    SRMux I__2297 (
            .O(N__13474),
            .I(N__13462));
    Span12Mux_s2_v I__2296 (
            .O(N__13471),
            .I(N__13455));
    Sp12to4 I__2295 (
            .O(N__13468),
            .I(N__13455));
    LocalMux I__2294 (
            .O(N__13465),
            .I(N__13455));
    LocalMux I__2293 (
            .O(N__13462),
            .I(N__13452));
    Span12Mux_v I__2292 (
            .O(N__13455),
            .I(N__13449));
    Span4Mux_v I__2291 (
            .O(N__13452),
            .I(N__13446));
    Span12Mux_h I__2290 (
            .O(N__13449),
            .I(N__13443));
    Span4Mux_h I__2289 (
            .O(N__13446),
            .I(N__13440));
    Odrv12 I__2288 (
            .O(N__13443),
            .I(n690));
    Odrv4 I__2287 (
            .O(N__13440),
            .I(n690));
    CascadeMux I__2286 (
            .O(N__13435),
            .I(N__13432));
    InMux I__2285 (
            .O(N__13432),
            .I(N__13429));
    LocalMux I__2284 (
            .O(N__13429),
            .I(\db5.COUNTER_3 ));
    InMux I__2283 (
            .O(N__13426),
            .I(N__13419));
    InMux I__2282 (
            .O(N__13425),
            .I(N__13419));
    InMux I__2281 (
            .O(N__13424),
            .I(N__13416));
    LocalMux I__2280 (
            .O(N__13419),
            .I(N__13413));
    LocalMux I__2279 (
            .O(N__13416),
            .I(\db5.NEXT_COUNTER_3 ));
    Odrv4 I__2278 (
            .O(N__13413),
            .I(\db5.NEXT_COUNTER_3 ));
    InMux I__2277 (
            .O(N__13408),
            .I(N__13404));
    InMux I__2276 (
            .O(N__13407),
            .I(N__13401));
    LocalMux I__2275 (
            .O(N__13404),
            .I(N__13396));
    LocalMux I__2274 (
            .O(N__13401),
            .I(N__13396));
    Odrv4 I__2273 (
            .O(N__13396),
            .I(\db5.COUNTER_2 ));
    CascadeMux I__2272 (
            .O(N__13393),
            .I(N__13390));
    InMux I__2271 (
            .O(N__13390),
            .I(N__13381));
    InMux I__2270 (
            .O(N__13389),
            .I(N__13381));
    InMux I__2269 (
            .O(N__13388),
            .I(N__13381));
    LocalMux I__2268 (
            .O(N__13381),
            .I(N__13378));
    Odrv4 I__2267 (
            .O(N__13378),
            .I(\db5.NEXT_COUNTER_2 ));
    InMux I__2266 (
            .O(N__13375),
            .I(N__13366));
    InMux I__2265 (
            .O(N__13374),
            .I(N__13366));
    InMux I__2264 (
            .O(N__13373),
            .I(N__13366));
    LocalMux I__2263 (
            .O(N__13366),
            .I(\db5.COUNTER_1 ));
    CascadeMux I__2262 (
            .O(N__13363),
            .I(N__13360));
    InMux I__2261 (
            .O(N__13360),
            .I(N__13357));
    LocalMux I__2260 (
            .O(N__13357),
            .I(N__13353));
    InMux I__2259 (
            .O(N__13356),
            .I(N__13350));
    Odrv4 I__2258 (
            .O(N__13353),
            .I(\db5.NEXT_COUNTER_1 ));
    LocalMux I__2257 (
            .O(N__13350),
            .I(\db5.NEXT_COUNTER_1 ));
    InMux I__2256 (
            .O(N__13345),
            .I(N__13333));
    InMux I__2255 (
            .O(N__13344),
            .I(N__13333));
    InMux I__2254 (
            .O(N__13343),
            .I(N__13333));
    InMux I__2253 (
            .O(N__13342),
            .I(N__13333));
    LocalMux I__2252 (
            .O(N__13333),
            .I(N__13330));
    Odrv4 I__2251 (
            .O(N__13330),
            .I(\db5.COUNTER_0 ));
    InMux I__2250 (
            .O(N__13327),
            .I(N__13321));
    InMux I__2249 (
            .O(N__13326),
            .I(N__13321));
    LocalMux I__2248 (
            .O(N__13321),
            .I(N__13318));
    Odrv4 I__2247 (
            .O(N__13318),
            .I(\db5.NEXT_COUNTER_0 ));
    SRMux I__2246 (
            .O(N__13315),
            .I(N__13312));
    LocalMux I__2245 (
            .O(N__13312),
            .I(N__13309));
    Span4Mux_v I__2244 (
            .O(N__13309),
            .I(N__13306));
    Odrv4 I__2243 (
            .O(N__13306),
            .I(\db5.n4221 ));
    CascadeMux I__2242 (
            .O(N__13303),
            .I(N__13300));
    InMux I__2241 (
            .O(N__13300),
            .I(N__13297));
    LocalMux I__2240 (
            .O(N__13297),
            .I(\transmit_module.video_signal_controller.n3997 ));
    InMux I__2239 (
            .O(N__13294),
            .I(N__13291));
    LocalMux I__2238 (
            .O(N__13291),
            .I(\transmit_module.video_signal_controller.n3196 ));
    InMux I__2237 (
            .O(N__13288),
            .I(N__13285));
    LocalMux I__2236 (
            .O(N__13285),
            .I(N__13282));
    Span4Mux_v I__2235 (
            .O(N__13282),
            .I(N__13279));
    Span4Mux_v I__2234 (
            .O(N__13279),
            .I(N__13276));
    Span4Mux_h I__2233 (
            .O(N__13276),
            .I(N__13273));
    Odrv4 I__2232 (
            .O(N__13273),
            .I(\line_buffer.n655 ));
    InMux I__2231 (
            .O(N__13270),
            .I(N__13267));
    LocalMux I__2230 (
            .O(N__13267),
            .I(N__13264));
    Span12Mux_v I__2229 (
            .O(N__13264),
            .I(N__13261));
    Span12Mux_h I__2228 (
            .O(N__13261),
            .I(N__13258));
    Odrv12 I__2227 (
            .O(N__13258),
            .I(\line_buffer.n647 ));
    InMux I__2226 (
            .O(N__13255),
            .I(N__13250));
    InMux I__2225 (
            .O(N__13254),
            .I(N__13245));
    InMux I__2224 (
            .O(N__13253),
            .I(N__13245));
    LocalMux I__2223 (
            .O(N__13250),
            .I(\transmit_module.video_signal_controller.VGA_X_0 ));
    LocalMux I__2222 (
            .O(N__13245),
            .I(\transmit_module.video_signal_controller.VGA_X_0 ));
    InMux I__2221 (
            .O(N__13240),
            .I(bfn_13_15_0_));
    InMux I__2220 (
            .O(N__13237),
            .I(N__13234));
    LocalMux I__2219 (
            .O(N__13234),
            .I(\receive_module.n7 ));
    CascadeMux I__2218 (
            .O(N__13231),
            .I(N__13228));
    InMux I__2217 (
            .O(N__13228),
            .I(N__13225));
    LocalMux I__2216 (
            .O(N__13225),
            .I(N__13222));
    Span4Mux_v I__2215 (
            .O(N__13222),
            .I(N__13217));
    InMux I__2214 (
            .O(N__13221),
            .I(N__13212));
    InMux I__2213 (
            .O(N__13220),
            .I(N__13212));
    Odrv4 I__2212 (
            .O(N__13217),
            .I(\receive_module.O_Y_3 ));
    LocalMux I__2211 (
            .O(N__13212),
            .I(\receive_module.O_Y_3 ));
    CascadeMux I__2210 (
            .O(N__13207),
            .I(N__13203));
    CascadeMux I__2209 (
            .O(N__13206),
            .I(N__13200));
    CascadeBuf I__2208 (
            .O(N__13203),
            .I(N__13197));
    CascadeBuf I__2207 (
            .O(N__13200),
            .I(N__13194));
    CascadeMux I__2206 (
            .O(N__13197),
            .I(N__13191));
    CascadeMux I__2205 (
            .O(N__13194),
            .I(N__13188));
    CascadeBuf I__2204 (
            .O(N__13191),
            .I(N__13185));
    CascadeBuf I__2203 (
            .O(N__13188),
            .I(N__13182));
    CascadeMux I__2202 (
            .O(N__13185),
            .I(N__13179));
    CascadeMux I__2201 (
            .O(N__13182),
            .I(N__13176));
    CascadeBuf I__2200 (
            .O(N__13179),
            .I(N__13173));
    CascadeBuf I__2199 (
            .O(N__13176),
            .I(N__13170));
    CascadeMux I__2198 (
            .O(N__13173),
            .I(N__13167));
    CascadeMux I__2197 (
            .O(N__13170),
            .I(N__13164));
    CascadeBuf I__2196 (
            .O(N__13167),
            .I(N__13161));
    CascadeBuf I__2195 (
            .O(N__13164),
            .I(N__13158));
    CascadeMux I__2194 (
            .O(N__13161),
            .I(N__13155));
    CascadeMux I__2193 (
            .O(N__13158),
            .I(N__13152));
    CascadeBuf I__2192 (
            .O(N__13155),
            .I(N__13149));
    CascadeBuf I__2191 (
            .O(N__13152),
            .I(N__13146));
    CascadeMux I__2190 (
            .O(N__13149),
            .I(N__13143));
    CascadeMux I__2189 (
            .O(N__13146),
            .I(N__13140));
    CascadeBuf I__2188 (
            .O(N__13143),
            .I(N__13137));
    CascadeBuf I__2187 (
            .O(N__13140),
            .I(N__13134));
    CascadeMux I__2186 (
            .O(N__13137),
            .I(N__13131));
    CascadeMux I__2185 (
            .O(N__13134),
            .I(N__13128));
    CascadeBuf I__2184 (
            .O(N__13131),
            .I(N__13125));
    CascadeBuf I__2183 (
            .O(N__13128),
            .I(N__13122));
    CascadeMux I__2182 (
            .O(N__13125),
            .I(N__13119));
    CascadeMux I__2181 (
            .O(N__13122),
            .I(N__13116));
    CascadeBuf I__2180 (
            .O(N__13119),
            .I(N__13113));
    CascadeBuf I__2179 (
            .O(N__13116),
            .I(N__13110));
    CascadeMux I__2178 (
            .O(N__13113),
            .I(N__13107));
    CascadeMux I__2177 (
            .O(N__13110),
            .I(N__13104));
    CascadeBuf I__2176 (
            .O(N__13107),
            .I(N__13101));
    CascadeBuf I__2175 (
            .O(N__13104),
            .I(N__13098));
    CascadeMux I__2174 (
            .O(N__13101),
            .I(N__13095));
    CascadeMux I__2173 (
            .O(N__13098),
            .I(N__13092));
    CascadeBuf I__2172 (
            .O(N__13095),
            .I(N__13089));
    CascadeBuf I__2171 (
            .O(N__13092),
            .I(N__13086));
    CascadeMux I__2170 (
            .O(N__13089),
            .I(N__13083));
    CascadeMux I__2169 (
            .O(N__13086),
            .I(N__13080));
    CascadeBuf I__2168 (
            .O(N__13083),
            .I(N__13077));
    CascadeBuf I__2167 (
            .O(N__13080),
            .I(N__13074));
    CascadeMux I__2166 (
            .O(N__13077),
            .I(N__13071));
    CascadeMux I__2165 (
            .O(N__13074),
            .I(N__13068));
    CascadeBuf I__2164 (
            .O(N__13071),
            .I(N__13065));
    CascadeBuf I__2163 (
            .O(N__13068),
            .I(N__13062));
    CascadeMux I__2162 (
            .O(N__13065),
            .I(N__13059));
    CascadeMux I__2161 (
            .O(N__13062),
            .I(N__13056));
    CascadeBuf I__2160 (
            .O(N__13059),
            .I(N__13053));
    CascadeBuf I__2159 (
            .O(N__13056),
            .I(N__13050));
    CascadeMux I__2158 (
            .O(N__13053),
            .I(N__13047));
    CascadeMux I__2157 (
            .O(N__13050),
            .I(N__13044));
    CascadeBuf I__2156 (
            .O(N__13047),
            .I(N__13041));
    CascadeBuf I__2155 (
            .O(N__13044),
            .I(N__13038));
    CascadeMux I__2154 (
            .O(N__13041),
            .I(N__13035));
    CascadeMux I__2153 (
            .O(N__13038),
            .I(N__13032));
    CascadeBuf I__2152 (
            .O(N__13035),
            .I(N__13029));
    CascadeBuf I__2151 (
            .O(N__13032),
            .I(N__13026));
    CascadeMux I__2150 (
            .O(N__13029),
            .I(N__13023));
    CascadeMux I__2149 (
            .O(N__13026),
            .I(N__13020));
    InMux I__2148 (
            .O(N__13023),
            .I(N__13017));
    InMux I__2147 (
            .O(N__13020),
            .I(N__13014));
    LocalMux I__2146 (
            .O(N__13017),
            .I(N__13011));
    LocalMux I__2145 (
            .O(N__13014),
            .I(N__13008));
    Span4Mux_h I__2144 (
            .O(N__13011),
            .I(N__13005));
    Span12Mux_s6_v I__2143 (
            .O(N__13008),
            .I(N__13002));
    Sp12to4 I__2142 (
            .O(N__13005),
            .I(N__12999));
    Span12Mux_v I__2141 (
            .O(N__13002),
            .I(N__12996));
    Span12Mux_s9_v I__2140 (
            .O(N__12999),
            .I(N__12993));
    Span12Mux_h I__2139 (
            .O(N__12996),
            .I(N__12990));
    Span12Mux_v I__2138 (
            .O(N__12993),
            .I(N__12987));
    Odrv12 I__2137 (
            .O(N__12990),
            .I(RX_ADDR_9));
    Odrv12 I__2136 (
            .O(N__12987),
            .I(RX_ADDR_9));
    InMux I__2135 (
            .O(N__12982),
            .I(\receive_module.n3701 ));
    InMux I__2134 (
            .O(N__12979),
            .I(N__12976));
    LocalMux I__2133 (
            .O(N__12976),
            .I(\receive_module.n6 ));
    CascadeMux I__2132 (
            .O(N__12973),
            .I(N__12970));
    InMux I__2131 (
            .O(N__12970),
            .I(N__12967));
    LocalMux I__2130 (
            .O(N__12967),
            .I(N__12964));
    Span4Mux_h I__2129 (
            .O(N__12964),
            .I(N__12960));
    InMux I__2128 (
            .O(N__12963),
            .I(N__12957));
    Odrv4 I__2127 (
            .O(N__12960),
            .I(\receive_module.O_Y_4 ));
    LocalMux I__2126 (
            .O(N__12957),
            .I(\receive_module.O_Y_4 ));
    CascadeMux I__2125 (
            .O(N__12952),
            .I(N__12949));
    CascadeBuf I__2124 (
            .O(N__12949),
            .I(N__12945));
    CascadeMux I__2123 (
            .O(N__12948),
            .I(N__12942));
    CascadeMux I__2122 (
            .O(N__12945),
            .I(N__12939));
    CascadeBuf I__2121 (
            .O(N__12942),
            .I(N__12936));
    CascadeBuf I__2120 (
            .O(N__12939),
            .I(N__12933));
    CascadeMux I__2119 (
            .O(N__12936),
            .I(N__12930));
    CascadeMux I__2118 (
            .O(N__12933),
            .I(N__12927));
    CascadeBuf I__2117 (
            .O(N__12930),
            .I(N__12924));
    CascadeBuf I__2116 (
            .O(N__12927),
            .I(N__12921));
    CascadeMux I__2115 (
            .O(N__12924),
            .I(N__12918));
    CascadeMux I__2114 (
            .O(N__12921),
            .I(N__12915));
    CascadeBuf I__2113 (
            .O(N__12918),
            .I(N__12912));
    CascadeBuf I__2112 (
            .O(N__12915),
            .I(N__12909));
    CascadeMux I__2111 (
            .O(N__12912),
            .I(N__12906));
    CascadeMux I__2110 (
            .O(N__12909),
            .I(N__12903));
    CascadeBuf I__2109 (
            .O(N__12906),
            .I(N__12900));
    CascadeBuf I__2108 (
            .O(N__12903),
            .I(N__12897));
    CascadeMux I__2107 (
            .O(N__12900),
            .I(N__12894));
    CascadeMux I__2106 (
            .O(N__12897),
            .I(N__12891));
    CascadeBuf I__2105 (
            .O(N__12894),
            .I(N__12888));
    CascadeBuf I__2104 (
            .O(N__12891),
            .I(N__12885));
    CascadeMux I__2103 (
            .O(N__12888),
            .I(N__12882));
    CascadeMux I__2102 (
            .O(N__12885),
            .I(N__12879));
    CascadeBuf I__2101 (
            .O(N__12882),
            .I(N__12876));
    CascadeBuf I__2100 (
            .O(N__12879),
            .I(N__12873));
    CascadeMux I__2099 (
            .O(N__12876),
            .I(N__12870));
    CascadeMux I__2098 (
            .O(N__12873),
            .I(N__12867));
    CascadeBuf I__2097 (
            .O(N__12870),
            .I(N__12864));
    CascadeBuf I__2096 (
            .O(N__12867),
            .I(N__12861));
    CascadeMux I__2095 (
            .O(N__12864),
            .I(N__12858));
    CascadeMux I__2094 (
            .O(N__12861),
            .I(N__12855));
    CascadeBuf I__2093 (
            .O(N__12858),
            .I(N__12852));
    CascadeBuf I__2092 (
            .O(N__12855),
            .I(N__12849));
    CascadeMux I__2091 (
            .O(N__12852),
            .I(N__12846));
    CascadeMux I__2090 (
            .O(N__12849),
            .I(N__12843));
    CascadeBuf I__2089 (
            .O(N__12846),
            .I(N__12840));
    CascadeBuf I__2088 (
            .O(N__12843),
            .I(N__12837));
    CascadeMux I__2087 (
            .O(N__12840),
            .I(N__12834));
    CascadeMux I__2086 (
            .O(N__12837),
            .I(N__12831));
    CascadeBuf I__2085 (
            .O(N__12834),
            .I(N__12828));
    CascadeBuf I__2084 (
            .O(N__12831),
            .I(N__12825));
    CascadeMux I__2083 (
            .O(N__12828),
            .I(N__12822));
    CascadeMux I__2082 (
            .O(N__12825),
            .I(N__12819));
    CascadeBuf I__2081 (
            .O(N__12822),
            .I(N__12816));
    CascadeBuf I__2080 (
            .O(N__12819),
            .I(N__12813));
    CascadeMux I__2079 (
            .O(N__12816),
            .I(N__12810));
    CascadeMux I__2078 (
            .O(N__12813),
            .I(N__12807));
    CascadeBuf I__2077 (
            .O(N__12810),
            .I(N__12804));
    CascadeBuf I__2076 (
            .O(N__12807),
            .I(N__12801));
    CascadeMux I__2075 (
            .O(N__12804),
            .I(N__12798));
    CascadeMux I__2074 (
            .O(N__12801),
            .I(N__12795));
    CascadeBuf I__2073 (
            .O(N__12798),
            .I(N__12792));
    CascadeBuf I__2072 (
            .O(N__12795),
            .I(N__12789));
    CascadeMux I__2071 (
            .O(N__12792),
            .I(N__12786));
    CascadeMux I__2070 (
            .O(N__12789),
            .I(N__12783));
    CascadeBuf I__2069 (
            .O(N__12786),
            .I(N__12780));
    CascadeBuf I__2068 (
            .O(N__12783),
            .I(N__12777));
    CascadeMux I__2067 (
            .O(N__12780),
            .I(N__12774));
    CascadeMux I__2066 (
            .O(N__12777),
            .I(N__12771));
    CascadeBuf I__2065 (
            .O(N__12774),
            .I(N__12768));
    InMux I__2064 (
            .O(N__12771),
            .I(N__12765));
    CascadeMux I__2063 (
            .O(N__12768),
            .I(N__12762));
    LocalMux I__2062 (
            .O(N__12765),
            .I(N__12759));
    InMux I__2061 (
            .O(N__12762),
            .I(N__12756));
    Span4Mux_s1_v I__2060 (
            .O(N__12759),
            .I(N__12753));
    LocalMux I__2059 (
            .O(N__12756),
            .I(N__12750));
    Span4Mux_h I__2058 (
            .O(N__12753),
            .I(N__12747));
    Span12Mux_s5_v I__2057 (
            .O(N__12750),
            .I(N__12744));
    Span4Mux_v I__2056 (
            .O(N__12747),
            .I(N__12741));
    Span12Mux_h I__2055 (
            .O(N__12744),
            .I(N__12736));
    Sp12to4 I__2054 (
            .O(N__12741),
            .I(N__12736));
    Span12Mux_v I__2053 (
            .O(N__12736),
            .I(N__12733));
    Odrv12 I__2052 (
            .O(N__12733),
            .I(RX_ADDR_10));
    InMux I__2051 (
            .O(N__12730),
            .I(\receive_module.n3702 ));
    InMux I__2050 (
            .O(N__12727),
            .I(N__12724));
    LocalMux I__2049 (
            .O(N__12724),
            .I(\receive_module.n5 ));
    CascadeMux I__2048 (
            .O(N__12721),
            .I(N__12718));
    InMux I__2047 (
            .O(N__12718),
            .I(N__12715));
    LocalMux I__2046 (
            .O(N__12715),
            .I(N__12712));
    Span4Mux_h I__2045 (
            .O(N__12712),
            .I(N__12709));
    Odrv4 I__2044 (
            .O(N__12709),
            .I(\receive_module.O_Y_5 ));
    InMux I__2043 (
            .O(N__12706),
            .I(\receive_module.n3703 ));
    InMux I__2042 (
            .O(N__12703),
            .I(N__12700));
    LocalMux I__2041 (
            .O(N__12700),
            .I(\receive_module.n4 ));
    CascadeMux I__2040 (
            .O(N__12697),
            .I(N__12694));
    InMux I__2039 (
            .O(N__12694),
            .I(N__12691));
    LocalMux I__2038 (
            .O(N__12691),
            .I(N__12688));
    Span4Mux_h I__2037 (
            .O(N__12688),
            .I(N__12685));
    Odrv4 I__2036 (
            .O(N__12685),
            .I(\receive_module.O_Y_6 ));
    InMux I__2035 (
            .O(N__12682),
            .I(\receive_module.n3704 ));
    InMux I__2034 (
            .O(N__12679),
            .I(N__12676));
    LocalMux I__2033 (
            .O(N__12676),
            .I(\receive_module.n3 ));
    InMux I__2032 (
            .O(N__12673),
            .I(N__12670));
    LocalMux I__2031 (
            .O(N__12670),
            .I(N__12667));
    Span4Mux_v I__2030 (
            .O(N__12667),
            .I(N__12664));
    Odrv4 I__2029 (
            .O(N__12664),
            .I(\receive_module.O_Y_7 ));
    InMux I__2028 (
            .O(N__12661),
            .I(\receive_module.n3705 ));
    SRMux I__2027 (
            .O(N__12658),
            .I(N__12653));
    SRMux I__2026 (
            .O(N__12657),
            .I(N__12650));
    SRMux I__2025 (
            .O(N__12656),
            .I(N__12647));
    LocalMux I__2024 (
            .O(N__12653),
            .I(N__12643));
    LocalMux I__2023 (
            .O(N__12650),
            .I(N__12638));
    LocalMux I__2022 (
            .O(N__12647),
            .I(N__12638));
    SRMux I__2021 (
            .O(N__12646),
            .I(N__12635));
    Span4Mux_v I__2020 (
            .O(N__12643),
            .I(N__12632));
    Span4Mux_s3_v I__2019 (
            .O(N__12638),
            .I(N__12627));
    LocalMux I__2018 (
            .O(N__12635),
            .I(N__12627));
    Span4Mux_h I__2017 (
            .O(N__12632),
            .I(N__12624));
    Span4Mux_v I__2016 (
            .O(N__12627),
            .I(N__12621));
    Span4Mux_v I__2015 (
            .O(N__12624),
            .I(N__12618));
    Span4Mux_h I__2014 (
            .O(N__12621),
            .I(N__12615));
    Odrv4 I__2013 (
            .O(N__12618),
            .I(\line_buffer.n627 ));
    Odrv4 I__2012 (
            .O(N__12615),
            .I(\line_buffer.n627 ));
    SRMux I__2011 (
            .O(N__12610),
            .I(N__12607));
    LocalMux I__2010 (
            .O(N__12607),
            .I(N__12602));
    SRMux I__2009 (
            .O(N__12606),
            .I(N__12599));
    SRMux I__2008 (
            .O(N__12605),
            .I(N__12595));
    Span4Mux_h I__2007 (
            .O(N__12602),
            .I(N__12592));
    LocalMux I__2006 (
            .O(N__12599),
            .I(N__12589));
    SRMux I__2005 (
            .O(N__12598),
            .I(N__12586));
    LocalMux I__2004 (
            .O(N__12595),
            .I(N__12583));
    Span4Mux_v I__2003 (
            .O(N__12592),
            .I(N__12578));
    Span4Mux_h I__2002 (
            .O(N__12589),
            .I(N__12578));
    LocalMux I__2001 (
            .O(N__12586),
            .I(N__12575));
    Span12Mux_s10_v I__2000 (
            .O(N__12583),
            .I(N__12570));
    Sp12to4 I__1999 (
            .O(N__12578),
            .I(N__12570));
    Span12Mux_v I__1998 (
            .O(N__12575),
            .I(N__12567));
    Span12Mux_h I__1997 (
            .O(N__12570),
            .I(N__12562));
    Span12Mux_h I__1996 (
            .O(N__12567),
            .I(N__12562));
    Odrv12 I__1995 (
            .O(N__12562),
            .I(\line_buffer.n562 ));
    InMux I__1994 (
            .O(N__12559),
            .I(\receive_module.rx_counter.n3652 ));
    InMux I__1993 (
            .O(N__12556),
            .I(\receive_module.rx_counter.n3653 ));
    InMux I__1992 (
            .O(N__12553),
            .I(\receive_module.rx_counter.n3654 ));
    InMux I__1991 (
            .O(N__12550),
            .I(\receive_module.rx_counter.n3655 ));
    InMux I__1990 (
            .O(N__12547),
            .I(N__12532));
    InMux I__1989 (
            .O(N__12546),
            .I(N__12532));
    InMux I__1988 (
            .O(N__12545),
            .I(N__12532));
    InMux I__1987 (
            .O(N__12544),
            .I(N__12532));
    InMux I__1986 (
            .O(N__12543),
            .I(N__12532));
    LocalMux I__1985 (
            .O(N__12532),
            .I(\receive_module.O_X_9 ));
    CascadeMux I__1984 (
            .O(N__12529),
            .I(N__12526));
    InMux I__1983 (
            .O(N__12526),
            .I(N__12523));
    LocalMux I__1982 (
            .O(N__12523),
            .I(\receive_module.rx_counter.n4 ));
    InMux I__1981 (
            .O(N__12520),
            .I(N__12517));
    LocalMux I__1980 (
            .O(N__12517),
            .I(N__12513));
    CascadeMux I__1979 (
            .O(N__12516),
            .I(N__12509));
    Span4Mux_h I__1978 (
            .O(N__12513),
            .I(N__12503));
    InMux I__1977 (
            .O(N__12512),
            .I(N__12500));
    InMux I__1976 (
            .O(N__12509),
            .I(N__12491));
    InMux I__1975 (
            .O(N__12508),
            .I(N__12491));
    InMux I__1974 (
            .O(N__12507),
            .I(N__12491));
    InMux I__1973 (
            .O(N__12506),
            .I(N__12491));
    Odrv4 I__1972 (
            .O(N__12503),
            .I(\receive_module.O_Y_0 ));
    LocalMux I__1971 (
            .O(N__12500),
            .I(\receive_module.O_Y_0 ));
    LocalMux I__1970 (
            .O(N__12491),
            .I(\receive_module.O_Y_0 ));
    CascadeMux I__1969 (
            .O(N__12484),
            .I(N__12481));
    InMux I__1968 (
            .O(N__12481),
            .I(N__12478));
    LocalMux I__1967 (
            .O(N__12478),
            .I(\receive_module.O_X_6 ));
    CascadeMux I__1966 (
            .O(N__12475),
            .I(N__12472));
    CascadeBuf I__1965 (
            .O(N__12472),
            .I(N__12469));
    CascadeMux I__1964 (
            .O(N__12469),
            .I(N__12465));
    CascadeMux I__1963 (
            .O(N__12468),
            .I(N__12462));
    CascadeBuf I__1962 (
            .O(N__12465),
            .I(N__12459));
    CascadeBuf I__1961 (
            .O(N__12462),
            .I(N__12456));
    CascadeMux I__1960 (
            .O(N__12459),
            .I(N__12453));
    CascadeMux I__1959 (
            .O(N__12456),
            .I(N__12450));
    CascadeBuf I__1958 (
            .O(N__12453),
            .I(N__12447));
    CascadeBuf I__1957 (
            .O(N__12450),
            .I(N__12444));
    CascadeMux I__1956 (
            .O(N__12447),
            .I(N__12441));
    CascadeMux I__1955 (
            .O(N__12444),
            .I(N__12438));
    CascadeBuf I__1954 (
            .O(N__12441),
            .I(N__12435));
    CascadeBuf I__1953 (
            .O(N__12438),
            .I(N__12432));
    CascadeMux I__1952 (
            .O(N__12435),
            .I(N__12429));
    CascadeMux I__1951 (
            .O(N__12432),
            .I(N__12426));
    CascadeBuf I__1950 (
            .O(N__12429),
            .I(N__12423));
    CascadeBuf I__1949 (
            .O(N__12426),
            .I(N__12420));
    CascadeMux I__1948 (
            .O(N__12423),
            .I(N__12417));
    CascadeMux I__1947 (
            .O(N__12420),
            .I(N__12414));
    CascadeBuf I__1946 (
            .O(N__12417),
            .I(N__12411));
    CascadeBuf I__1945 (
            .O(N__12414),
            .I(N__12408));
    CascadeMux I__1944 (
            .O(N__12411),
            .I(N__12405));
    CascadeMux I__1943 (
            .O(N__12408),
            .I(N__12402));
    CascadeBuf I__1942 (
            .O(N__12405),
            .I(N__12399));
    CascadeBuf I__1941 (
            .O(N__12402),
            .I(N__12396));
    CascadeMux I__1940 (
            .O(N__12399),
            .I(N__12393));
    CascadeMux I__1939 (
            .O(N__12396),
            .I(N__12390));
    CascadeBuf I__1938 (
            .O(N__12393),
            .I(N__12387));
    CascadeBuf I__1937 (
            .O(N__12390),
            .I(N__12384));
    CascadeMux I__1936 (
            .O(N__12387),
            .I(N__12381));
    CascadeMux I__1935 (
            .O(N__12384),
            .I(N__12378));
    CascadeBuf I__1934 (
            .O(N__12381),
            .I(N__12375));
    CascadeBuf I__1933 (
            .O(N__12378),
            .I(N__12372));
    CascadeMux I__1932 (
            .O(N__12375),
            .I(N__12369));
    CascadeMux I__1931 (
            .O(N__12372),
            .I(N__12366));
    CascadeBuf I__1930 (
            .O(N__12369),
            .I(N__12363));
    CascadeBuf I__1929 (
            .O(N__12366),
            .I(N__12360));
    CascadeMux I__1928 (
            .O(N__12363),
            .I(N__12357));
    CascadeMux I__1927 (
            .O(N__12360),
            .I(N__12354));
    CascadeBuf I__1926 (
            .O(N__12357),
            .I(N__12351));
    CascadeBuf I__1925 (
            .O(N__12354),
            .I(N__12348));
    CascadeMux I__1924 (
            .O(N__12351),
            .I(N__12345));
    CascadeMux I__1923 (
            .O(N__12348),
            .I(N__12342));
    CascadeBuf I__1922 (
            .O(N__12345),
            .I(N__12339));
    CascadeBuf I__1921 (
            .O(N__12342),
            .I(N__12336));
    CascadeMux I__1920 (
            .O(N__12339),
            .I(N__12333));
    CascadeMux I__1919 (
            .O(N__12336),
            .I(N__12330));
    CascadeBuf I__1918 (
            .O(N__12333),
            .I(N__12327));
    CascadeBuf I__1917 (
            .O(N__12330),
            .I(N__12324));
    CascadeMux I__1916 (
            .O(N__12327),
            .I(N__12321));
    CascadeMux I__1915 (
            .O(N__12324),
            .I(N__12318));
    CascadeBuf I__1914 (
            .O(N__12321),
            .I(N__12315));
    CascadeBuf I__1913 (
            .O(N__12318),
            .I(N__12312));
    CascadeMux I__1912 (
            .O(N__12315),
            .I(N__12309));
    CascadeMux I__1911 (
            .O(N__12312),
            .I(N__12306));
    CascadeBuf I__1910 (
            .O(N__12309),
            .I(N__12303));
    CascadeBuf I__1909 (
            .O(N__12306),
            .I(N__12300));
    CascadeMux I__1908 (
            .O(N__12303),
            .I(N__12297));
    CascadeMux I__1907 (
            .O(N__12300),
            .I(N__12294));
    InMux I__1906 (
            .O(N__12297),
            .I(N__12291));
    CascadeBuf I__1905 (
            .O(N__12294),
            .I(N__12288));
    LocalMux I__1904 (
            .O(N__12291),
            .I(N__12285));
    CascadeMux I__1903 (
            .O(N__12288),
            .I(N__12282));
    Span4Mux_s1_v I__1902 (
            .O(N__12285),
            .I(N__12279));
    InMux I__1901 (
            .O(N__12282),
            .I(N__12276));
    Span4Mux_h I__1900 (
            .O(N__12279),
            .I(N__12273));
    LocalMux I__1899 (
            .O(N__12276),
            .I(N__12270));
    Sp12to4 I__1898 (
            .O(N__12273),
            .I(N__12267));
    Sp12to4 I__1897 (
            .O(N__12270),
            .I(N__12264));
    Span12Mux_s9_v I__1896 (
            .O(N__12267),
            .I(N__12261));
    Span12Mux_s9_v I__1895 (
            .O(N__12264),
            .I(N__12258));
    Span12Mux_v I__1894 (
            .O(N__12261),
            .I(N__12253));
    Span12Mux_v I__1893 (
            .O(N__12258),
            .I(N__12253));
    Odrv12 I__1892 (
            .O(N__12253),
            .I(RX_ADDR_6));
    InMux I__1891 (
            .O(N__12250),
            .I(N__12247));
    LocalMux I__1890 (
            .O(N__12247),
            .I(\receive_module.O_X_7 ));
    CascadeMux I__1889 (
            .O(N__12244),
            .I(N__12241));
    InMux I__1888 (
            .O(N__12241),
            .I(N__12238));
    LocalMux I__1887 (
            .O(N__12238),
            .I(N__12231));
    InMux I__1886 (
            .O(N__12237),
            .I(N__12222));
    InMux I__1885 (
            .O(N__12236),
            .I(N__12222));
    InMux I__1884 (
            .O(N__12235),
            .I(N__12222));
    InMux I__1883 (
            .O(N__12234),
            .I(N__12222));
    Span4Mux_h I__1882 (
            .O(N__12231),
            .I(N__12219));
    LocalMux I__1881 (
            .O(N__12222),
            .I(\receive_module.O_Y_1 ));
    Odrv4 I__1880 (
            .O(N__12219),
            .I(\receive_module.O_Y_1 ));
    CascadeMux I__1879 (
            .O(N__12214),
            .I(N__12210));
    CascadeMux I__1878 (
            .O(N__12213),
            .I(N__12207));
    CascadeBuf I__1877 (
            .O(N__12210),
            .I(N__12204));
    CascadeBuf I__1876 (
            .O(N__12207),
            .I(N__12201));
    CascadeMux I__1875 (
            .O(N__12204),
            .I(N__12198));
    CascadeMux I__1874 (
            .O(N__12201),
            .I(N__12195));
    CascadeBuf I__1873 (
            .O(N__12198),
            .I(N__12192));
    CascadeBuf I__1872 (
            .O(N__12195),
            .I(N__12189));
    CascadeMux I__1871 (
            .O(N__12192),
            .I(N__12186));
    CascadeMux I__1870 (
            .O(N__12189),
            .I(N__12183));
    CascadeBuf I__1869 (
            .O(N__12186),
            .I(N__12180));
    CascadeBuf I__1868 (
            .O(N__12183),
            .I(N__12177));
    CascadeMux I__1867 (
            .O(N__12180),
            .I(N__12174));
    CascadeMux I__1866 (
            .O(N__12177),
            .I(N__12171));
    CascadeBuf I__1865 (
            .O(N__12174),
            .I(N__12168));
    CascadeBuf I__1864 (
            .O(N__12171),
            .I(N__12165));
    CascadeMux I__1863 (
            .O(N__12168),
            .I(N__12162));
    CascadeMux I__1862 (
            .O(N__12165),
            .I(N__12159));
    CascadeBuf I__1861 (
            .O(N__12162),
            .I(N__12156));
    CascadeBuf I__1860 (
            .O(N__12159),
            .I(N__12153));
    CascadeMux I__1859 (
            .O(N__12156),
            .I(N__12150));
    CascadeMux I__1858 (
            .O(N__12153),
            .I(N__12147));
    CascadeBuf I__1857 (
            .O(N__12150),
            .I(N__12144));
    CascadeBuf I__1856 (
            .O(N__12147),
            .I(N__12141));
    CascadeMux I__1855 (
            .O(N__12144),
            .I(N__12138));
    CascadeMux I__1854 (
            .O(N__12141),
            .I(N__12135));
    CascadeBuf I__1853 (
            .O(N__12138),
            .I(N__12132));
    CascadeBuf I__1852 (
            .O(N__12135),
            .I(N__12129));
    CascadeMux I__1851 (
            .O(N__12132),
            .I(N__12126));
    CascadeMux I__1850 (
            .O(N__12129),
            .I(N__12123));
    CascadeBuf I__1849 (
            .O(N__12126),
            .I(N__12120));
    CascadeBuf I__1848 (
            .O(N__12123),
            .I(N__12117));
    CascadeMux I__1847 (
            .O(N__12120),
            .I(N__12114));
    CascadeMux I__1846 (
            .O(N__12117),
            .I(N__12111));
    CascadeBuf I__1845 (
            .O(N__12114),
            .I(N__12108));
    CascadeBuf I__1844 (
            .O(N__12111),
            .I(N__12105));
    CascadeMux I__1843 (
            .O(N__12108),
            .I(N__12102));
    CascadeMux I__1842 (
            .O(N__12105),
            .I(N__12099));
    CascadeBuf I__1841 (
            .O(N__12102),
            .I(N__12096));
    CascadeBuf I__1840 (
            .O(N__12099),
            .I(N__12093));
    CascadeMux I__1839 (
            .O(N__12096),
            .I(N__12090));
    CascadeMux I__1838 (
            .O(N__12093),
            .I(N__12087));
    CascadeBuf I__1837 (
            .O(N__12090),
            .I(N__12084));
    CascadeBuf I__1836 (
            .O(N__12087),
            .I(N__12081));
    CascadeMux I__1835 (
            .O(N__12084),
            .I(N__12078));
    CascadeMux I__1834 (
            .O(N__12081),
            .I(N__12075));
    CascadeBuf I__1833 (
            .O(N__12078),
            .I(N__12072));
    CascadeBuf I__1832 (
            .O(N__12075),
            .I(N__12069));
    CascadeMux I__1831 (
            .O(N__12072),
            .I(N__12066));
    CascadeMux I__1830 (
            .O(N__12069),
            .I(N__12063));
    CascadeBuf I__1829 (
            .O(N__12066),
            .I(N__12060));
    CascadeBuf I__1828 (
            .O(N__12063),
            .I(N__12057));
    CascadeMux I__1827 (
            .O(N__12060),
            .I(N__12054));
    CascadeMux I__1826 (
            .O(N__12057),
            .I(N__12051));
    CascadeBuf I__1825 (
            .O(N__12054),
            .I(N__12048));
    CascadeBuf I__1824 (
            .O(N__12051),
            .I(N__12045));
    CascadeMux I__1823 (
            .O(N__12048),
            .I(N__12042));
    CascadeMux I__1822 (
            .O(N__12045),
            .I(N__12039));
    CascadeBuf I__1821 (
            .O(N__12042),
            .I(N__12036));
    CascadeBuf I__1820 (
            .O(N__12039),
            .I(N__12033));
    CascadeMux I__1819 (
            .O(N__12036),
            .I(N__12030));
    CascadeMux I__1818 (
            .O(N__12033),
            .I(N__12027));
    InMux I__1817 (
            .O(N__12030),
            .I(N__12024));
    InMux I__1816 (
            .O(N__12027),
            .I(N__12021));
    LocalMux I__1815 (
            .O(N__12024),
            .I(N__12018));
    LocalMux I__1814 (
            .O(N__12021),
            .I(N__12015));
    Span12Mux_v I__1813 (
            .O(N__12018),
            .I(N__12012));
    Span12Mux_s9_v I__1812 (
            .O(N__12015),
            .I(N__12009));
    Span12Mux_h I__1811 (
            .O(N__12012),
            .I(N__12006));
    Span12Mux_v I__1810 (
            .O(N__12009),
            .I(N__12003));
    Odrv12 I__1809 (
            .O(N__12006),
            .I(RX_ADDR_7));
    Odrv12 I__1808 (
            .O(N__12003),
            .I(RX_ADDR_7));
    InMux I__1807 (
            .O(N__11998),
            .I(\receive_module.n3699 ));
    InMux I__1806 (
            .O(N__11995),
            .I(N__11992));
    LocalMux I__1805 (
            .O(N__11992),
            .I(N__11989));
    Span4Mux_v I__1804 (
            .O(N__11989),
            .I(N__11983));
    InMux I__1803 (
            .O(N__11988),
            .I(N__11978));
    InMux I__1802 (
            .O(N__11987),
            .I(N__11978));
    InMux I__1801 (
            .O(N__11986),
            .I(N__11975));
    Odrv4 I__1800 (
            .O(N__11983),
            .I(\receive_module.O_Y_2 ));
    LocalMux I__1799 (
            .O(N__11978),
            .I(\receive_module.O_Y_2 ));
    LocalMux I__1798 (
            .O(N__11975),
            .I(\receive_module.O_Y_2 ));
    CascadeMux I__1797 (
            .O(N__11968),
            .I(N__11965));
    InMux I__1796 (
            .O(N__11965),
            .I(N__11962));
    LocalMux I__1795 (
            .O(N__11962),
            .I(\receive_module.O_X_8 ));
    CascadeMux I__1794 (
            .O(N__11959),
            .I(N__11955));
    CascadeMux I__1793 (
            .O(N__11958),
            .I(N__11952));
    CascadeBuf I__1792 (
            .O(N__11955),
            .I(N__11949));
    CascadeBuf I__1791 (
            .O(N__11952),
            .I(N__11946));
    CascadeMux I__1790 (
            .O(N__11949),
            .I(N__11943));
    CascadeMux I__1789 (
            .O(N__11946),
            .I(N__11940));
    CascadeBuf I__1788 (
            .O(N__11943),
            .I(N__11937));
    CascadeBuf I__1787 (
            .O(N__11940),
            .I(N__11934));
    CascadeMux I__1786 (
            .O(N__11937),
            .I(N__11931));
    CascadeMux I__1785 (
            .O(N__11934),
            .I(N__11928));
    CascadeBuf I__1784 (
            .O(N__11931),
            .I(N__11925));
    CascadeBuf I__1783 (
            .O(N__11928),
            .I(N__11922));
    CascadeMux I__1782 (
            .O(N__11925),
            .I(N__11919));
    CascadeMux I__1781 (
            .O(N__11922),
            .I(N__11916));
    CascadeBuf I__1780 (
            .O(N__11919),
            .I(N__11913));
    CascadeBuf I__1779 (
            .O(N__11916),
            .I(N__11910));
    CascadeMux I__1778 (
            .O(N__11913),
            .I(N__11907));
    CascadeMux I__1777 (
            .O(N__11910),
            .I(N__11904));
    CascadeBuf I__1776 (
            .O(N__11907),
            .I(N__11901));
    CascadeBuf I__1775 (
            .O(N__11904),
            .I(N__11898));
    CascadeMux I__1774 (
            .O(N__11901),
            .I(N__11895));
    CascadeMux I__1773 (
            .O(N__11898),
            .I(N__11892));
    CascadeBuf I__1772 (
            .O(N__11895),
            .I(N__11889));
    CascadeBuf I__1771 (
            .O(N__11892),
            .I(N__11886));
    CascadeMux I__1770 (
            .O(N__11889),
            .I(N__11883));
    CascadeMux I__1769 (
            .O(N__11886),
            .I(N__11880));
    CascadeBuf I__1768 (
            .O(N__11883),
            .I(N__11877));
    CascadeBuf I__1767 (
            .O(N__11880),
            .I(N__11874));
    CascadeMux I__1766 (
            .O(N__11877),
            .I(N__11871));
    CascadeMux I__1765 (
            .O(N__11874),
            .I(N__11868));
    CascadeBuf I__1764 (
            .O(N__11871),
            .I(N__11865));
    CascadeBuf I__1763 (
            .O(N__11868),
            .I(N__11862));
    CascadeMux I__1762 (
            .O(N__11865),
            .I(N__11859));
    CascadeMux I__1761 (
            .O(N__11862),
            .I(N__11856));
    CascadeBuf I__1760 (
            .O(N__11859),
            .I(N__11853));
    CascadeBuf I__1759 (
            .O(N__11856),
            .I(N__11850));
    CascadeMux I__1758 (
            .O(N__11853),
            .I(N__11847));
    CascadeMux I__1757 (
            .O(N__11850),
            .I(N__11844));
    CascadeBuf I__1756 (
            .O(N__11847),
            .I(N__11841));
    CascadeBuf I__1755 (
            .O(N__11844),
            .I(N__11838));
    CascadeMux I__1754 (
            .O(N__11841),
            .I(N__11835));
    CascadeMux I__1753 (
            .O(N__11838),
            .I(N__11832));
    CascadeBuf I__1752 (
            .O(N__11835),
            .I(N__11829));
    CascadeBuf I__1751 (
            .O(N__11832),
            .I(N__11826));
    CascadeMux I__1750 (
            .O(N__11829),
            .I(N__11823));
    CascadeMux I__1749 (
            .O(N__11826),
            .I(N__11820));
    CascadeBuf I__1748 (
            .O(N__11823),
            .I(N__11817));
    CascadeBuf I__1747 (
            .O(N__11820),
            .I(N__11814));
    CascadeMux I__1746 (
            .O(N__11817),
            .I(N__11811));
    CascadeMux I__1745 (
            .O(N__11814),
            .I(N__11808));
    CascadeBuf I__1744 (
            .O(N__11811),
            .I(N__11805));
    CascadeBuf I__1743 (
            .O(N__11808),
            .I(N__11802));
    CascadeMux I__1742 (
            .O(N__11805),
            .I(N__11799));
    CascadeMux I__1741 (
            .O(N__11802),
            .I(N__11796));
    CascadeBuf I__1740 (
            .O(N__11799),
            .I(N__11793));
    CascadeBuf I__1739 (
            .O(N__11796),
            .I(N__11790));
    CascadeMux I__1738 (
            .O(N__11793),
            .I(N__11787));
    CascadeMux I__1737 (
            .O(N__11790),
            .I(N__11784));
    CascadeBuf I__1736 (
            .O(N__11787),
            .I(N__11781));
    CascadeBuf I__1735 (
            .O(N__11784),
            .I(N__11778));
    CascadeMux I__1734 (
            .O(N__11781),
            .I(N__11775));
    CascadeMux I__1733 (
            .O(N__11778),
            .I(N__11772));
    InMux I__1732 (
            .O(N__11775),
            .I(N__11769));
    InMux I__1731 (
            .O(N__11772),
            .I(N__11766));
    LocalMux I__1730 (
            .O(N__11769),
            .I(N__11763));
    LocalMux I__1729 (
            .O(N__11766),
            .I(N__11760));
    Span4Mux_s1_v I__1728 (
            .O(N__11763),
            .I(N__11757));
    Span12Mux_s7_v I__1727 (
            .O(N__11760),
            .I(N__11754));
    Span4Mux_h I__1726 (
            .O(N__11757),
            .I(N__11751));
    Span12Mux_h I__1725 (
            .O(N__11754),
            .I(N__11748));
    Sp12to4 I__1724 (
            .O(N__11751),
            .I(N__11745));
    Span12Mux_v I__1723 (
            .O(N__11748),
            .I(N__11742));
    Span12Mux_s11_v I__1722 (
            .O(N__11745),
            .I(N__11739));
    Odrv12 I__1721 (
            .O(N__11742),
            .I(RX_ADDR_8));
    Odrv12 I__1720 (
            .O(N__11739),
            .I(RX_ADDR_8));
    InMux I__1719 (
            .O(N__11734),
            .I(\receive_module.n3700 ));
    InMux I__1718 (
            .O(N__11731),
            .I(N__11728));
    LocalMux I__1717 (
            .O(N__11728),
            .I(\transmit_module.ADDR_Y_COMPONENT_10 ));
    InMux I__1716 (
            .O(N__11725),
            .I(N__11722));
    LocalMux I__1715 (
            .O(N__11722),
            .I(N__11719));
    Span4Mux_v I__1714 (
            .O(N__11719),
            .I(N__11716));
    Odrv4 I__1713 (
            .O(N__11716),
            .I(\transmit_module.n209 ));
    InMux I__1712 (
            .O(N__11713),
            .I(N__11710));
    LocalMux I__1711 (
            .O(N__11710),
            .I(N__11706));
    InMux I__1710 (
            .O(N__11709),
            .I(N__11703));
    Span4Mux_v I__1709 (
            .O(N__11706),
            .I(N__11700));
    LocalMux I__1708 (
            .O(N__11703),
            .I(\transmit_module.n178 ));
    Odrv4 I__1707 (
            .O(N__11700),
            .I(\transmit_module.n178 ));
    CascadeMux I__1706 (
            .O(N__11695),
            .I(\transmit_module.n209_cascade_ ));
    CEMux I__1705 (
            .O(N__11692),
            .I(N__11688));
    CEMux I__1704 (
            .O(N__11691),
            .I(N__11685));
    LocalMux I__1703 (
            .O(N__11688),
            .I(N__11682));
    LocalMux I__1702 (
            .O(N__11685),
            .I(N__11679));
    Span4Mux_h I__1701 (
            .O(N__11682),
            .I(N__11676));
    Span4Mux_h I__1700 (
            .O(N__11679),
            .I(N__11673));
    Odrv4 I__1699 (
            .O(N__11676),
            .I(n2283));
    Odrv4 I__1698 (
            .O(N__11673),
            .I(n2283));
    InMux I__1697 (
            .O(N__11668),
            .I(N__11665));
    LocalMux I__1696 (
            .O(N__11665),
            .I(old_HS));
    CascadeMux I__1695 (
            .O(N__11662),
            .I(N__11659));
    CascadeBuf I__1694 (
            .O(N__11659),
            .I(N__11656));
    CascadeMux I__1693 (
            .O(N__11656),
            .I(N__11652));
    CascadeMux I__1692 (
            .O(N__11655),
            .I(N__11649));
    CascadeBuf I__1691 (
            .O(N__11652),
            .I(N__11646));
    CascadeBuf I__1690 (
            .O(N__11649),
            .I(N__11643));
    CascadeMux I__1689 (
            .O(N__11646),
            .I(N__11640));
    CascadeMux I__1688 (
            .O(N__11643),
            .I(N__11637));
    CascadeBuf I__1687 (
            .O(N__11640),
            .I(N__11634));
    CascadeBuf I__1686 (
            .O(N__11637),
            .I(N__11631));
    CascadeMux I__1685 (
            .O(N__11634),
            .I(N__11628));
    CascadeMux I__1684 (
            .O(N__11631),
            .I(N__11625));
    CascadeBuf I__1683 (
            .O(N__11628),
            .I(N__11622));
    CascadeBuf I__1682 (
            .O(N__11625),
            .I(N__11619));
    CascadeMux I__1681 (
            .O(N__11622),
            .I(N__11616));
    CascadeMux I__1680 (
            .O(N__11619),
            .I(N__11613));
    CascadeBuf I__1679 (
            .O(N__11616),
            .I(N__11610));
    CascadeBuf I__1678 (
            .O(N__11613),
            .I(N__11607));
    CascadeMux I__1677 (
            .O(N__11610),
            .I(N__11604));
    CascadeMux I__1676 (
            .O(N__11607),
            .I(N__11601));
    CascadeBuf I__1675 (
            .O(N__11604),
            .I(N__11598));
    CascadeBuf I__1674 (
            .O(N__11601),
            .I(N__11595));
    CascadeMux I__1673 (
            .O(N__11598),
            .I(N__11592));
    CascadeMux I__1672 (
            .O(N__11595),
            .I(N__11589));
    CascadeBuf I__1671 (
            .O(N__11592),
            .I(N__11586));
    CascadeBuf I__1670 (
            .O(N__11589),
            .I(N__11583));
    CascadeMux I__1669 (
            .O(N__11586),
            .I(N__11580));
    CascadeMux I__1668 (
            .O(N__11583),
            .I(N__11577));
    CascadeBuf I__1667 (
            .O(N__11580),
            .I(N__11574));
    CascadeBuf I__1666 (
            .O(N__11577),
            .I(N__11571));
    CascadeMux I__1665 (
            .O(N__11574),
            .I(N__11568));
    CascadeMux I__1664 (
            .O(N__11571),
            .I(N__11565));
    CascadeBuf I__1663 (
            .O(N__11568),
            .I(N__11562));
    CascadeBuf I__1662 (
            .O(N__11565),
            .I(N__11559));
    CascadeMux I__1661 (
            .O(N__11562),
            .I(N__11556));
    CascadeMux I__1660 (
            .O(N__11559),
            .I(N__11553));
    CascadeBuf I__1659 (
            .O(N__11556),
            .I(N__11550));
    CascadeBuf I__1658 (
            .O(N__11553),
            .I(N__11547));
    CascadeMux I__1657 (
            .O(N__11550),
            .I(N__11544));
    CascadeMux I__1656 (
            .O(N__11547),
            .I(N__11541));
    CascadeBuf I__1655 (
            .O(N__11544),
            .I(N__11538));
    CascadeBuf I__1654 (
            .O(N__11541),
            .I(N__11535));
    CascadeMux I__1653 (
            .O(N__11538),
            .I(N__11532));
    CascadeMux I__1652 (
            .O(N__11535),
            .I(N__11529));
    CascadeBuf I__1651 (
            .O(N__11532),
            .I(N__11526));
    CascadeBuf I__1650 (
            .O(N__11529),
            .I(N__11523));
    CascadeMux I__1649 (
            .O(N__11526),
            .I(N__11520));
    CascadeMux I__1648 (
            .O(N__11523),
            .I(N__11517));
    CascadeBuf I__1647 (
            .O(N__11520),
            .I(N__11514));
    CascadeBuf I__1646 (
            .O(N__11517),
            .I(N__11511));
    CascadeMux I__1645 (
            .O(N__11514),
            .I(N__11508));
    CascadeMux I__1644 (
            .O(N__11511),
            .I(N__11505));
    CascadeBuf I__1643 (
            .O(N__11508),
            .I(N__11502));
    CascadeBuf I__1642 (
            .O(N__11505),
            .I(N__11499));
    CascadeMux I__1641 (
            .O(N__11502),
            .I(N__11496));
    CascadeMux I__1640 (
            .O(N__11499),
            .I(N__11493));
    CascadeBuf I__1639 (
            .O(N__11496),
            .I(N__11490));
    CascadeBuf I__1638 (
            .O(N__11493),
            .I(N__11487));
    CascadeMux I__1637 (
            .O(N__11490),
            .I(N__11484));
    CascadeMux I__1636 (
            .O(N__11487),
            .I(N__11481));
    InMux I__1635 (
            .O(N__11484),
            .I(N__11478));
    CascadeBuf I__1634 (
            .O(N__11481),
            .I(N__11475));
    LocalMux I__1633 (
            .O(N__11478),
            .I(N__11472));
    CascadeMux I__1632 (
            .O(N__11475),
            .I(N__11469));
    Span4Mux_s2_v I__1631 (
            .O(N__11472),
            .I(N__11466));
    InMux I__1630 (
            .O(N__11469),
            .I(N__11463));
    Span4Mux_h I__1629 (
            .O(N__11466),
            .I(N__11460));
    LocalMux I__1628 (
            .O(N__11463),
            .I(N__11457));
    Sp12to4 I__1627 (
            .O(N__11460),
            .I(N__11454));
    Span4Mux_s2_v I__1626 (
            .O(N__11457),
            .I(N__11451));
    Span12Mux_s10_v I__1625 (
            .O(N__11454),
            .I(N__11448));
    Sp12to4 I__1624 (
            .O(N__11451),
            .I(N__11445));
    Span12Mux_h I__1623 (
            .O(N__11448),
            .I(N__11440));
    Span12Mux_s10_v I__1622 (
            .O(N__11445),
            .I(N__11440));
    Span12Mux_v I__1621 (
            .O(N__11440),
            .I(N__11437));
    Odrv12 I__1620 (
            .O(N__11437),
            .I(RX_ADDR_3));
    InMux I__1619 (
            .O(N__11434),
            .I(bfn_13_10_0_));
    CascadeMux I__1618 (
            .O(N__11431),
            .I(N__11428));
    CascadeBuf I__1617 (
            .O(N__11428),
            .I(N__11424));
    CascadeMux I__1616 (
            .O(N__11427),
            .I(N__11421));
    CascadeMux I__1615 (
            .O(N__11424),
            .I(N__11418));
    CascadeBuf I__1614 (
            .O(N__11421),
            .I(N__11415));
    CascadeBuf I__1613 (
            .O(N__11418),
            .I(N__11412));
    CascadeMux I__1612 (
            .O(N__11415),
            .I(N__11409));
    CascadeMux I__1611 (
            .O(N__11412),
            .I(N__11406));
    CascadeBuf I__1610 (
            .O(N__11409),
            .I(N__11403));
    CascadeBuf I__1609 (
            .O(N__11406),
            .I(N__11400));
    CascadeMux I__1608 (
            .O(N__11403),
            .I(N__11397));
    CascadeMux I__1607 (
            .O(N__11400),
            .I(N__11394));
    CascadeBuf I__1606 (
            .O(N__11397),
            .I(N__11391));
    CascadeBuf I__1605 (
            .O(N__11394),
            .I(N__11388));
    CascadeMux I__1604 (
            .O(N__11391),
            .I(N__11385));
    CascadeMux I__1603 (
            .O(N__11388),
            .I(N__11382));
    CascadeBuf I__1602 (
            .O(N__11385),
            .I(N__11379));
    CascadeBuf I__1601 (
            .O(N__11382),
            .I(N__11376));
    CascadeMux I__1600 (
            .O(N__11379),
            .I(N__11373));
    CascadeMux I__1599 (
            .O(N__11376),
            .I(N__11370));
    CascadeBuf I__1598 (
            .O(N__11373),
            .I(N__11367));
    CascadeBuf I__1597 (
            .O(N__11370),
            .I(N__11364));
    CascadeMux I__1596 (
            .O(N__11367),
            .I(N__11361));
    CascadeMux I__1595 (
            .O(N__11364),
            .I(N__11358));
    CascadeBuf I__1594 (
            .O(N__11361),
            .I(N__11355));
    CascadeBuf I__1593 (
            .O(N__11358),
            .I(N__11352));
    CascadeMux I__1592 (
            .O(N__11355),
            .I(N__11349));
    CascadeMux I__1591 (
            .O(N__11352),
            .I(N__11346));
    CascadeBuf I__1590 (
            .O(N__11349),
            .I(N__11343));
    CascadeBuf I__1589 (
            .O(N__11346),
            .I(N__11340));
    CascadeMux I__1588 (
            .O(N__11343),
            .I(N__11337));
    CascadeMux I__1587 (
            .O(N__11340),
            .I(N__11334));
    CascadeBuf I__1586 (
            .O(N__11337),
            .I(N__11331));
    CascadeBuf I__1585 (
            .O(N__11334),
            .I(N__11328));
    CascadeMux I__1584 (
            .O(N__11331),
            .I(N__11325));
    CascadeMux I__1583 (
            .O(N__11328),
            .I(N__11322));
    CascadeBuf I__1582 (
            .O(N__11325),
            .I(N__11319));
    CascadeBuf I__1581 (
            .O(N__11322),
            .I(N__11316));
    CascadeMux I__1580 (
            .O(N__11319),
            .I(N__11313));
    CascadeMux I__1579 (
            .O(N__11316),
            .I(N__11310));
    CascadeBuf I__1578 (
            .O(N__11313),
            .I(N__11307));
    CascadeBuf I__1577 (
            .O(N__11310),
            .I(N__11304));
    CascadeMux I__1576 (
            .O(N__11307),
            .I(N__11301));
    CascadeMux I__1575 (
            .O(N__11304),
            .I(N__11298));
    CascadeBuf I__1574 (
            .O(N__11301),
            .I(N__11295));
    CascadeBuf I__1573 (
            .O(N__11298),
            .I(N__11292));
    CascadeMux I__1572 (
            .O(N__11295),
            .I(N__11289));
    CascadeMux I__1571 (
            .O(N__11292),
            .I(N__11286));
    CascadeBuf I__1570 (
            .O(N__11289),
            .I(N__11283));
    CascadeBuf I__1569 (
            .O(N__11286),
            .I(N__11280));
    CascadeMux I__1568 (
            .O(N__11283),
            .I(N__11277));
    CascadeMux I__1567 (
            .O(N__11280),
            .I(N__11274));
    CascadeBuf I__1566 (
            .O(N__11277),
            .I(N__11271));
    CascadeBuf I__1565 (
            .O(N__11274),
            .I(N__11268));
    CascadeMux I__1564 (
            .O(N__11271),
            .I(N__11265));
    CascadeMux I__1563 (
            .O(N__11268),
            .I(N__11262));
    CascadeBuf I__1562 (
            .O(N__11265),
            .I(N__11259));
    CascadeBuf I__1561 (
            .O(N__11262),
            .I(N__11256));
    CascadeMux I__1560 (
            .O(N__11259),
            .I(N__11253));
    CascadeMux I__1559 (
            .O(N__11256),
            .I(N__11250));
    CascadeBuf I__1558 (
            .O(N__11253),
            .I(N__11247));
    InMux I__1557 (
            .O(N__11250),
            .I(N__11244));
    CascadeMux I__1556 (
            .O(N__11247),
            .I(N__11241));
    LocalMux I__1555 (
            .O(N__11244),
            .I(N__11238));
    InMux I__1554 (
            .O(N__11241),
            .I(N__11235));
    Span12Mux_s1_v I__1553 (
            .O(N__11238),
            .I(N__11232));
    LocalMux I__1552 (
            .O(N__11235),
            .I(N__11229));
    Span12Mux_h I__1551 (
            .O(N__11232),
            .I(N__11226));
    Span12Mux_s10_v I__1550 (
            .O(N__11229),
            .I(N__11223));
    Span12Mux_v I__1549 (
            .O(N__11226),
            .I(N__11220));
    Span12Mux_v I__1548 (
            .O(N__11223),
            .I(N__11217));
    Odrv12 I__1547 (
            .O(N__11220),
            .I(RX_ADDR_4));
    Odrv12 I__1546 (
            .O(N__11217),
            .I(RX_ADDR_4));
    InMux I__1545 (
            .O(N__11212),
            .I(\receive_module.rx_counter.n3650 ));
    CascadeMux I__1544 (
            .O(N__11209),
            .I(N__11205));
    CascadeMux I__1543 (
            .O(N__11208),
            .I(N__11202));
    CascadeBuf I__1542 (
            .O(N__11205),
            .I(N__11199));
    CascadeBuf I__1541 (
            .O(N__11202),
            .I(N__11196));
    CascadeMux I__1540 (
            .O(N__11199),
            .I(N__11193));
    CascadeMux I__1539 (
            .O(N__11196),
            .I(N__11190));
    CascadeBuf I__1538 (
            .O(N__11193),
            .I(N__11187));
    CascadeBuf I__1537 (
            .O(N__11190),
            .I(N__11184));
    CascadeMux I__1536 (
            .O(N__11187),
            .I(N__11181));
    CascadeMux I__1535 (
            .O(N__11184),
            .I(N__11178));
    CascadeBuf I__1534 (
            .O(N__11181),
            .I(N__11175));
    CascadeBuf I__1533 (
            .O(N__11178),
            .I(N__11172));
    CascadeMux I__1532 (
            .O(N__11175),
            .I(N__11169));
    CascadeMux I__1531 (
            .O(N__11172),
            .I(N__11166));
    CascadeBuf I__1530 (
            .O(N__11169),
            .I(N__11163));
    CascadeBuf I__1529 (
            .O(N__11166),
            .I(N__11160));
    CascadeMux I__1528 (
            .O(N__11163),
            .I(N__11157));
    CascadeMux I__1527 (
            .O(N__11160),
            .I(N__11154));
    CascadeBuf I__1526 (
            .O(N__11157),
            .I(N__11151));
    CascadeBuf I__1525 (
            .O(N__11154),
            .I(N__11148));
    CascadeMux I__1524 (
            .O(N__11151),
            .I(N__11145));
    CascadeMux I__1523 (
            .O(N__11148),
            .I(N__11142));
    CascadeBuf I__1522 (
            .O(N__11145),
            .I(N__11139));
    CascadeBuf I__1521 (
            .O(N__11142),
            .I(N__11136));
    CascadeMux I__1520 (
            .O(N__11139),
            .I(N__11133));
    CascadeMux I__1519 (
            .O(N__11136),
            .I(N__11130));
    CascadeBuf I__1518 (
            .O(N__11133),
            .I(N__11127));
    CascadeBuf I__1517 (
            .O(N__11130),
            .I(N__11124));
    CascadeMux I__1516 (
            .O(N__11127),
            .I(N__11121));
    CascadeMux I__1515 (
            .O(N__11124),
            .I(N__11118));
    CascadeBuf I__1514 (
            .O(N__11121),
            .I(N__11115));
    CascadeBuf I__1513 (
            .O(N__11118),
            .I(N__11112));
    CascadeMux I__1512 (
            .O(N__11115),
            .I(N__11109));
    CascadeMux I__1511 (
            .O(N__11112),
            .I(N__11106));
    CascadeBuf I__1510 (
            .O(N__11109),
            .I(N__11103));
    CascadeBuf I__1509 (
            .O(N__11106),
            .I(N__11100));
    CascadeMux I__1508 (
            .O(N__11103),
            .I(N__11097));
    CascadeMux I__1507 (
            .O(N__11100),
            .I(N__11094));
    CascadeBuf I__1506 (
            .O(N__11097),
            .I(N__11091));
    CascadeBuf I__1505 (
            .O(N__11094),
            .I(N__11088));
    CascadeMux I__1504 (
            .O(N__11091),
            .I(N__11085));
    CascadeMux I__1503 (
            .O(N__11088),
            .I(N__11082));
    CascadeBuf I__1502 (
            .O(N__11085),
            .I(N__11079));
    CascadeBuf I__1501 (
            .O(N__11082),
            .I(N__11076));
    CascadeMux I__1500 (
            .O(N__11079),
            .I(N__11073));
    CascadeMux I__1499 (
            .O(N__11076),
            .I(N__11070));
    CascadeBuf I__1498 (
            .O(N__11073),
            .I(N__11067));
    CascadeBuf I__1497 (
            .O(N__11070),
            .I(N__11064));
    CascadeMux I__1496 (
            .O(N__11067),
            .I(N__11061));
    CascadeMux I__1495 (
            .O(N__11064),
            .I(N__11058));
    CascadeBuf I__1494 (
            .O(N__11061),
            .I(N__11055));
    CascadeBuf I__1493 (
            .O(N__11058),
            .I(N__11052));
    CascadeMux I__1492 (
            .O(N__11055),
            .I(N__11049));
    CascadeMux I__1491 (
            .O(N__11052),
            .I(N__11046));
    CascadeBuf I__1490 (
            .O(N__11049),
            .I(N__11043));
    CascadeBuf I__1489 (
            .O(N__11046),
            .I(N__11040));
    CascadeMux I__1488 (
            .O(N__11043),
            .I(N__11037));
    CascadeMux I__1487 (
            .O(N__11040),
            .I(N__11034));
    CascadeBuf I__1486 (
            .O(N__11037),
            .I(N__11031));
    CascadeBuf I__1485 (
            .O(N__11034),
            .I(N__11028));
    CascadeMux I__1484 (
            .O(N__11031),
            .I(N__11025));
    CascadeMux I__1483 (
            .O(N__11028),
            .I(N__11022));
    InMux I__1482 (
            .O(N__11025),
            .I(N__11019));
    InMux I__1481 (
            .O(N__11022),
            .I(N__11016));
    LocalMux I__1480 (
            .O(N__11019),
            .I(N__11013));
    LocalMux I__1479 (
            .O(N__11016),
            .I(N__11010));
    Span12Mux_v I__1478 (
            .O(N__11013),
            .I(N__11007));
    Span12Mux_h I__1477 (
            .O(N__11010),
            .I(N__11004));
    Span12Mux_h I__1476 (
            .O(N__11007),
            .I(N__10999));
    Span12Mux_v I__1475 (
            .O(N__11004),
            .I(N__10999));
    Odrv12 I__1474 (
            .O(N__10999),
            .I(RX_ADDR_5));
    InMux I__1473 (
            .O(N__10996),
            .I(\receive_module.rx_counter.n3651 ));
    InMux I__1472 (
            .O(N__10993),
            .I(N__10990));
    LocalMux I__1471 (
            .O(N__10990),
            .I(N__10987));
    Span4Mux_v I__1470 (
            .O(N__10987),
            .I(N__10984));
    Odrv4 I__1469 (
            .O(N__10984),
            .I(\transmit_module.Y_DELTA_PATTERN_81 ));
    InMux I__1468 (
            .O(N__10981),
            .I(N__10978));
    LocalMux I__1467 (
            .O(N__10978),
            .I(\transmit_module.Y_DELTA_PATTERN_69 ));
    InMux I__1466 (
            .O(N__10975),
            .I(N__10972));
    LocalMux I__1465 (
            .O(N__10972),
            .I(\transmit_module.Y_DELTA_PATTERN_68 ));
    InMux I__1464 (
            .O(N__10969),
            .I(N__10966));
    LocalMux I__1463 (
            .O(N__10966),
            .I(N__10963));
    Odrv4 I__1462 (
            .O(N__10963),
            .I(\transmit_module.Y_DELTA_PATTERN_78 ));
    InMux I__1461 (
            .O(N__10960),
            .I(N__10957));
    LocalMux I__1460 (
            .O(N__10957),
            .I(\transmit_module.Y_DELTA_PATTERN_62 ));
    InMux I__1459 (
            .O(N__10954),
            .I(N__10951));
    LocalMux I__1458 (
            .O(N__10951),
            .I(\transmit_module.Y_DELTA_PATTERN_66 ));
    InMux I__1457 (
            .O(N__10948),
            .I(N__10945));
    LocalMux I__1456 (
            .O(N__10945),
            .I(\transmit_module.Y_DELTA_PATTERN_65 ));
    InMux I__1455 (
            .O(N__10942),
            .I(N__10939));
    LocalMux I__1454 (
            .O(N__10939),
            .I(\transmit_module.Y_DELTA_PATTERN_80 ));
    InMux I__1453 (
            .O(N__10936),
            .I(N__10933));
    LocalMux I__1452 (
            .O(N__10933),
            .I(\transmit_module.Y_DELTA_PATTERN_79 ));
    InMux I__1451 (
            .O(N__10930),
            .I(N__10927));
    LocalMux I__1450 (
            .O(N__10927),
            .I(\transmit_module.Y_DELTA_PATTERN_57 ));
    CascadeMux I__1449 (
            .O(N__10924),
            .I(N__10919));
    InMux I__1448 (
            .O(N__10923),
            .I(N__10916));
    InMux I__1447 (
            .O(N__10922),
            .I(N__10913));
    InMux I__1446 (
            .O(N__10919),
            .I(N__10910));
    LocalMux I__1445 (
            .O(N__10916),
            .I(\transmit_module.video_signal_controller.VGA_Y_11 ));
    LocalMux I__1444 (
            .O(N__10913),
            .I(\transmit_module.video_signal_controller.VGA_Y_11 ));
    LocalMux I__1443 (
            .O(N__10910),
            .I(\transmit_module.video_signal_controller.VGA_Y_11 ));
    InMux I__1442 (
            .O(N__10903),
            .I(N__10898));
    InMux I__1441 (
            .O(N__10902),
            .I(N__10895));
    InMux I__1440 (
            .O(N__10901),
            .I(N__10892));
    LocalMux I__1439 (
            .O(N__10898),
            .I(\transmit_module.video_signal_controller.VGA_Y_10 ));
    LocalMux I__1438 (
            .O(N__10895),
            .I(\transmit_module.video_signal_controller.VGA_Y_10 ));
    LocalMux I__1437 (
            .O(N__10892),
            .I(\transmit_module.video_signal_controller.VGA_Y_10 ));
    InMux I__1436 (
            .O(N__10885),
            .I(N__10882));
    LocalMux I__1435 (
            .O(N__10882),
            .I(\transmit_module.video_signal_controller.n4218 ));
    CascadeMux I__1434 (
            .O(N__10879),
            .I(\transmit_module.n219_cascade_ ));
    CascadeMux I__1433 (
            .O(N__10876),
            .I(N__10873));
    CascadeBuf I__1432 (
            .O(N__10873),
            .I(N__10870));
    CascadeMux I__1431 (
            .O(N__10870),
            .I(N__10866));
    CascadeMux I__1430 (
            .O(N__10869),
            .I(N__10863));
    CascadeBuf I__1429 (
            .O(N__10866),
            .I(N__10860));
    CascadeBuf I__1428 (
            .O(N__10863),
            .I(N__10857));
    CascadeMux I__1427 (
            .O(N__10860),
            .I(N__10854));
    CascadeMux I__1426 (
            .O(N__10857),
            .I(N__10851));
    CascadeBuf I__1425 (
            .O(N__10854),
            .I(N__10848));
    CascadeBuf I__1424 (
            .O(N__10851),
            .I(N__10845));
    CascadeMux I__1423 (
            .O(N__10848),
            .I(N__10842));
    CascadeMux I__1422 (
            .O(N__10845),
            .I(N__10839));
    CascadeBuf I__1421 (
            .O(N__10842),
            .I(N__10836));
    CascadeBuf I__1420 (
            .O(N__10839),
            .I(N__10833));
    CascadeMux I__1419 (
            .O(N__10836),
            .I(N__10830));
    CascadeMux I__1418 (
            .O(N__10833),
            .I(N__10827));
    CascadeBuf I__1417 (
            .O(N__10830),
            .I(N__10824));
    CascadeBuf I__1416 (
            .O(N__10827),
            .I(N__10821));
    CascadeMux I__1415 (
            .O(N__10824),
            .I(N__10818));
    CascadeMux I__1414 (
            .O(N__10821),
            .I(N__10815));
    CascadeBuf I__1413 (
            .O(N__10818),
            .I(N__10812));
    CascadeBuf I__1412 (
            .O(N__10815),
            .I(N__10809));
    CascadeMux I__1411 (
            .O(N__10812),
            .I(N__10806));
    CascadeMux I__1410 (
            .O(N__10809),
            .I(N__10803));
    CascadeBuf I__1409 (
            .O(N__10806),
            .I(N__10800));
    CascadeBuf I__1408 (
            .O(N__10803),
            .I(N__10797));
    CascadeMux I__1407 (
            .O(N__10800),
            .I(N__10794));
    CascadeMux I__1406 (
            .O(N__10797),
            .I(N__10791));
    CascadeBuf I__1405 (
            .O(N__10794),
            .I(N__10788));
    CascadeBuf I__1404 (
            .O(N__10791),
            .I(N__10785));
    CascadeMux I__1403 (
            .O(N__10788),
            .I(N__10782));
    CascadeMux I__1402 (
            .O(N__10785),
            .I(N__10779));
    CascadeBuf I__1401 (
            .O(N__10782),
            .I(N__10776));
    CascadeBuf I__1400 (
            .O(N__10779),
            .I(N__10773));
    CascadeMux I__1399 (
            .O(N__10776),
            .I(N__10770));
    CascadeMux I__1398 (
            .O(N__10773),
            .I(N__10767));
    CascadeBuf I__1397 (
            .O(N__10770),
            .I(N__10764));
    CascadeBuf I__1396 (
            .O(N__10767),
            .I(N__10761));
    CascadeMux I__1395 (
            .O(N__10764),
            .I(N__10758));
    CascadeMux I__1394 (
            .O(N__10761),
            .I(N__10755));
    CascadeBuf I__1393 (
            .O(N__10758),
            .I(N__10752));
    CascadeBuf I__1392 (
            .O(N__10755),
            .I(N__10749));
    CascadeMux I__1391 (
            .O(N__10752),
            .I(N__10746));
    CascadeMux I__1390 (
            .O(N__10749),
            .I(N__10743));
    CascadeBuf I__1389 (
            .O(N__10746),
            .I(N__10740));
    CascadeBuf I__1388 (
            .O(N__10743),
            .I(N__10737));
    CascadeMux I__1387 (
            .O(N__10740),
            .I(N__10734));
    CascadeMux I__1386 (
            .O(N__10737),
            .I(N__10731));
    CascadeBuf I__1385 (
            .O(N__10734),
            .I(N__10728));
    CascadeBuf I__1384 (
            .O(N__10731),
            .I(N__10725));
    CascadeMux I__1383 (
            .O(N__10728),
            .I(N__10722));
    CascadeMux I__1382 (
            .O(N__10725),
            .I(N__10719));
    CascadeBuf I__1381 (
            .O(N__10722),
            .I(N__10716));
    CascadeBuf I__1380 (
            .O(N__10719),
            .I(N__10713));
    CascadeMux I__1379 (
            .O(N__10716),
            .I(N__10710));
    CascadeMux I__1378 (
            .O(N__10713),
            .I(N__10707));
    CascadeBuf I__1377 (
            .O(N__10710),
            .I(N__10704));
    CascadeBuf I__1376 (
            .O(N__10707),
            .I(N__10701));
    CascadeMux I__1375 (
            .O(N__10704),
            .I(N__10698));
    CascadeMux I__1374 (
            .O(N__10701),
            .I(N__10695));
    InMux I__1373 (
            .O(N__10698),
            .I(N__10692));
    CascadeBuf I__1372 (
            .O(N__10695),
            .I(N__10689));
    LocalMux I__1371 (
            .O(N__10692),
            .I(N__10686));
    CascadeMux I__1370 (
            .O(N__10689),
            .I(N__10683));
    Span4Mux_h I__1369 (
            .O(N__10686),
            .I(N__10680));
    InMux I__1368 (
            .O(N__10683),
            .I(N__10677));
    Sp12to4 I__1367 (
            .O(N__10680),
            .I(N__10674));
    LocalMux I__1366 (
            .O(N__10677),
            .I(N__10671));
    Span12Mux_v I__1365 (
            .O(N__10674),
            .I(N__10668));
    Span4Mux_h I__1364 (
            .O(N__10671),
            .I(N__10665));
    Span12Mux_h I__1363 (
            .O(N__10668),
            .I(N__10660));
    Sp12to4 I__1362 (
            .O(N__10665),
            .I(N__10660));
    Odrv12 I__1361 (
            .O(N__10660),
            .I(n28));
    IoInMux I__1360 (
            .O(N__10657),
            .I(N__10654));
    LocalMux I__1359 (
            .O(N__10654),
            .I(N__10651));
    IoSpan4Mux I__1358 (
            .O(N__10651),
            .I(N__10648));
    Span4Mux_s2_h I__1357 (
            .O(N__10648),
            .I(N__10645));
    Sp12to4 I__1356 (
            .O(N__10645),
            .I(N__10642));
    Odrv12 I__1355 (
            .O(N__10642),
            .I(n4210));
    CascadeMux I__1354 (
            .O(N__10639),
            .I(n4210_cascade_));
    InMux I__1353 (
            .O(N__10636),
            .I(N__10633));
    LocalMux I__1352 (
            .O(N__10633),
            .I(\transmit_module.Y_DELTA_PATTERN_64 ));
    InMux I__1351 (
            .O(N__10630),
            .I(N__10627));
    LocalMux I__1350 (
            .O(N__10627),
            .I(\transmit_module.Y_DELTA_PATTERN_67 ));
    InMux I__1349 (
            .O(N__10624),
            .I(N__10620));
    InMux I__1348 (
            .O(N__10623),
            .I(N__10617));
    LocalMux I__1347 (
            .O(N__10620),
            .I(\transmit_module.video_signal_controller.VGA_Y_7 ));
    LocalMux I__1346 (
            .O(N__10617),
            .I(\transmit_module.video_signal_controller.VGA_Y_7 ));
    InMux I__1345 (
            .O(N__10612),
            .I(\transmit_module.video_signal_controller.n3683 ));
    InMux I__1344 (
            .O(N__10609),
            .I(N__10605));
    InMux I__1343 (
            .O(N__10608),
            .I(N__10602));
    LocalMux I__1342 (
            .O(N__10605),
            .I(\transmit_module.video_signal_controller.VGA_Y_8 ));
    LocalMux I__1341 (
            .O(N__10602),
            .I(\transmit_module.video_signal_controller.VGA_Y_8 ));
    InMux I__1340 (
            .O(N__10597),
            .I(bfn_12_17_0_));
    InMux I__1339 (
            .O(N__10594),
            .I(\transmit_module.video_signal_controller.n3685 ));
    InMux I__1338 (
            .O(N__10591),
            .I(\transmit_module.video_signal_controller.n3686 ));
    InMux I__1337 (
            .O(N__10588),
            .I(\transmit_module.video_signal_controller.n3687 ));
    SRMux I__1336 (
            .O(N__10585),
            .I(N__10581));
    SRMux I__1335 (
            .O(N__10584),
            .I(N__10578));
    LocalMux I__1334 (
            .O(N__10581),
            .I(N__10575));
    LocalMux I__1333 (
            .O(N__10578),
            .I(N__10572));
    Span4Mux_h I__1332 (
            .O(N__10575),
            .I(N__10569));
    Span4Mux_v I__1331 (
            .O(N__10572),
            .I(N__10566));
    Odrv4 I__1330 (
            .O(N__10569),
            .I(\transmit_module.video_signal_controller.n2594 ));
    Odrv4 I__1329 (
            .O(N__10566),
            .I(\transmit_module.video_signal_controller.n2594 ));
    InMux I__1328 (
            .O(N__10561),
            .I(N__10556));
    InMux I__1327 (
            .O(N__10560),
            .I(N__10552));
    InMux I__1326 (
            .O(N__10559),
            .I(N__10549));
    LocalMux I__1325 (
            .O(N__10556),
            .I(N__10546));
    InMux I__1324 (
            .O(N__10555),
            .I(N__10543));
    LocalMux I__1323 (
            .O(N__10552),
            .I(\transmit_module.video_signal_controller.VGA_Y_3 ));
    LocalMux I__1322 (
            .O(N__10549),
            .I(\transmit_module.video_signal_controller.VGA_Y_3 ));
    Odrv4 I__1321 (
            .O(N__10546),
            .I(\transmit_module.video_signal_controller.VGA_Y_3 ));
    LocalMux I__1320 (
            .O(N__10543),
            .I(\transmit_module.video_signal_controller.VGA_Y_3 ));
    InMux I__1319 (
            .O(N__10534),
            .I(N__10531));
    LocalMux I__1318 (
            .O(N__10531),
            .I(\transmit_module.video_signal_controller.n4215 ));
    CascadeMux I__1317 (
            .O(N__10528),
            .I(N__10524));
    CascadeMux I__1316 (
            .O(N__10527),
            .I(N__10521));
    InMux I__1315 (
            .O(N__10524),
            .I(N__10517));
    InMux I__1314 (
            .O(N__10521),
            .I(N__10513));
    InMux I__1313 (
            .O(N__10520),
            .I(N__10510));
    LocalMux I__1312 (
            .O(N__10517),
            .I(N__10507));
    InMux I__1311 (
            .O(N__10516),
            .I(N__10504));
    LocalMux I__1310 (
            .O(N__10513),
            .I(\transmit_module.video_signal_controller.VGA_Y_4 ));
    LocalMux I__1309 (
            .O(N__10510),
            .I(\transmit_module.video_signal_controller.VGA_Y_4 ));
    Odrv4 I__1308 (
            .O(N__10507),
            .I(\transmit_module.video_signal_controller.VGA_Y_4 ));
    LocalMux I__1307 (
            .O(N__10504),
            .I(\transmit_module.video_signal_controller.VGA_Y_4 ));
    InMux I__1306 (
            .O(N__10495),
            .I(N__10491));
    InMux I__1305 (
            .O(N__10494),
            .I(N__10488));
    LocalMux I__1304 (
            .O(N__10491),
            .I(\transmit_module.video_signal_controller.n3892 ));
    LocalMux I__1303 (
            .O(N__10488),
            .I(\transmit_module.video_signal_controller.n3892 ));
    InMux I__1302 (
            .O(N__10483),
            .I(N__10478));
    InMux I__1301 (
            .O(N__10482),
            .I(N__10475));
    InMux I__1300 (
            .O(N__10481),
            .I(N__10472));
    LocalMux I__1299 (
            .O(N__10478),
            .I(\transmit_module.video_signal_controller.VGA_Y_9 ));
    LocalMux I__1298 (
            .O(N__10475),
            .I(\transmit_module.video_signal_controller.VGA_Y_9 ));
    LocalMux I__1297 (
            .O(N__10472),
            .I(\transmit_module.video_signal_controller.VGA_Y_9 ));
    CascadeMux I__1296 (
            .O(N__10465),
            .I(\transmit_module.video_signal_controller.VGA_VISIBLE_Y_N_553_cascade_ ));
    InMux I__1295 (
            .O(N__10462),
            .I(N__10459));
    LocalMux I__1294 (
            .O(N__10459),
            .I(\transmit_module.video_signal_controller.n3936 ));
    CascadeMux I__1293 (
            .O(N__10456),
            .I(\transmit_module.n3926_cascade_ ));
    CascadeMux I__1292 (
            .O(N__10453),
            .I(\transmit_module.video_signal_controller.n18_cascade_ ));
    InMux I__1291 (
            .O(N__10450),
            .I(N__10447));
    LocalMux I__1290 (
            .O(N__10447),
            .I(\transmit_module.video_signal_controller.n2219 ));
    InMux I__1289 (
            .O(N__10444),
            .I(N__10440));
    InMux I__1288 (
            .O(N__10443),
            .I(N__10437));
    LocalMux I__1287 (
            .O(N__10440),
            .I(\transmit_module.video_signal_controller.VGA_Y_0 ));
    LocalMux I__1286 (
            .O(N__10437),
            .I(\transmit_module.video_signal_controller.VGA_Y_0 ));
    InMux I__1285 (
            .O(N__10432),
            .I(bfn_12_16_0_));
    CascadeMux I__1284 (
            .O(N__10429),
            .I(N__10424));
    InMux I__1283 (
            .O(N__10428),
            .I(N__10420));
    InMux I__1282 (
            .O(N__10427),
            .I(N__10417));
    InMux I__1281 (
            .O(N__10424),
            .I(N__10412));
    InMux I__1280 (
            .O(N__10423),
            .I(N__10412));
    LocalMux I__1279 (
            .O(N__10420),
            .I(\transmit_module.video_signal_controller.VGA_Y_1 ));
    LocalMux I__1278 (
            .O(N__10417),
            .I(\transmit_module.video_signal_controller.VGA_Y_1 ));
    LocalMux I__1277 (
            .O(N__10412),
            .I(\transmit_module.video_signal_controller.VGA_Y_1 ));
    InMux I__1276 (
            .O(N__10405),
            .I(\transmit_module.video_signal_controller.n3677 ));
    InMux I__1275 (
            .O(N__10402),
            .I(N__10396));
    InMux I__1274 (
            .O(N__10401),
            .I(N__10393));
    InMux I__1273 (
            .O(N__10400),
            .I(N__10388));
    InMux I__1272 (
            .O(N__10399),
            .I(N__10388));
    LocalMux I__1271 (
            .O(N__10396),
            .I(\transmit_module.video_signal_controller.VGA_Y_2 ));
    LocalMux I__1270 (
            .O(N__10393),
            .I(\transmit_module.video_signal_controller.VGA_Y_2 ));
    LocalMux I__1269 (
            .O(N__10388),
            .I(\transmit_module.video_signal_controller.VGA_Y_2 ));
    InMux I__1268 (
            .O(N__10381),
            .I(\transmit_module.video_signal_controller.n3678 ));
    InMux I__1267 (
            .O(N__10378),
            .I(\transmit_module.video_signal_controller.n3679 ));
    InMux I__1266 (
            .O(N__10375),
            .I(\transmit_module.video_signal_controller.n3680 ));
    InMux I__1265 (
            .O(N__10372),
            .I(N__10367));
    InMux I__1264 (
            .O(N__10371),
            .I(N__10364));
    InMux I__1263 (
            .O(N__10370),
            .I(N__10361));
    LocalMux I__1262 (
            .O(N__10367),
            .I(\transmit_module.video_signal_controller.VGA_Y_5 ));
    LocalMux I__1261 (
            .O(N__10364),
            .I(\transmit_module.video_signal_controller.VGA_Y_5 ));
    LocalMux I__1260 (
            .O(N__10361),
            .I(\transmit_module.video_signal_controller.VGA_Y_5 ));
    InMux I__1259 (
            .O(N__10354),
            .I(\transmit_module.video_signal_controller.n3681 ));
    InMux I__1258 (
            .O(N__10351),
            .I(N__10346));
    InMux I__1257 (
            .O(N__10350),
            .I(N__10341));
    InMux I__1256 (
            .O(N__10349),
            .I(N__10341));
    LocalMux I__1255 (
            .O(N__10346),
            .I(\transmit_module.video_signal_controller.VGA_Y_6 ));
    LocalMux I__1254 (
            .O(N__10341),
            .I(\transmit_module.video_signal_controller.VGA_Y_6 ));
    InMux I__1253 (
            .O(N__10336),
            .I(\transmit_module.video_signal_controller.n3682 ));
    InMux I__1252 (
            .O(N__10333),
            .I(N__10330));
    LocalMux I__1251 (
            .O(N__10330),
            .I(\transmit_module.video_signal_controller.n4052 ));
    CascadeMux I__1250 (
            .O(N__10327),
            .I(\transmit_module.video_signal_controller.n4216_cascade_ ));
    InMux I__1249 (
            .O(N__10324),
            .I(N__10321));
    LocalMux I__1248 (
            .O(N__10321),
            .I(\transmit_module.video_signal_controller.n12 ));
    CascadeMux I__1247 (
            .O(N__10318),
            .I(\transmit_module.video_signal_controller.n2274_cascade_ ));
    InMux I__1246 (
            .O(N__10315),
            .I(N__10312));
    LocalMux I__1245 (
            .O(N__10312),
            .I(\transmit_module.video_signal_controller.SYNC_BUFF2 ));
    CascadeMux I__1244 (
            .O(N__10309),
            .I(N__10306));
    InMux I__1243 (
            .O(N__10306),
            .I(N__10303));
    LocalMux I__1242 (
            .O(N__10303),
            .I(\transmit_module.video_signal_controller.n3226 ));
    CascadeMux I__1241 (
            .O(N__10300),
            .I(N__10297));
    InMux I__1240 (
            .O(N__10297),
            .I(N__10294));
    LocalMux I__1239 (
            .O(N__10294),
            .I(\transmit_module.video_signal_controller.n2260 ));
    InMux I__1238 (
            .O(N__10291),
            .I(N__10285));
    InMux I__1237 (
            .O(N__10290),
            .I(N__10285));
    LocalMux I__1236 (
            .O(N__10285),
            .I(\transmit_module.video_signal_controller.n3917 ));
    CascadeMux I__1235 (
            .O(N__10282),
            .I(\transmit_module.video_signal_controller.n2260_cascade_ ));
    InMux I__1234 (
            .O(N__10279),
            .I(N__10276));
    LocalMux I__1233 (
            .O(N__10276),
            .I(\transmit_module.video_signal_controller.n4217 ));
    SRMux I__1232 (
            .O(N__10273),
            .I(N__10270));
    LocalMux I__1231 (
            .O(N__10270),
            .I(N__10266));
    SRMux I__1230 (
            .O(N__10269),
            .I(N__10263));
    Span4Mux_v I__1229 (
            .O(N__10266),
            .I(N__10257));
    LocalMux I__1228 (
            .O(N__10263),
            .I(N__10257));
    SRMux I__1227 (
            .O(N__10262),
            .I(N__10254));
    Span4Mux_v I__1226 (
            .O(N__10257),
            .I(N__10248));
    LocalMux I__1225 (
            .O(N__10254),
            .I(N__10248));
    SRMux I__1224 (
            .O(N__10253),
            .I(N__10245));
    Span4Mux_v I__1223 (
            .O(N__10248),
            .I(N__10240));
    LocalMux I__1222 (
            .O(N__10245),
            .I(N__10240));
    Span4Mux_h I__1221 (
            .O(N__10240),
            .I(N__10237));
    Odrv4 I__1220 (
            .O(N__10237),
            .I(n691));
    SRMux I__1219 (
            .O(N__10234),
            .I(N__10231));
    LocalMux I__1218 (
            .O(N__10231),
            .I(N__10228));
    Span4Mux_s2_v I__1217 (
            .O(N__10228),
            .I(N__10222));
    SRMux I__1216 (
            .O(N__10227),
            .I(N__10219));
    SRMux I__1215 (
            .O(N__10226),
            .I(N__10216));
    SRMux I__1214 (
            .O(N__10225),
            .I(N__10213));
    Span4Mux_v I__1213 (
            .O(N__10222),
            .I(N__10206));
    LocalMux I__1212 (
            .O(N__10219),
            .I(N__10206));
    LocalMux I__1211 (
            .O(N__10216),
            .I(N__10206));
    LocalMux I__1210 (
            .O(N__10213),
            .I(N__10203));
    Span4Mux_v I__1209 (
            .O(N__10206),
            .I(N__10198));
    Span4Mux_v I__1208 (
            .O(N__10203),
            .I(N__10198));
    Span4Mux_h I__1207 (
            .O(N__10198),
            .I(N__10195));
    Sp12to4 I__1206 (
            .O(N__10195),
            .I(N__10192));
    Odrv12 I__1205 (
            .O(N__10192),
            .I(\line_buffer.n626 ));
    SRMux I__1204 (
            .O(N__10189),
            .I(N__10185));
    SRMux I__1203 (
            .O(N__10188),
            .I(N__10182));
    LocalMux I__1202 (
            .O(N__10185),
            .I(N__10175));
    LocalMux I__1201 (
            .O(N__10182),
            .I(N__10175));
    SRMux I__1200 (
            .O(N__10181),
            .I(N__10172));
    SRMux I__1199 (
            .O(N__10180),
            .I(N__10169));
    Span4Mux_v I__1198 (
            .O(N__10175),
            .I(N__10164));
    LocalMux I__1197 (
            .O(N__10172),
            .I(N__10164));
    LocalMux I__1196 (
            .O(N__10169),
            .I(N__10161));
    Span4Mux_v I__1195 (
            .O(N__10164),
            .I(N__10158));
    Span4Mux_h I__1194 (
            .O(N__10161),
            .I(N__10155));
    Span4Mux_v I__1193 (
            .O(N__10158),
            .I(N__10152));
    Sp12to4 I__1192 (
            .O(N__10155),
            .I(N__10149));
    Span4Mux_v I__1191 (
            .O(N__10152),
            .I(N__10146));
    Span12Mux_h I__1190 (
            .O(N__10149),
            .I(N__10143));
    Span4Mux_v I__1189 (
            .O(N__10146),
            .I(N__10140));
    Odrv12 I__1188 (
            .O(N__10143),
            .I(\line_buffer.n561 ));
    Odrv4 I__1187 (
            .O(N__10140),
            .I(\line_buffer.n561 ));
    CascadeMux I__1186 (
            .O(N__10135),
            .I(\transmit_module.video_signal_controller.n3978_cascade_ ));
    CascadeMux I__1185 (
            .O(N__10132),
            .I(\receive_module.n4212_cascade_ ));
    CascadeMux I__1184 (
            .O(N__10129),
            .I(\receive_module.n4213_cascade_ ));
    InMux I__1183 (
            .O(N__10126),
            .I(N__10123));
    LocalMux I__1182 (
            .O(N__10123),
            .I(\receive_module.rx_counter.n3204 ));
    SRMux I__1181 (
            .O(N__10120),
            .I(N__10117));
    LocalMux I__1180 (
            .O(N__10117),
            .I(N__10114));
    Span4Mux_v I__1179 (
            .O(N__10114),
            .I(N__10109));
    SRMux I__1178 (
            .O(N__10113),
            .I(N__10106));
    SRMux I__1177 (
            .O(N__10112),
            .I(N__10102));
    Span4Mux_v I__1176 (
            .O(N__10109),
            .I(N__10099));
    LocalMux I__1175 (
            .O(N__10106),
            .I(N__10096));
    SRMux I__1174 (
            .O(N__10105),
            .I(N__10093));
    LocalMux I__1173 (
            .O(N__10102),
            .I(N__10090));
    Span4Mux_v I__1172 (
            .O(N__10099),
            .I(N__10083));
    Span4Mux_v I__1171 (
            .O(N__10096),
            .I(N__10083));
    LocalMux I__1170 (
            .O(N__10093),
            .I(N__10083));
    Span4Mux_h I__1169 (
            .O(N__10090),
            .I(N__10078));
    Span4Mux_h I__1168 (
            .O(N__10083),
            .I(N__10078));
    Odrv4 I__1167 (
            .O(N__10078),
            .I(n659));
    IoInMux I__1166 (
            .O(N__10075),
            .I(N__10072));
    LocalMux I__1165 (
            .O(N__10072),
            .I(N__10069));
    Span4Mux_s3_h I__1164 (
            .O(N__10069),
            .I(N__10066));
    Span4Mux_v I__1163 (
            .O(N__10066),
            .I(N__10063));
    Span4Mux_h I__1162 (
            .O(N__10063),
            .I(N__10060));
    Span4Mux_h I__1161 (
            .O(N__10060),
            .I(N__10057));
    Odrv4 I__1160 (
            .O(N__10057),
            .I(DEBUG_c_0));
    IoInMux I__1159 (
            .O(N__10054),
            .I(N__10051));
    LocalMux I__1158 (
            .O(N__10051),
            .I(N__10048));
    IoSpan4Mux I__1157 (
            .O(N__10048),
            .I(N__10044));
    IoInMux I__1156 (
            .O(N__10047),
            .I(N__10041));
    Span4Mux_s1_v I__1155 (
            .O(N__10044),
            .I(N__10037));
    LocalMux I__1154 (
            .O(N__10041),
            .I(N__10034));
    IoInMux I__1153 (
            .O(N__10040),
            .I(N__10031));
    Span4Mux_v I__1152 (
            .O(N__10037),
            .I(N__10026));
    Span4Mux_s2_h I__1151 (
            .O(N__10034),
            .I(N__10026));
    LocalMux I__1150 (
            .O(N__10031),
            .I(N__10023));
    Span4Mux_h I__1149 (
            .O(N__10026),
            .I(N__10020));
    Span4Mux_s1_v I__1148 (
            .O(N__10023),
            .I(N__10017));
    Span4Mux_h I__1147 (
            .O(N__10020),
            .I(N__10012));
    Span4Mux_v I__1146 (
            .O(N__10017),
            .I(N__10012));
    Span4Mux_v I__1145 (
            .O(N__10012),
            .I(N__10009));
    Odrv4 I__1144 (
            .O(N__10009),
            .I(n1996));
    InMux I__1143 (
            .O(N__10006),
            .I(N__10003));
    LocalMux I__1142 (
            .O(N__10003),
            .I(\transmit_module.Y_DELTA_PATTERN_70 ));
    InMux I__1141 (
            .O(N__10000),
            .I(N__9997));
    LocalMux I__1140 (
            .O(N__9997),
            .I(N__9994));
    Odrv4 I__1139 (
            .O(N__9994),
            .I(\transmit_module.Y_DELTA_PATTERN_72 ));
    InMux I__1138 (
            .O(N__9991),
            .I(N__9988));
    LocalMux I__1137 (
            .O(N__9988),
            .I(\transmit_module.Y_DELTA_PATTERN_71 ));
    InMux I__1136 (
            .O(N__9985),
            .I(N__9982));
    LocalMux I__1135 (
            .O(N__9982),
            .I(\transmit_module.Y_DELTA_PATTERN_63 ));
    CascadeMux I__1134 (
            .O(N__9979),
            .I(N__9976));
    CascadeBuf I__1133 (
            .O(N__9976),
            .I(N__9972));
    CascadeMux I__1132 (
            .O(N__9975),
            .I(N__9969));
    CascadeMux I__1131 (
            .O(N__9972),
            .I(N__9966));
    CascadeBuf I__1130 (
            .O(N__9969),
            .I(N__9963));
    CascadeBuf I__1129 (
            .O(N__9966),
            .I(N__9960));
    CascadeMux I__1128 (
            .O(N__9963),
            .I(N__9957));
    CascadeMux I__1127 (
            .O(N__9960),
            .I(N__9954));
    CascadeBuf I__1126 (
            .O(N__9957),
            .I(N__9951));
    CascadeBuf I__1125 (
            .O(N__9954),
            .I(N__9948));
    CascadeMux I__1124 (
            .O(N__9951),
            .I(N__9945));
    CascadeMux I__1123 (
            .O(N__9948),
            .I(N__9942));
    CascadeBuf I__1122 (
            .O(N__9945),
            .I(N__9939));
    CascadeBuf I__1121 (
            .O(N__9942),
            .I(N__9936));
    CascadeMux I__1120 (
            .O(N__9939),
            .I(N__9933));
    CascadeMux I__1119 (
            .O(N__9936),
            .I(N__9930));
    CascadeBuf I__1118 (
            .O(N__9933),
            .I(N__9927));
    CascadeBuf I__1117 (
            .O(N__9930),
            .I(N__9924));
    CascadeMux I__1116 (
            .O(N__9927),
            .I(N__9921));
    CascadeMux I__1115 (
            .O(N__9924),
            .I(N__9918));
    CascadeBuf I__1114 (
            .O(N__9921),
            .I(N__9915));
    CascadeBuf I__1113 (
            .O(N__9918),
            .I(N__9912));
    CascadeMux I__1112 (
            .O(N__9915),
            .I(N__9909));
    CascadeMux I__1111 (
            .O(N__9912),
            .I(N__9906));
    CascadeBuf I__1110 (
            .O(N__9909),
            .I(N__9903));
    CascadeBuf I__1109 (
            .O(N__9906),
            .I(N__9900));
    CascadeMux I__1108 (
            .O(N__9903),
            .I(N__9897));
    CascadeMux I__1107 (
            .O(N__9900),
            .I(N__9894));
    CascadeBuf I__1106 (
            .O(N__9897),
            .I(N__9891));
    CascadeBuf I__1105 (
            .O(N__9894),
            .I(N__9888));
    CascadeMux I__1104 (
            .O(N__9891),
            .I(N__9885));
    CascadeMux I__1103 (
            .O(N__9888),
            .I(N__9882));
    CascadeBuf I__1102 (
            .O(N__9885),
            .I(N__9879));
    CascadeBuf I__1101 (
            .O(N__9882),
            .I(N__9876));
    CascadeMux I__1100 (
            .O(N__9879),
            .I(N__9873));
    CascadeMux I__1099 (
            .O(N__9876),
            .I(N__9870));
    CascadeBuf I__1098 (
            .O(N__9873),
            .I(N__9867));
    CascadeBuf I__1097 (
            .O(N__9870),
            .I(N__9864));
    CascadeMux I__1096 (
            .O(N__9867),
            .I(N__9861));
    CascadeMux I__1095 (
            .O(N__9864),
            .I(N__9858));
    CascadeBuf I__1094 (
            .O(N__9861),
            .I(N__9855));
    CascadeBuf I__1093 (
            .O(N__9858),
            .I(N__9852));
    CascadeMux I__1092 (
            .O(N__9855),
            .I(N__9849));
    CascadeMux I__1091 (
            .O(N__9852),
            .I(N__9846));
    CascadeBuf I__1090 (
            .O(N__9849),
            .I(N__9843));
    CascadeBuf I__1089 (
            .O(N__9846),
            .I(N__9840));
    CascadeMux I__1088 (
            .O(N__9843),
            .I(N__9837));
    CascadeMux I__1087 (
            .O(N__9840),
            .I(N__9834));
    CascadeBuf I__1086 (
            .O(N__9837),
            .I(N__9831));
    CascadeBuf I__1085 (
            .O(N__9834),
            .I(N__9828));
    CascadeMux I__1084 (
            .O(N__9831),
            .I(N__9825));
    CascadeMux I__1083 (
            .O(N__9828),
            .I(N__9822));
    CascadeBuf I__1082 (
            .O(N__9825),
            .I(N__9819));
    CascadeBuf I__1081 (
            .O(N__9822),
            .I(N__9816));
    CascadeMux I__1080 (
            .O(N__9819),
            .I(N__9813));
    CascadeMux I__1079 (
            .O(N__9816),
            .I(N__9810));
    CascadeBuf I__1078 (
            .O(N__9813),
            .I(N__9807));
    CascadeBuf I__1077 (
            .O(N__9810),
            .I(N__9804));
    CascadeMux I__1076 (
            .O(N__9807),
            .I(N__9801));
    CascadeMux I__1075 (
            .O(N__9804),
            .I(N__9798));
    CascadeBuf I__1074 (
            .O(N__9801),
            .I(N__9795));
    InMux I__1073 (
            .O(N__9798),
            .I(N__9792));
    CascadeMux I__1072 (
            .O(N__9795),
            .I(N__9789));
    LocalMux I__1071 (
            .O(N__9792),
            .I(N__9786));
    InMux I__1070 (
            .O(N__9789),
            .I(N__9783));
    Span12Mux_h I__1069 (
            .O(N__9786),
            .I(N__9780));
    LocalMux I__1068 (
            .O(N__9783),
            .I(N__9777));
    Odrv12 I__1067 (
            .O(N__9780),
            .I(n18));
    Odrv4 I__1066 (
            .O(N__9777),
            .I(n18));
    SRMux I__1065 (
            .O(N__9772),
            .I(N__9769));
    LocalMux I__1064 (
            .O(N__9769),
            .I(N__9765));
    SRMux I__1063 (
            .O(N__9768),
            .I(N__9762));
    Span4Mux_v I__1062 (
            .O(N__9765),
            .I(N__9757));
    LocalMux I__1061 (
            .O(N__9762),
            .I(N__9757));
    Span4Mux_h I__1060 (
            .O(N__9757),
            .I(N__9754));
    Sp12to4 I__1059 (
            .O(N__9754),
            .I(N__9751));
    Odrv12 I__1058 (
            .O(N__9751),
            .I(\receive_module.rx_counter.PULSE_1HZ_N_97 ));
    CascadeMux I__1057 (
            .O(N__9748),
            .I(\transmit_module.video_signal_controller.n3935_cascade_ ));
    InMux I__1056 (
            .O(N__9745),
            .I(N__9742));
    LocalMux I__1055 (
            .O(N__9742),
            .I(\transmit_module.video_signal_controller.n6 ));
    InMux I__1054 (
            .O(N__9739),
            .I(N__9736));
    LocalMux I__1053 (
            .O(N__9736),
            .I(\transmit_module.Y_DELTA_PATTERN_98 ));
    InMux I__1052 (
            .O(N__9733),
            .I(N__9730));
    LocalMux I__1051 (
            .O(N__9730),
            .I(\transmit_module.Y_DELTA_PATTERN_76 ));
    InMux I__1050 (
            .O(N__9727),
            .I(N__9724));
    LocalMux I__1049 (
            .O(N__9724),
            .I(\transmit_module.Y_DELTA_PATTERN_73 ));
    InMux I__1048 (
            .O(N__9721),
            .I(N__9718));
    LocalMux I__1047 (
            .O(N__9718),
            .I(N__9715));
    Span4Mux_v I__1046 (
            .O(N__9715),
            .I(N__9712));
    Odrv4 I__1045 (
            .O(N__9712),
            .I(\transmit_module.Y_DELTA_PATTERN_82 ));
    InMux I__1044 (
            .O(N__9709),
            .I(N__9706));
    LocalMux I__1043 (
            .O(N__9706),
            .I(\transmit_module.Y_DELTA_PATTERN_75 ));
    InMux I__1042 (
            .O(N__9703),
            .I(N__9700));
    LocalMux I__1041 (
            .O(N__9700),
            .I(\transmit_module.Y_DELTA_PATTERN_74 ));
    InMux I__1040 (
            .O(N__9697),
            .I(N__9694));
    LocalMux I__1039 (
            .O(N__9694),
            .I(\transmit_module.Y_DELTA_PATTERN_77 ));
    CascadeMux I__1038 (
            .O(N__9691),
            .I(N__9688));
    InMux I__1037 (
            .O(N__9688),
            .I(N__9685));
    LocalMux I__1036 (
            .O(N__9685),
            .I(N__9682));
    Odrv4 I__1035 (
            .O(N__9682),
            .I(\receive_module.rx_counter.n3979 ));
    InMux I__1034 (
            .O(N__9679),
            .I(\receive_module.rx_counter.O_VISIBLE_N_89 ));
    IoInMux I__1033 (
            .O(N__9676),
            .I(N__9673));
    LocalMux I__1032 (
            .O(N__9673),
            .I(N__9669));
    InMux I__1031 (
            .O(N__9672),
            .I(N__9666));
    Span4Mux_s1_h I__1030 (
            .O(N__9669),
            .I(N__9663));
    LocalMux I__1029 (
            .O(N__9666),
            .I(N__9660));
    Sp12to4 I__1028 (
            .O(N__9663),
            .I(N__9657));
    Span4Mux_h I__1027 (
            .O(N__9660),
            .I(N__9654));
    Span12Mux_v I__1026 (
            .O(N__9657),
            .I(N__9651));
    Sp12to4 I__1025 (
            .O(N__9654),
            .I(N__9648));
    Odrv12 I__1024 (
            .O(N__9651),
            .I(DEBUG_c_6));
    Odrv12 I__1023 (
            .O(N__9648),
            .I(DEBUG_c_6));
    InMux I__1022 (
            .O(N__9643),
            .I(N__9640));
    LocalMux I__1021 (
            .O(N__9640),
            .I(\transmit_module.video_signal_controller.SYNC_BUFF1 ));
    CascadeMux I__1020 (
            .O(N__9637),
            .I(\transmit_module.video_signal_controller.n3987_cascade_ ));
    CascadeMux I__1019 (
            .O(N__9634),
            .I(\transmit_module.video_signal_controller.n4_cascade_ ));
    InMux I__1018 (
            .O(N__9631),
            .I(N__9628));
    LocalMux I__1017 (
            .O(N__9628),
            .I(\transmit_module.video_signal_controller.n3935 ));
    CascadeMux I__1016 (
            .O(N__9625),
            .I(N__9622));
    InMux I__1015 (
            .O(N__9622),
            .I(N__9616));
    InMux I__1014 (
            .O(N__9621),
            .I(N__9613));
    InMux I__1013 (
            .O(N__9620),
            .I(N__9610));
    InMux I__1012 (
            .O(N__9619),
            .I(N__9607));
    LocalMux I__1011 (
            .O(N__9616),
            .I(\receive_module.rx_counter.Y_1 ));
    LocalMux I__1010 (
            .O(N__9613),
            .I(\receive_module.rx_counter.Y_1 ));
    LocalMux I__1009 (
            .O(N__9610),
            .I(\receive_module.rx_counter.Y_1 ));
    LocalMux I__1008 (
            .O(N__9607),
            .I(\receive_module.rx_counter.Y_1 ));
    InMux I__1007 (
            .O(N__9598),
            .I(\receive_module.rx_counter.n3711 ));
    CascadeMux I__1006 (
            .O(N__9595),
            .I(N__9589));
    InMux I__1005 (
            .O(N__9594),
            .I(N__9586));
    InMux I__1004 (
            .O(N__9593),
            .I(N__9583));
    InMux I__1003 (
            .O(N__9592),
            .I(N__9580));
    InMux I__1002 (
            .O(N__9589),
            .I(N__9577));
    LocalMux I__1001 (
            .O(N__9586),
            .I(\receive_module.rx_counter.Y_2 ));
    LocalMux I__1000 (
            .O(N__9583),
            .I(\receive_module.rx_counter.Y_2 ));
    LocalMux I__999 (
            .O(N__9580),
            .I(\receive_module.rx_counter.Y_2 ));
    LocalMux I__998 (
            .O(N__9577),
            .I(\receive_module.rx_counter.Y_2 ));
    InMux I__997 (
            .O(N__9568),
            .I(\receive_module.rx_counter.n3712 ));
    InMux I__996 (
            .O(N__9565),
            .I(N__9559));
    InMux I__995 (
            .O(N__9564),
            .I(N__9556));
    InMux I__994 (
            .O(N__9563),
            .I(N__9553));
    InMux I__993 (
            .O(N__9562),
            .I(N__9550));
    LocalMux I__992 (
            .O(N__9559),
            .I(\receive_module.rx_counter.Y_3 ));
    LocalMux I__991 (
            .O(N__9556),
            .I(\receive_module.rx_counter.Y_3 ));
    LocalMux I__990 (
            .O(N__9553),
            .I(\receive_module.rx_counter.Y_3 ));
    LocalMux I__989 (
            .O(N__9550),
            .I(\receive_module.rx_counter.Y_3 ));
    InMux I__988 (
            .O(N__9541),
            .I(\receive_module.rx_counter.n3713 ));
    InMux I__987 (
            .O(N__9538),
            .I(N__9532));
    InMux I__986 (
            .O(N__9537),
            .I(N__9527));
    InMux I__985 (
            .O(N__9536),
            .I(N__9527));
    InMux I__984 (
            .O(N__9535),
            .I(N__9524));
    LocalMux I__983 (
            .O(N__9532),
            .I(\receive_module.rx_counter.Y_4 ));
    LocalMux I__982 (
            .O(N__9527),
            .I(\receive_module.rx_counter.Y_4 ));
    LocalMux I__981 (
            .O(N__9524),
            .I(\receive_module.rx_counter.Y_4 ));
    InMux I__980 (
            .O(N__9517),
            .I(\receive_module.rx_counter.n3714 ));
    InMux I__979 (
            .O(N__9514),
            .I(N__9509));
    InMux I__978 (
            .O(N__9513),
            .I(N__9506));
    InMux I__977 (
            .O(N__9512),
            .I(N__9503));
    LocalMux I__976 (
            .O(N__9509),
            .I(\receive_module.rx_counter.Y_5 ));
    LocalMux I__975 (
            .O(N__9506),
            .I(\receive_module.rx_counter.Y_5 ));
    LocalMux I__974 (
            .O(N__9503),
            .I(\receive_module.rx_counter.Y_5 ));
    InMux I__973 (
            .O(N__9496),
            .I(\receive_module.rx_counter.n3715 ));
    CascadeMux I__972 (
            .O(N__9493),
            .I(N__9489));
    InMux I__971 (
            .O(N__9492),
            .I(N__9485));
    InMux I__970 (
            .O(N__9489),
            .I(N__9482));
    InMux I__969 (
            .O(N__9488),
            .I(N__9479));
    LocalMux I__968 (
            .O(N__9485),
            .I(\receive_module.rx_counter.Y_6 ));
    LocalMux I__967 (
            .O(N__9482),
            .I(\receive_module.rx_counter.Y_6 ));
    LocalMux I__966 (
            .O(N__9479),
            .I(\receive_module.rx_counter.Y_6 ));
    InMux I__965 (
            .O(N__9472),
            .I(\receive_module.rx_counter.n3716 ));
    InMux I__964 (
            .O(N__9469),
            .I(N__9463));
    InMux I__963 (
            .O(N__9468),
            .I(N__9458));
    InMux I__962 (
            .O(N__9467),
            .I(N__9458));
    InMux I__961 (
            .O(N__9466),
            .I(N__9455));
    LocalMux I__960 (
            .O(N__9463),
            .I(\receive_module.rx_counter.Y_7 ));
    LocalMux I__959 (
            .O(N__9458),
            .I(\receive_module.rx_counter.Y_7 ));
    LocalMux I__958 (
            .O(N__9455),
            .I(\receive_module.rx_counter.Y_7 ));
    InMux I__957 (
            .O(N__9448),
            .I(\receive_module.rx_counter.n3717 ));
    InMux I__956 (
            .O(N__9445),
            .I(N__9439));
    InMux I__955 (
            .O(N__9444),
            .I(N__9436));
    InMux I__954 (
            .O(N__9443),
            .I(N__9433));
    InMux I__953 (
            .O(N__9442),
            .I(N__9430));
    LocalMux I__952 (
            .O(N__9439),
            .I(\receive_module.rx_counter.Y_8 ));
    LocalMux I__951 (
            .O(N__9436),
            .I(\receive_module.rx_counter.Y_8 ));
    LocalMux I__950 (
            .O(N__9433),
            .I(\receive_module.rx_counter.Y_8 ));
    LocalMux I__949 (
            .O(N__9430),
            .I(\receive_module.rx_counter.Y_8 ));
    InMux I__948 (
            .O(N__9421),
            .I(N__9418));
    LocalMux I__947 (
            .O(N__9418),
            .I(\transmit_module.Y_DELTA_PATTERN_89 ));
    InMux I__946 (
            .O(N__9415),
            .I(N__9412));
    LocalMux I__945 (
            .O(N__9412),
            .I(\transmit_module.Y_DELTA_PATTERN_88 ));
    InMux I__944 (
            .O(N__9409),
            .I(N__9406));
    LocalMux I__943 (
            .O(N__9406),
            .I(\transmit_module.Y_DELTA_PATTERN_87 ));
    InMux I__942 (
            .O(N__9403),
            .I(N__9400));
    LocalMux I__941 (
            .O(N__9400),
            .I(\transmit_module.Y_DELTA_PATTERN_92 ));
    InMux I__940 (
            .O(N__9397),
            .I(N__9394));
    LocalMux I__939 (
            .O(N__9394),
            .I(\transmit_module.Y_DELTA_PATTERN_91 ));
    InMux I__938 (
            .O(N__9391),
            .I(N__9388));
    LocalMux I__937 (
            .O(N__9388),
            .I(\transmit_module.Y_DELTA_PATTERN_86 ));
    InMux I__936 (
            .O(N__9385),
            .I(N__9382));
    LocalMux I__935 (
            .O(N__9382),
            .I(N__9379));
    Odrv4 I__934 (
            .O(N__9379),
            .I(\transmit_module.Y_DELTA_PATTERN_85 ));
    InMux I__933 (
            .O(N__9376),
            .I(N__9373));
    LocalMux I__932 (
            .O(N__9373),
            .I(\transmit_module.Y_DELTA_PATTERN_94 ));
    InMux I__931 (
            .O(N__9370),
            .I(N__9367));
    LocalMux I__930 (
            .O(N__9367),
            .I(\transmit_module.Y_DELTA_PATTERN_93 ));
    InMux I__929 (
            .O(N__9364),
            .I(N__9361));
    LocalMux I__928 (
            .O(N__9361),
            .I(\transmit_module.Y_DELTA_PATTERN_96 ));
    InMux I__927 (
            .O(N__9358),
            .I(N__9355));
    LocalMux I__926 (
            .O(N__9355),
            .I(\transmit_module.Y_DELTA_PATTERN_97 ));
    InMux I__925 (
            .O(N__9352),
            .I(N__9349));
    LocalMux I__924 (
            .O(N__9349),
            .I(N__9346));
    Odrv4 I__923 (
            .O(N__9346),
            .I(\line_buffer.n624 ));
    InMux I__922 (
            .O(N__9343),
            .I(N__9340));
    LocalMux I__921 (
            .O(N__9340),
            .I(\line_buffer.n4122 ));
    CascadeMux I__920 (
            .O(N__9337),
            .I(N__9334));
    InMux I__919 (
            .O(N__9334),
            .I(N__9331));
    LocalMux I__918 (
            .O(N__9331),
            .I(N__9328));
    Span4Mux_h I__917 (
            .O(N__9328),
            .I(N__9325));
    Span4Mux_h I__916 (
            .O(N__9325),
            .I(N__9322));
    Sp12to4 I__915 (
            .O(N__9322),
            .I(N__9319));
    Span12Mux_v I__914 (
            .O(N__9319),
            .I(N__9316));
    Span12Mux_v I__913 (
            .O(N__9316),
            .I(N__9313));
    Odrv12 I__912 (
            .O(N__9313),
            .I(\line_buffer.n616 ));
    InMux I__911 (
            .O(N__9310),
            .I(N__9304));
    InMux I__910 (
            .O(N__9309),
            .I(N__9301));
    InMux I__909 (
            .O(N__9308),
            .I(N__9298));
    InMux I__908 (
            .O(N__9307),
            .I(N__9295));
    LocalMux I__907 (
            .O(N__9304),
            .I(\receive_module.rx_counter.Y_0 ));
    LocalMux I__906 (
            .O(N__9301),
            .I(\receive_module.rx_counter.Y_0 ));
    LocalMux I__905 (
            .O(N__9298),
            .I(\receive_module.rx_counter.Y_0 ));
    LocalMux I__904 (
            .O(N__9295),
            .I(\receive_module.rx_counter.Y_0 ));
    InMux I__903 (
            .O(N__9286),
            .I(bfn_11_9_0_));
    InMux I__902 (
            .O(N__9283),
            .I(\receive_module.rx_counter.n3674 ));
    InMux I__901 (
            .O(N__9280),
            .I(\receive_module.rx_counter.n3675 ));
    InMux I__900 (
            .O(N__9277),
            .I(bfn_10_10_0_));
    InMux I__899 (
            .O(N__9274),
            .I(N__9271));
    LocalMux I__898 (
            .O(N__9271),
            .I(\transmit_module.Y_DELTA_PATTERN_84 ));
    InMux I__897 (
            .O(N__9268),
            .I(N__9265));
    LocalMux I__896 (
            .O(N__9265),
            .I(\transmit_module.Y_DELTA_PATTERN_83 ));
    InMux I__895 (
            .O(N__9262),
            .I(N__9259));
    LocalMux I__894 (
            .O(N__9259),
            .I(\transmit_module.Y_DELTA_PATTERN_90 ));
    InMux I__893 (
            .O(N__9256),
            .I(N__9253));
    LocalMux I__892 (
            .O(N__9253),
            .I(\transmit_module.Y_DELTA_PATTERN_95 ));
    InMux I__891 (
            .O(N__9250),
            .I(N__9247));
    LocalMux I__890 (
            .O(N__9247),
            .I(N__9244));
    Span4Mux_v I__889 (
            .O(N__9244),
            .I(N__9241));
    Odrv4 I__888 (
            .O(N__9241),
            .I(\line_buffer.n680 ));
    CascadeMux I__887 (
            .O(N__9238),
            .I(N__9235));
    InMux I__886 (
            .O(N__9235),
            .I(N__9232));
    LocalMux I__885 (
            .O(N__9232),
            .I(N__9229));
    Span4Mux_h I__884 (
            .O(N__9229),
            .I(N__9226));
    Odrv4 I__883 (
            .O(N__9226),
            .I(\line_buffer.n688 ));
    InMux I__882 (
            .O(N__9223),
            .I(bfn_10_9_0_));
    InMux I__881 (
            .O(N__9220),
            .I(\receive_module.rx_counter.n3669 ));
    InMux I__880 (
            .O(N__9217),
            .I(\receive_module.rx_counter.n3670 ));
    InMux I__879 (
            .O(N__9214),
            .I(\receive_module.rx_counter.n3671 ));
    InMux I__878 (
            .O(N__9211),
            .I(\receive_module.rx_counter.n3672 ));
    InMux I__877 (
            .O(N__9208),
            .I(\receive_module.rx_counter.n3673 ));
    CascadeMux I__876 (
            .O(N__9205),
            .I(\receive_module.rx_counter.n3176_cascade_ ));
    InMux I__875 (
            .O(N__9202),
            .I(N__9199));
    LocalMux I__874 (
            .O(N__9199),
            .I(\receive_module.rx_counter.n3208 ));
    InMux I__873 (
            .O(N__9196),
            .I(N__9193));
    LocalMux I__872 (
            .O(N__9193),
            .I(N__9190));
    Span4Mux_v I__871 (
            .O(N__9190),
            .I(N__9187));
    Sp12to4 I__870 (
            .O(N__9187),
            .I(N__9184));
    Span12Mux_h I__869 (
            .O(N__9184),
            .I(N__9181));
    Span12Mux_v I__868 (
            .O(N__9181),
            .I(N__9178));
    Odrv12 I__867 (
            .O(N__9178),
            .I(\line_buffer.n675 ));
    InMux I__866 (
            .O(N__9175),
            .I(N__9172));
    LocalMux I__865 (
            .O(N__9172),
            .I(N__9169));
    Odrv4 I__864 (
            .O(N__9169),
            .I(\line_buffer.n683 ));
    InMux I__863 (
            .O(N__9166),
            .I(N__9163));
    LocalMux I__862 (
            .O(N__9163),
            .I(N__9160));
    Span4Mux_v I__861 (
            .O(N__9160),
            .I(N__9157));
    Span4Mux_h I__860 (
            .O(N__9157),
            .I(N__9154));
    Sp12to4 I__859 (
            .O(N__9154),
            .I(N__9151));
    Span12Mux_h I__858 (
            .O(N__9151),
            .I(N__9148));
    Odrv12 I__857 (
            .O(N__9148),
            .I(\line_buffer.n611 ));
    CascadeMux I__856 (
            .O(N__9145),
            .I(\line_buffer.n4170_cascade_ ));
    InMux I__855 (
            .O(N__9142),
            .I(N__9139));
    LocalMux I__854 (
            .O(N__9139),
            .I(N__9136));
    Span4Mux_v I__853 (
            .O(N__9136),
            .I(N__9133));
    Span4Mux_v I__852 (
            .O(N__9133),
            .I(N__9130));
    Odrv4 I__851 (
            .O(N__9130),
            .I(\line_buffer.n619 ));
    InMux I__850 (
            .O(N__9127),
            .I(N__9124));
    LocalMux I__849 (
            .O(N__9124),
            .I(N__9121));
    Span4Mux_v I__848 (
            .O(N__9121),
            .I(N__9118));
    Sp12to4 I__847 (
            .O(N__9118),
            .I(N__9115));
    Span12Mux_h I__846 (
            .O(N__9115),
            .I(N__9112));
    Odrv12 I__845 (
            .O(N__9112),
            .I(\line_buffer.n643 ));
    CascadeMux I__844 (
            .O(N__9109),
            .I(N__9106));
    InMux I__843 (
            .O(N__9106),
            .I(N__9103));
    LocalMux I__842 (
            .O(N__9103),
            .I(N__9100));
    Span4Mux_v I__841 (
            .O(N__9100),
            .I(N__9097));
    Odrv4 I__840 (
            .O(N__9097),
            .I(\line_buffer.n651 ));
    InMux I__839 (
            .O(N__9094),
            .I(N__9091));
    LocalMux I__838 (
            .O(N__9091),
            .I(N__9088));
    Span4Mux_v I__837 (
            .O(N__9088),
            .I(N__9085));
    Span4Mux_v I__836 (
            .O(N__9085),
            .I(N__9082));
    Odrv4 I__835 (
            .O(N__9082),
            .I(\line_buffer.n687 ));
    InMux I__834 (
            .O(N__9079),
            .I(N__9076));
    LocalMux I__833 (
            .O(N__9076),
            .I(\line_buffer.n679 ));
    InMux I__832 (
            .O(N__9073),
            .I(N__9070));
    LocalMux I__831 (
            .O(N__9070),
            .I(\line_buffer.n4152 ));
    InMux I__830 (
            .O(N__9067),
            .I(N__9064));
    LocalMux I__829 (
            .O(N__9064),
            .I(N__9061));
    Span4Mux_h I__828 (
            .O(N__9061),
            .I(N__9058));
    Sp12to4 I__827 (
            .O(N__9058),
            .I(N__9055));
    Span12Mux_v I__826 (
            .O(N__9055),
            .I(N__9052));
    Span12Mux_h I__825 (
            .O(N__9052),
            .I(N__9049));
    Odrv12 I__824 (
            .O(N__9049),
            .I(\line_buffer.n554 ));
    CascadeMux I__823 (
            .O(N__9046),
            .I(N__9043));
    InMux I__822 (
            .O(N__9043),
            .I(N__9040));
    LocalMux I__821 (
            .O(N__9040),
            .I(N__9037));
    Span4Mux_h I__820 (
            .O(N__9037),
            .I(N__9034));
    Sp12to4 I__819 (
            .O(N__9034),
            .I(N__9031));
    Span12Mux_v I__818 (
            .O(N__9031),
            .I(N__9028));
    Odrv12 I__817 (
            .O(N__9028),
            .I(\line_buffer.n546 ));
    CascadeMux I__816 (
            .O(N__9025),
            .I(\line_buffer.n4155_cascade_ ));
    InMux I__815 (
            .O(N__9022),
            .I(N__9019));
    LocalMux I__814 (
            .O(N__9019),
            .I(\line_buffer.n4173 ));
    InMux I__813 (
            .O(N__9016),
            .I(N__9013));
    LocalMux I__812 (
            .O(N__9013),
            .I(N__9010));
    Span4Mux_s2_v I__811 (
            .O(N__9010),
            .I(N__9006));
    InMux I__810 (
            .O(N__9009),
            .I(N__9003));
    Span4Mux_v I__809 (
            .O(N__9006),
            .I(N__8998));
    LocalMux I__808 (
            .O(N__9003),
            .I(N__8998));
    Span4Mux_v I__807 (
            .O(N__8998),
            .I(N__8994));
    InMux I__806 (
            .O(N__8997),
            .I(N__8991));
    Span4Mux_v I__805 (
            .O(N__8994),
            .I(N__8985));
    LocalMux I__804 (
            .O(N__8991),
            .I(N__8985));
    InMux I__803 (
            .O(N__8990),
            .I(N__8982));
    Span4Mux_v I__802 (
            .O(N__8985),
            .I(N__8979));
    LocalMux I__801 (
            .O(N__8982),
            .I(N__8976));
    Span4Mux_v I__800 (
            .O(N__8979),
            .I(N__8969));
    Span4Mux_v I__799 (
            .O(N__8976),
            .I(N__8969));
    InMux I__798 (
            .O(N__8975),
            .I(N__8966));
    InMux I__797 (
            .O(N__8974),
            .I(N__8963));
    Span4Mux_v I__796 (
            .O(N__8969),
            .I(N__8958));
    LocalMux I__795 (
            .O(N__8966),
            .I(N__8958));
    LocalMux I__794 (
            .O(N__8963),
            .I(N__8955));
    Span4Mux_h I__793 (
            .O(N__8958),
            .I(N__8951));
    Span4Mux_h I__792 (
            .O(N__8955),
            .I(N__8948));
    InMux I__791 (
            .O(N__8954),
            .I(N__8945));
    Span4Mux_h I__790 (
            .O(N__8951),
            .I(N__8942));
    Span4Mux_v I__789 (
            .O(N__8948),
            .I(N__8938));
    LocalMux I__788 (
            .O(N__8945),
            .I(N__8935));
    Span4Mux_h I__787 (
            .O(N__8942),
            .I(N__8932));
    InMux I__786 (
            .O(N__8941),
            .I(N__8929));
    Span4Mux_v I__785 (
            .O(N__8938),
            .I(N__8924));
    Span4Mux_h I__784 (
            .O(N__8935),
            .I(N__8924));
    Span4Mux_h I__783 (
            .O(N__8932),
            .I(N__8919));
    LocalMux I__782 (
            .O(N__8929),
            .I(N__8919));
    Span4Mux_v I__781 (
            .O(N__8924),
            .I(N__8916));
    Span4Mux_h I__780 (
            .O(N__8919),
            .I(N__8913));
    Span4Mux_v I__779 (
            .O(N__8916),
            .I(N__8910));
    Span4Mux_v I__778 (
            .O(N__8913),
            .I(N__8907));
    Odrv4 I__777 (
            .O(N__8910),
            .I(TVP_VIDEO_c_2));
    Odrv4 I__776 (
            .O(N__8907),
            .I(TVP_VIDEO_c_2));
    CascadeMux I__775 (
            .O(N__8902),
            .I(\receive_module.rx_counter.n12_cascade_ ));
    CascadeMux I__774 (
            .O(N__8899),
            .I(\receive_module.rx_counter.n3938_cascade_ ));
    InMux I__773 (
            .O(N__8896),
            .I(N__8893));
    LocalMux I__772 (
            .O(N__8893),
            .I(\receive_module.rx_counter.n3938 ));
    InMux I__771 (
            .O(N__8890),
            .I(N__8887));
    LocalMux I__770 (
            .O(N__8887),
            .I(\receive_module.rx_counter.n13 ));
    InMux I__769 (
            .O(N__8884),
            .I(N__8880));
    InMux I__768 (
            .O(N__8883),
            .I(N__8877));
    LocalMux I__767 (
            .O(N__8880),
            .I(N__8870));
    LocalMux I__766 (
            .O(N__8877),
            .I(N__8870));
    InMux I__765 (
            .O(N__8876),
            .I(N__8867));
    InMux I__764 (
            .O(N__8875),
            .I(N__8864));
    Span4Mux_v I__763 (
            .O(N__8870),
            .I(N__8857));
    LocalMux I__762 (
            .O(N__8867),
            .I(N__8857));
    LocalMux I__761 (
            .O(N__8864),
            .I(N__8857));
    Span4Mux_v I__760 (
            .O(N__8857),
            .I(N__8852));
    InMux I__759 (
            .O(N__8856),
            .I(N__8849));
    InMux I__758 (
            .O(N__8855),
            .I(N__8846));
    Span4Mux_v I__757 (
            .O(N__8852),
            .I(N__8841));
    LocalMux I__756 (
            .O(N__8849),
            .I(N__8841));
    LocalMux I__755 (
            .O(N__8846),
            .I(N__8836));
    Span4Mux_h I__754 (
            .O(N__8841),
            .I(N__8833));
    InMux I__753 (
            .O(N__8840),
            .I(N__8830));
    InMux I__752 (
            .O(N__8839),
            .I(N__8827));
    Span4Mux_v I__751 (
            .O(N__8836),
            .I(N__8824));
    Span4Mux_h I__750 (
            .O(N__8833),
            .I(N__8821));
    LocalMux I__749 (
            .O(N__8830),
            .I(N__8818));
    LocalMux I__748 (
            .O(N__8827),
            .I(N__8815));
    Sp12to4 I__747 (
            .O(N__8824),
            .I(N__8812));
    Span4Mux_v I__746 (
            .O(N__8821),
            .I(N__8809));
    Span4Mux_h I__745 (
            .O(N__8818),
            .I(N__8806));
    Span4Mux_h I__744 (
            .O(N__8815),
            .I(N__8803));
    Span12Mux_h I__743 (
            .O(N__8812),
            .I(N__8800));
    Span4Mux_v I__742 (
            .O(N__8809),
            .I(N__8797));
    Span4Mux_h I__741 (
            .O(N__8806),
            .I(N__8794));
    Span4Mux_h I__740 (
            .O(N__8803),
            .I(N__8791));
    Span12Mux_v I__739 (
            .O(N__8800),
            .I(N__8788));
    Span4Mux_v I__738 (
            .O(N__8797),
            .I(N__8783));
    Span4Mux_h I__737 (
            .O(N__8794),
            .I(N__8783));
    Span4Mux_h I__736 (
            .O(N__8791),
            .I(N__8780));
    Odrv12 I__735 (
            .O(N__8788),
            .I(TVP_VIDEO_c_8));
    Odrv4 I__734 (
            .O(N__8783),
            .I(TVP_VIDEO_c_8));
    Odrv4 I__733 (
            .O(N__8780),
            .I(TVP_VIDEO_c_8));
    InMux I__732 (
            .O(N__8773),
            .I(N__8769));
    InMux I__731 (
            .O(N__8772),
            .I(N__8766));
    LocalMux I__730 (
            .O(N__8769),
            .I(N__8760));
    LocalMux I__729 (
            .O(N__8766),
            .I(N__8760));
    InMux I__728 (
            .O(N__8765),
            .I(N__8757));
    Span4Mux_v I__727 (
            .O(N__8760),
            .I(N__8752));
    LocalMux I__726 (
            .O(N__8757),
            .I(N__8752));
    Span4Mux_v I__725 (
            .O(N__8752),
            .I(N__8747));
    InMux I__724 (
            .O(N__8751),
            .I(N__8744));
    InMux I__723 (
            .O(N__8750),
            .I(N__8740));
    Span4Mux_v I__722 (
            .O(N__8747),
            .I(N__8735));
    LocalMux I__721 (
            .O(N__8744),
            .I(N__8735));
    InMux I__720 (
            .O(N__8743),
            .I(N__8732));
    LocalMux I__719 (
            .O(N__8740),
            .I(N__8729));
    Span4Mux_h I__718 (
            .O(N__8735),
            .I(N__8726));
    LocalMux I__717 (
            .O(N__8732),
            .I(N__8723));
    Span12Mux_s11_h I__716 (
            .O(N__8729),
            .I(N__8719));
    Sp12to4 I__715 (
            .O(N__8726),
            .I(N__8716));
    Span12Mux_s8_h I__714 (
            .O(N__8723),
            .I(N__8713));
    InMux I__713 (
            .O(N__8722),
            .I(N__8710));
    Span12Mux_h I__712 (
            .O(N__8719),
            .I(N__8707));
    Span12Mux_v I__711 (
            .O(N__8716),
            .I(N__8704));
    Span12Mux_v I__710 (
            .O(N__8713),
            .I(N__8701));
    LocalMux I__709 (
            .O(N__8710),
            .I(N__8698));
    Span12Mux_v I__708 (
            .O(N__8707),
            .I(N__8694));
    Span12Mux_h I__707 (
            .O(N__8704),
            .I(N__8691));
    Span12Mux_v I__706 (
            .O(N__8701),
            .I(N__8688));
    Span4Mux_h I__705 (
            .O(N__8698),
            .I(N__8685));
    InMux I__704 (
            .O(N__8697),
            .I(N__8682));
    Odrv12 I__703 (
            .O(N__8694),
            .I(TVP_VIDEO_c_9));
    Odrv12 I__702 (
            .O(N__8691),
            .I(TVP_VIDEO_c_9));
    Odrv12 I__701 (
            .O(N__8688),
            .I(TVP_VIDEO_c_9));
    Odrv4 I__700 (
            .O(N__8685),
            .I(TVP_VIDEO_c_9));
    LocalMux I__699 (
            .O(N__8682),
            .I(TVP_VIDEO_c_9));
    InMux I__698 (
            .O(N__8671),
            .I(N__8668));
    LocalMux I__697 (
            .O(N__8668),
            .I(N__8662));
    InMux I__696 (
            .O(N__8667),
            .I(N__8659));
    InMux I__695 (
            .O(N__8666),
            .I(N__8656));
    InMux I__694 (
            .O(N__8665),
            .I(N__8653));
    Span4Mux_h I__693 (
            .O(N__8662),
            .I(N__8650));
    LocalMux I__692 (
            .O(N__8659),
            .I(N__8646));
    LocalMux I__691 (
            .O(N__8656),
            .I(N__8643));
    LocalMux I__690 (
            .O(N__8653),
            .I(N__8639));
    Span4Mux_h I__689 (
            .O(N__8650),
            .I(N__8636));
    InMux I__688 (
            .O(N__8649),
            .I(N__8633));
    Span4Mux_h I__687 (
            .O(N__8646),
            .I(N__8630));
    Span4Mux_v I__686 (
            .O(N__8643),
            .I(N__8627));
    InMux I__685 (
            .O(N__8642),
            .I(N__8622));
    Span12Mux_h I__684 (
            .O(N__8639),
            .I(N__8619));
    Sp12to4 I__683 (
            .O(N__8636),
            .I(N__8616));
    LocalMux I__682 (
            .O(N__8633),
            .I(N__8613));
    Span4Mux_h I__681 (
            .O(N__8630),
            .I(N__8610));
    Span4Mux_v I__680 (
            .O(N__8627),
            .I(N__8607));
    InMux I__679 (
            .O(N__8626),
            .I(N__8604));
    InMux I__678 (
            .O(N__8625),
            .I(N__8601));
    LocalMux I__677 (
            .O(N__8622),
            .I(N__8598));
    Span12Mux_v I__676 (
            .O(N__8619),
            .I(N__8595));
    Span12Mux_v I__675 (
            .O(N__8616),
            .I(N__8588));
    Span12Mux_h I__674 (
            .O(N__8613),
            .I(N__8588));
    Sp12to4 I__673 (
            .O(N__8610),
            .I(N__8588));
    Sp12to4 I__672 (
            .O(N__8607),
            .I(N__8583));
    LocalMux I__671 (
            .O(N__8604),
            .I(N__8583));
    LocalMux I__670 (
            .O(N__8601),
            .I(N__8580));
    Span4Mux_h I__669 (
            .O(N__8598),
            .I(N__8577));
    Span12Mux_v I__668 (
            .O(N__8595),
            .I(N__8574));
    Span12Mux_v I__667 (
            .O(N__8588),
            .I(N__8567));
    Span12Mux_h I__666 (
            .O(N__8583),
            .I(N__8567));
    Span12Mux_h I__665 (
            .O(N__8580),
            .I(N__8567));
    Span4Mux_h I__664 (
            .O(N__8577),
            .I(N__8564));
    Odrv12 I__663 (
            .O(N__8574),
            .I(TVP_VIDEO_c_7));
    Odrv12 I__662 (
            .O(N__8567),
            .I(TVP_VIDEO_c_7));
    Odrv4 I__661 (
            .O(N__8564),
            .I(TVP_VIDEO_c_7));
    InMux I__660 (
            .O(N__8557),
            .I(N__8553));
    InMux I__659 (
            .O(N__8556),
            .I(N__8550));
    LocalMux I__658 (
            .O(N__8553),
            .I(N__8547));
    LocalMux I__657 (
            .O(N__8550),
            .I(N__8543));
    Span4Mux_v I__656 (
            .O(N__8547),
            .I(N__8540));
    InMux I__655 (
            .O(N__8546),
            .I(N__8537));
    Span4Mux_v I__654 (
            .O(N__8543),
            .I(N__8533));
    Span4Mux_v I__653 (
            .O(N__8540),
            .I(N__8528));
    LocalMux I__652 (
            .O(N__8537),
            .I(N__8528));
    InMux I__651 (
            .O(N__8536),
            .I(N__8525));
    Span4Mux_v I__650 (
            .O(N__8533),
            .I(N__8522));
    Span4Mux_v I__649 (
            .O(N__8528),
            .I(N__8516));
    LocalMux I__648 (
            .O(N__8525),
            .I(N__8516));
    Span4Mux_v I__647 (
            .O(N__8522),
            .I(N__8512));
    InMux I__646 (
            .O(N__8521),
            .I(N__8509));
    Span4Mux_v I__645 (
            .O(N__8516),
            .I(N__8505));
    InMux I__644 (
            .O(N__8515),
            .I(N__8502));
    Span4Mux_v I__643 (
            .O(N__8512),
            .I(N__8497));
    LocalMux I__642 (
            .O(N__8509),
            .I(N__8497));
    InMux I__641 (
            .O(N__8508),
            .I(N__8494));
    Span4Mux_v I__640 (
            .O(N__8505),
            .I(N__8489));
    LocalMux I__639 (
            .O(N__8502),
            .I(N__8489));
    Span4Mux_v I__638 (
            .O(N__8497),
            .I(N__8484));
    LocalMux I__637 (
            .O(N__8494),
            .I(N__8484));
    Span4Mux_v I__636 (
            .O(N__8489),
            .I(N__8480));
    Span4Mux_v I__635 (
            .O(N__8484),
            .I(N__8477));
    InMux I__634 (
            .O(N__8483),
            .I(N__8474));
    Sp12to4 I__633 (
            .O(N__8480),
            .I(N__8471));
    Span4Mux_v I__632 (
            .O(N__8477),
            .I(N__8466));
    LocalMux I__631 (
            .O(N__8474),
            .I(N__8466));
    Span12Mux_h I__630 (
            .O(N__8471),
            .I(N__8463));
    Span4Mux_h I__629 (
            .O(N__8466),
            .I(N__8460));
    Odrv12 I__628 (
            .O(N__8463),
            .I(TVP_VIDEO_c_6));
    Odrv4 I__627 (
            .O(N__8460),
            .I(TVP_VIDEO_c_6));
    InMux I__626 (
            .O(N__8455),
            .I(N__8452));
    LocalMux I__625 (
            .O(N__8452),
            .I(N__8448));
    InMux I__624 (
            .O(N__8451),
            .I(N__8444));
    Span4Mux_v I__623 (
            .O(N__8448),
            .I(N__8441));
    InMux I__622 (
            .O(N__8447),
            .I(N__8437));
    LocalMux I__621 (
            .O(N__8444),
            .I(N__8434));
    Span4Mux_v I__620 (
            .O(N__8441),
            .I(N__8430));
    InMux I__619 (
            .O(N__8440),
            .I(N__8427));
    LocalMux I__618 (
            .O(N__8437),
            .I(N__8424));
    Span4Mux_v I__617 (
            .O(N__8434),
            .I(N__8421));
    InMux I__616 (
            .O(N__8433),
            .I(N__8418));
    Span4Mux_v I__615 (
            .O(N__8430),
            .I(N__8412));
    LocalMux I__614 (
            .O(N__8427),
            .I(N__8412));
    Span4Mux_h I__613 (
            .O(N__8424),
            .I(N__8408));
    Span4Mux_v I__612 (
            .O(N__8421),
            .I(N__8403));
    LocalMux I__611 (
            .O(N__8418),
            .I(N__8403));
    InMux I__610 (
            .O(N__8417),
            .I(N__8400));
    Span4Mux_v I__609 (
            .O(N__8412),
            .I(N__8397));
    InMux I__608 (
            .O(N__8411),
            .I(N__8394));
    Sp12to4 I__607 (
            .O(N__8408),
            .I(N__8391));
    Span4Mux_v I__606 (
            .O(N__8403),
            .I(N__8386));
    LocalMux I__605 (
            .O(N__8400),
            .I(N__8386));
    Span4Mux_v I__604 (
            .O(N__8397),
            .I(N__8381));
    LocalMux I__603 (
            .O(N__8394),
            .I(N__8381));
    Span12Mux_v I__602 (
            .O(N__8391),
            .I(N__8377));
    Span4Mux_v I__601 (
            .O(N__8386),
            .I(N__8374));
    Span4Mux_v I__600 (
            .O(N__8381),
            .I(N__8371));
    InMux I__599 (
            .O(N__8380),
            .I(N__8368));
    Span12Mux_v I__598 (
            .O(N__8377),
            .I(N__8363));
    Sp12to4 I__597 (
            .O(N__8374),
            .I(N__8363));
    Span4Mux_v I__596 (
            .O(N__8371),
            .I(N__8358));
    LocalMux I__595 (
            .O(N__8368),
            .I(N__8358));
    Span12Mux_h I__594 (
            .O(N__8363),
            .I(N__8355));
    Span4Mux_h I__593 (
            .O(N__8358),
            .I(N__8352));
    Odrv12 I__592 (
            .O(N__8355),
            .I(TVP_VIDEO_c_5));
    Odrv4 I__591 (
            .O(N__8352),
            .I(TVP_VIDEO_c_5));
    InMux I__590 (
            .O(N__8347),
            .I(N__8343));
    InMux I__589 (
            .O(N__8346),
            .I(N__8340));
    LocalMux I__588 (
            .O(N__8343),
            .I(N__8337));
    LocalMux I__587 (
            .O(N__8340),
            .I(N__8332));
    Span4Mux_v I__586 (
            .O(N__8337),
            .I(N__8329));
    InMux I__585 (
            .O(N__8336),
            .I(N__8326));
    InMux I__584 (
            .O(N__8335),
            .I(N__8322));
    Span4Mux_s1_v I__583 (
            .O(N__8332),
            .I(N__8318));
    Span4Mux_v I__582 (
            .O(N__8329),
            .I(N__8313));
    LocalMux I__581 (
            .O(N__8326),
            .I(N__8313));
    InMux I__580 (
            .O(N__8325),
            .I(N__8310));
    LocalMux I__579 (
            .O(N__8322),
            .I(N__8307));
    InMux I__578 (
            .O(N__8321),
            .I(N__8304));
    Span4Mux_h I__577 (
            .O(N__8318),
            .I(N__8301));
    Span4Mux_v I__576 (
            .O(N__8313),
            .I(N__8296));
    LocalMux I__575 (
            .O(N__8310),
            .I(N__8296));
    Span4Mux_h I__574 (
            .O(N__8307),
            .I(N__8293));
    LocalMux I__573 (
            .O(N__8304),
            .I(N__8290));
    Span4Mux_v I__572 (
            .O(N__8301),
            .I(N__8286));
    Span4Mux_v I__571 (
            .O(N__8296),
            .I(N__8283));
    Span4Mux_h I__570 (
            .O(N__8293),
            .I(N__8280));
    Span4Mux_h I__569 (
            .O(N__8290),
            .I(N__8277));
    InMux I__568 (
            .O(N__8289),
            .I(N__8274));
    Sp12to4 I__567 (
            .O(N__8286),
            .I(N__8271));
    Span4Mux_h I__566 (
            .O(N__8283),
            .I(N__8268));
    Span4Mux_h I__565 (
            .O(N__8280),
            .I(N__8265));
    Span4Mux_v I__564 (
            .O(N__8277),
            .I(N__8262));
    LocalMux I__563 (
            .O(N__8274),
            .I(N__8259));
    Span12Mux_h I__562 (
            .O(N__8271),
            .I(N__8255));
    Sp12to4 I__561 (
            .O(N__8268),
            .I(N__8252));
    Span4Mux_h I__560 (
            .O(N__8265),
            .I(N__8245));
    Span4Mux_v I__559 (
            .O(N__8262),
            .I(N__8245));
    Span4Mux_h I__558 (
            .O(N__8259),
            .I(N__8245));
    InMux I__557 (
            .O(N__8258),
            .I(N__8242));
    Span12Mux_v I__556 (
            .O(N__8255),
            .I(N__8237));
    Span12Mux_h I__555 (
            .O(N__8252),
            .I(N__8237));
    Span4Mux_v I__554 (
            .O(N__8245),
            .I(N__8234));
    LocalMux I__553 (
            .O(N__8242),
            .I(N__8231));
    Span12Mux_v I__552 (
            .O(N__8237),
            .I(N__8228));
    Span4Mux_v I__551 (
            .O(N__8234),
            .I(N__8225));
    Span4Mux_h I__550 (
            .O(N__8231),
            .I(N__8222));
    Odrv12 I__549 (
            .O(N__8228),
            .I(TVP_VIDEO_c_4));
    Odrv4 I__548 (
            .O(N__8225),
            .I(TVP_VIDEO_c_4));
    Odrv4 I__547 (
            .O(N__8222),
            .I(TVP_VIDEO_c_4));
    InMux I__546 (
            .O(N__8215),
            .I(N__8211));
    InMux I__545 (
            .O(N__8214),
            .I(N__8208));
    LocalMux I__544 (
            .O(N__8211),
            .I(N__8203));
    LocalMux I__543 (
            .O(N__8208),
            .I(N__8200));
    InMux I__542 (
            .O(N__8207),
            .I(N__8197));
    InMux I__541 (
            .O(N__8206),
            .I(N__8194));
    Sp12to4 I__540 (
            .O(N__8203),
            .I(N__8190));
    Span4Mux_h I__539 (
            .O(N__8200),
            .I(N__8187));
    LocalMux I__538 (
            .O(N__8197),
            .I(N__8184));
    LocalMux I__537 (
            .O(N__8194),
            .I(N__8179));
    InMux I__536 (
            .O(N__8193),
            .I(N__8176));
    Span12Mux_h I__535 (
            .O(N__8190),
            .I(N__8172));
    Span4Mux_h I__534 (
            .O(N__8187),
            .I(N__8169));
    Span4Mux_v I__533 (
            .O(N__8184),
            .I(N__8166));
    InMux I__532 (
            .O(N__8183),
            .I(N__8163));
    InMux I__531 (
            .O(N__8182),
            .I(N__8160));
    Span12Mux_h I__530 (
            .O(N__8179),
            .I(N__8157));
    LocalMux I__529 (
            .O(N__8176),
            .I(N__8154));
    InMux I__528 (
            .O(N__8175),
            .I(N__8151));
    Span12Mux_v I__527 (
            .O(N__8172),
            .I(N__8146));
    Sp12to4 I__526 (
            .O(N__8169),
            .I(N__8146));
    Sp12to4 I__525 (
            .O(N__8166),
            .I(N__8143));
    LocalMux I__524 (
            .O(N__8163),
            .I(N__8140));
    LocalMux I__523 (
            .O(N__8160),
            .I(N__8137));
    Span12Mux_v I__522 (
            .O(N__8157),
            .I(N__8130));
    Span12Mux_h I__521 (
            .O(N__8154),
            .I(N__8130));
    LocalMux I__520 (
            .O(N__8151),
            .I(N__8130));
    Span12Mux_v I__519 (
            .O(N__8146),
            .I(N__8125));
    Span12Mux_h I__518 (
            .O(N__8143),
            .I(N__8125));
    Span12Mux_h I__517 (
            .O(N__8140),
            .I(N__8122));
    Span4Mux_h I__516 (
            .O(N__8137),
            .I(N__8119));
    Span12Mux_h I__515 (
            .O(N__8130),
            .I(N__8116));
    Span12Mux_h I__514 (
            .O(N__8125),
            .I(N__8109));
    Span12Mux_v I__513 (
            .O(N__8122),
            .I(N__8109));
    Sp12to4 I__512 (
            .O(N__8119),
            .I(N__8109));
    Odrv12 I__511 (
            .O(N__8116),
            .I(TVP_VIDEO_c_3));
    Odrv12 I__510 (
            .O(N__8109),
            .I(TVP_VIDEO_c_3));
    INV INVADV_R__i2C (
            .O(INVADV_R__i2C_net),
            .I(N__22547));
    INV \INVdb5.NEXT_COUNTER__i3C  (
            .O(\INVdb5.NEXT_COUNTER__i3C_net ),
            .I(N__19340));
    INV INVADV_R__i1C (
            .O(INVADV_R__i1C_net),
            .I(N__22535));
    defparam IN_MUX_bfv_12_16_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_16_0_));
    defparam IN_MUX_bfv_12_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_17_0_ (
            .carryinitin(\transmit_module.video_signal_controller.n3684 ),
            .carryinitout(bfn_12_17_0_));
    defparam IN_MUX_bfv_13_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_15_0_));
    defparam IN_MUX_bfv_13_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_16_0_ (
            .carryinitin(\transmit_module.video_signal_controller.n3695 ),
            .carryinitout(bfn_13_16_0_));
    defparam IN_MUX_bfv_15_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_17_0_));
    defparam IN_MUX_bfv_15_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_18_0_ (
            .carryinitin(\transmit_module.n3663 ),
            .carryinitout(bfn_15_18_0_));
    defparam IN_MUX_bfv_13_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_10_0_));
    defparam IN_MUX_bfv_11_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_9_0_));
    defparam IN_MUX_bfv_11_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_10_0_ (
            .carryinitin(\receive_module.rx_counter.n3718 ),
            .carryinitout(bfn_11_10_0_));
    defparam IN_MUX_bfv_10_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_9_0_));
    defparam IN_MUX_bfv_10_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_10_0_ (
            .carryinitin(\receive_module.rx_counter.n3676 ),
            .carryinitout(bfn_10_10_0_));
    defparam IN_MUX_bfv_14_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_9_0_));
    defparam IN_MUX_bfv_14_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_10_0_ (
            .carryinitin(\receive_module.rx_counter.n3727 ),
            .carryinitout(bfn_14_10_0_));
    defparam IN_MUX_bfv_15_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_8_0_));
    defparam IN_MUX_bfv_13_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_11_0_));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \receive_module.rx_counter.i4_2_lut_LC_9_9_2 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i4_2_lut_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i4_2_lut_LC_9_9_2 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \receive_module.rx_counter.i4_2_lut_LC_9_9_2  (
            .in0(_gnd_net_),
            .in1(N__9444),
            .in2(_gnd_net_),
            .in3(N__9565),
            .lcout(),
            .ltout(\receive_module.rx_counter.n12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.SYNC_45_LC_9_9_3 .C_ON=1'b0;
    defparam \receive_module.rx_counter.SYNC_45_LC_9_9_3 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.SYNC_45_LC_9_9_3 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \receive_module.rx_counter.SYNC_45_LC_9_9_3  (
            .in0(N__8890),
            .in1(N__9594),
            .in2(N__8902),
            .in3(N__9310),
            .lcout(DEBUG_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19342),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i1_2_lut_LC_9_10_0 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i1_2_lut_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i1_2_lut_LC_9_10_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \receive_module.rx_counter.i1_2_lut_LC_9_10_0  (
            .in0(_gnd_net_),
            .in1(N__9488),
            .in2(_gnd_net_),
            .in3(N__9513),
            .lcout(\receive_module.rx_counter.n3938 ),
            .ltout(\receive_module.rx_counter.n3938_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i2_4_lut_LC_9_10_1 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i2_4_lut_LC_9_10_1 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i2_4_lut_LC_9_10_1 .LUT_INIT=16'b1000100010000000;
    LogicCell40 \receive_module.rx_counter.i2_4_lut_LC_9_10_1  (
            .in0(N__9467),
            .in1(N__9442),
            .in2(N__8899),
            .in3(N__9202),
            .lcout(\receive_module.rx_counter.n3979 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i5_4_lut_LC_9_10_2 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i5_4_lut_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i5_4_lut_LC_9_10_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \receive_module.rx_counter.i5_4_lut_LC_9_10_2  (
            .in0(N__8896),
            .in1(N__9537),
            .in2(N__9625),
            .in3(N__9468),
            .lcout(\receive_module.rx_counter.n13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i1803_2_lut_LC_9_10_6 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i1803_2_lut_LC_9_10_6 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i1803_2_lut_LC_9_10_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \receive_module.rx_counter.i1803_2_lut_LC_9_10_6  (
            .in0(_gnd_net_),
            .in1(N__9620),
            .in2(_gnd_net_),
            .in3(N__9308),
            .lcout(),
            .ltout(\receive_module.rx_counter.n3176_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i1835_4_lut_LC_9_10_7 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i1835_4_lut_LC_9_10_7 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i1835_4_lut_LC_9_10_7 .LUT_INIT=16'b1010101010101000;
    LogicCell40 \receive_module.rx_counter.i1835_4_lut_LC_9_10_7  (
            .in0(N__9536),
            .in1(N__9563),
            .in2(N__9205),
            .in3(N__9592),
            .lcout(\receive_module.rx_counter.n3208 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2693_LC_9_15_3 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2693_LC_9_15_3 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2693_LC_9_15_3 .LUT_INIT=16'b1111100000111000;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_2693_LC_9_15_3  (
            .in0(N__9196),
            .in1(N__23838),
            .in2(N__23613),
            .in3(N__9175),
            .lcout(),
            .ltout(\line_buffer.n4170_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n4170_bdd_4_lut_LC_9_15_4 .C_ON=1'b0;
    defparam \line_buffer.n4170_bdd_4_lut_LC_9_15_4 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n4170_bdd_4_lut_LC_9_15_4 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \line_buffer.n4170_bdd_4_lut_LC_9_15_4  (
            .in0(N__23839),
            .in1(N__9166),
            .in2(N__9145),
            .in3(N__9142),
            .lcout(\line_buffer.n4173 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2678_LC_9_15_5 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2678_LC_9_15_5 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2678_LC_9_15_5 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_2678_LC_9_15_5  (
            .in0(N__9127),
            .in1(N__23837),
            .in2(N__9109),
            .in3(N__23604),
            .lcout(\line_buffer.n4152 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2598_3_lut_LC_9_15_6 .C_ON=1'b0;
    defparam \line_buffer.i2598_3_lut_LC_9_15_6 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2598_3_lut_LC_9_15_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \line_buffer.i2598_3_lut_LC_9_15_6  (
            .in0(N__23603),
            .in1(N__9094),
            .in2(_gnd_net_),
            .in3(N__9079),
            .lcout(\line_buffer.n4072 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n4152_bdd_4_lut_LC_9_16_2 .C_ON=1'b0;
    defparam \line_buffer.n4152_bdd_4_lut_LC_9_16_2 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n4152_bdd_4_lut_LC_9_16_2 .LUT_INIT=16'b1010101011011000;
    LogicCell40 \line_buffer.n4152_bdd_4_lut_LC_9_16_2  (
            .in0(N__9073),
            .in1(N__9067),
            .in2(N__9046),
            .in3(N__23863),
            .lcout(),
            .ltout(\line_buffer.n4155_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i2_LC_9_16_3 .C_ON=1'b0;
    defparam \line_buffer.dout_i2_LC_9_16_3 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i2_LC_9_16_3 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \line_buffer.dout_i2_LC_9_16_3  (
            .in0(_gnd_net_),
            .in1(N__22846),
            .in2(N__9025),
            .in3(N__9022),
            .lcout(TX_DATA_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22650),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.Y_DELTA_PATTERN_i90_LC_9_17_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i90_LC_9_17_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i90_LC_9_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i90_LC_9_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9397),
            .lcout(\transmit_module.Y_DELTA_PATTERN_90 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22581),
            .ce(N__16039),
            .sr(N__21279));
    defparam \transmit_module.Y_DELTA_PATTERN_i94_LC_9_18_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i94_LC_9_18_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i94_LC_9_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i94_LC_9_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9256),
            .lcout(\transmit_module.Y_DELTA_PATTERN_94 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22563),
            .ce(N__16037),
            .sr(N__21151));
    defparam \transmit_module.Y_DELTA_PATTERN_i95_LC_9_18_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i95_LC_9_18_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i95_LC_9_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i95_LC_9_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9364),
            .lcout(\transmit_module.Y_DELTA_PATTERN_95 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22563),
            .ce(N__16037),
            .sr(N__21151));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2668_LC_9_21_0 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2668_LC_9_21_0 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2668_LC_9_21_0 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_2668_LC_9_21_0  (
            .in0(N__9250),
            .in1(N__23844),
            .in2(N__9238),
            .in3(N__23543),
            .lcout(\line_buffer.n4122 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.Y__i0_LC_10_9_0 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i0_LC_10_9_0 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i0_LC_10_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i0_LC_10_9_0  (
            .in0(_gnd_net_),
            .in1(N__9309),
            .in2(_gnd_net_),
            .in3(N__9223),
            .lcout(\receive_module.rx_counter.Y_0 ),
            .ltout(),
            .carryin(bfn_10_9_0_),
            .carryout(\receive_module.rx_counter.n3669 ),
            .clk(N__19334),
            .ce(N__11691),
            .sr(N__9768));
    defparam \receive_module.rx_counter.Y__i1_LC_10_9_1 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i1_LC_10_9_1 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i1_LC_10_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i1_LC_10_9_1  (
            .in0(_gnd_net_),
            .in1(N__9621),
            .in2(_gnd_net_),
            .in3(N__9220),
            .lcout(\receive_module.rx_counter.Y_1 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3669 ),
            .carryout(\receive_module.rx_counter.n3670 ),
            .clk(N__19334),
            .ce(N__11691),
            .sr(N__9768));
    defparam \receive_module.rx_counter.Y__i2_LC_10_9_2 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i2_LC_10_9_2 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i2_LC_10_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i2_LC_10_9_2  (
            .in0(_gnd_net_),
            .in1(N__9593),
            .in2(_gnd_net_),
            .in3(N__9217),
            .lcout(\receive_module.rx_counter.Y_2 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3670 ),
            .carryout(\receive_module.rx_counter.n3671 ),
            .clk(N__19334),
            .ce(N__11691),
            .sr(N__9768));
    defparam \receive_module.rx_counter.Y__i3_LC_10_9_3 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i3_LC_10_9_3 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i3_LC_10_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i3_LC_10_9_3  (
            .in0(_gnd_net_),
            .in1(N__9564),
            .in2(_gnd_net_),
            .in3(N__9214),
            .lcout(\receive_module.rx_counter.Y_3 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3671 ),
            .carryout(\receive_module.rx_counter.n3672 ),
            .clk(N__19334),
            .ce(N__11691),
            .sr(N__9768));
    defparam \receive_module.rx_counter.Y__i4_LC_10_9_4 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i4_LC_10_9_4 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i4_LC_10_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i4_LC_10_9_4  (
            .in0(_gnd_net_),
            .in1(N__9538),
            .in2(_gnd_net_),
            .in3(N__9211),
            .lcout(\receive_module.rx_counter.Y_4 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3672 ),
            .carryout(\receive_module.rx_counter.n3673 ),
            .clk(N__19334),
            .ce(N__11691),
            .sr(N__9768));
    defparam \receive_module.rx_counter.Y__i5_LC_10_9_5 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i5_LC_10_9_5 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i5_LC_10_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i5_LC_10_9_5  (
            .in0(_gnd_net_),
            .in1(N__9514),
            .in2(_gnd_net_),
            .in3(N__9208),
            .lcout(\receive_module.rx_counter.Y_5 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3673 ),
            .carryout(\receive_module.rx_counter.n3674 ),
            .clk(N__19334),
            .ce(N__11691),
            .sr(N__9768));
    defparam \receive_module.rx_counter.Y__i6_LC_10_9_6 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i6_LC_10_9_6 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i6_LC_10_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i6_LC_10_9_6  (
            .in0(_gnd_net_),
            .in1(N__9492),
            .in2(_gnd_net_),
            .in3(N__9283),
            .lcout(\receive_module.rx_counter.Y_6 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3674 ),
            .carryout(\receive_module.rx_counter.n3675 ),
            .clk(N__19334),
            .ce(N__11691),
            .sr(N__9768));
    defparam \receive_module.rx_counter.Y__i7_LC_10_9_7 .C_ON=1'b1;
    defparam \receive_module.rx_counter.Y__i7_LC_10_9_7 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i7_LC_10_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i7_LC_10_9_7  (
            .in0(_gnd_net_),
            .in1(N__9469),
            .in2(_gnd_net_),
            .in3(N__9280),
            .lcout(\receive_module.rx_counter.Y_7 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3675 ),
            .carryout(\receive_module.rx_counter.n3676 ),
            .clk(N__19334),
            .ce(N__11691),
            .sr(N__9768));
    defparam \receive_module.rx_counter.Y__i8_LC_10_10_0 .C_ON=1'b0;
    defparam \receive_module.rx_counter.Y__i8_LC_10_10_0 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.Y__i8_LC_10_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.Y__i8_LC_10_10_0  (
            .in0(_gnd_net_),
            .in1(N__9445),
            .in2(_gnd_net_),
            .in3(N__9277),
            .lcout(\receive_module.rx_counter.Y_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19338),
            .ce(N__11692),
            .sr(N__9772));
    defparam \transmit_module.Y_DELTA_PATTERN_i84_LC_10_15_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i84_LC_10_15_2 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i84_LC_10_15_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i84_LC_10_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9385),
            .lcout(\transmit_module.Y_DELTA_PATTERN_84 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22537),
            .ce(N__16036),
            .sr(N__21056));
    defparam \transmit_module.Y_DELTA_PATTERN_i83_LC_10_15_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i83_LC_10_15_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i83_LC_10_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i83_LC_10_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9274),
            .lcout(\transmit_module.Y_DELTA_PATTERN_83 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22537),
            .ce(N__16036),
            .sr(N__21056));
    defparam \transmit_module.Y_DELTA_PATTERN_i82_LC_10_16_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i82_LC_10_16_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i82_LC_10_16_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i82_LC_10_16_1  (
            .in0(N__9268),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.Y_DELTA_PATTERN_82 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22649),
            .ce(N__21457),
            .sr(N__20955));
    defparam \transmit_module.Y_DELTA_PATTERN_i87_LC_10_17_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i87_LC_10_17_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i87_LC_10_17_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i87_LC_10_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9415),
            .lcout(\transmit_module.Y_DELTA_PATTERN_87 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22578),
            .ce(N__16029),
            .sr(N__21321));
    defparam \transmit_module.Y_DELTA_PATTERN_i92_LC_10_17_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i92_LC_10_17_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i92_LC_10_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i92_LC_10_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9370),
            .lcout(\transmit_module.Y_DELTA_PATTERN_92 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22578),
            .ce(N__16029),
            .sr(N__21321));
    defparam \transmit_module.Y_DELTA_PATTERN_i89_LC_10_17_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i89_LC_10_17_2 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i89_LC_10_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i89_LC_10_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9262),
            .lcout(\transmit_module.Y_DELTA_PATTERN_89 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22578),
            .ce(N__16029),
            .sr(N__21321));
    defparam \transmit_module.Y_DELTA_PATTERN_i88_LC_10_17_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i88_LC_10_17_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i88_LC_10_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i88_LC_10_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9421),
            .lcout(\transmit_module.Y_DELTA_PATTERN_88 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22578),
            .ce(N__16029),
            .sr(N__21321));
    defparam \transmit_module.Y_DELTA_PATTERN_i86_LC_10_17_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i86_LC_10_17_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i86_LC_10_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i86_LC_10_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9409),
            .lcout(\transmit_module.Y_DELTA_PATTERN_86 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22578),
            .ce(N__16029),
            .sr(N__21321));
    defparam \transmit_module.Y_DELTA_PATTERN_i91_LC_10_17_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i91_LC_10_17_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i91_LC_10_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i91_LC_10_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9403),
            .lcout(\transmit_module.Y_DELTA_PATTERN_91 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22578),
            .ce(N__16029),
            .sr(N__21321));
    defparam \transmit_module.Y_DELTA_PATTERN_i85_LC_10_17_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i85_LC_10_17_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i85_LC_10_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i85_LC_10_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9391),
            .lcout(\transmit_module.Y_DELTA_PATTERN_85 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22578),
            .ce(N__16029),
            .sr(N__21321));
    defparam \transmit_module.Y_DELTA_PATTERN_i93_LC_10_18_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i93_LC_10_18_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i93_LC_10_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i93_LC_10_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9376),
            .lcout(\transmit_module.Y_DELTA_PATTERN_93 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22564),
            .ce(N__20596),
            .sr(N__21251));
    defparam \transmit_module.Y_DELTA_PATTERN_i96_LC_10_19_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i96_LC_10_19_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i96_LC_10_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i96_LC_10_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9358),
            .lcout(\transmit_module.Y_DELTA_PATTERN_96 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22435),
            .ce(N__21480),
            .sr(N__21055));
    defparam \transmit_module.Y_DELTA_PATTERN_i97_LC_10_19_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i97_LC_10_19_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i97_LC_10_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i97_LC_10_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9739),
            .lcout(\transmit_module.Y_DELTA_PATTERN_97 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22435),
            .ce(N__21480),
            .sr(N__21055));
    defparam \line_buffer.n4122_bdd_4_lut_LC_10_21_2 .C_ON=1'b0;
    defparam \line_buffer.n4122_bdd_4_lut_LC_10_21_2 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n4122_bdd_4_lut_LC_10_21_2 .LUT_INIT=16'b1100110010111000;
    LogicCell40 \line_buffer.n4122_bdd_4_lut_LC_10_21_2  (
            .in0(N__9352),
            .in1(N__9343),
            .in2(N__9337),
            .in3(N__23845),
            .lcout(\line_buffer.n4125 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.sub_23_add_2_2_lut_LC_11_9_0 .C_ON=1'b1;
    defparam \receive_module.rx_counter.sub_23_add_2_2_lut_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.sub_23_add_2_2_lut_LC_11_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.sub_23_add_2_2_lut_LC_11_9_0  (
            .in0(_gnd_net_),
            .in1(N__9307),
            .in2(_gnd_net_),
            .in3(N__9286),
            .lcout(\receive_module.O_Y_0 ),
            .ltout(),
            .carryin(bfn_11_9_0_),
            .carryout(\receive_module.rx_counter.n3711 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.sub_23_add_2_3_lut_LC_11_9_1 .C_ON=1'b1;
    defparam \receive_module.rx_counter.sub_23_add_2_3_lut_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.sub_23_add_2_3_lut_LC_11_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.sub_23_add_2_3_lut_LC_11_9_1  (
            .in0(_gnd_net_),
            .in1(N__9619),
            .in2(N__23307),
            .in3(N__9598),
            .lcout(\receive_module.O_Y_1 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3711 ),
            .carryout(\receive_module.rx_counter.n3712 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.sub_23_add_2_4_lut_LC_11_9_2 .C_ON=1'b1;
    defparam \receive_module.rx_counter.sub_23_add_2_4_lut_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.sub_23_add_2_4_lut_LC_11_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.sub_23_add_2_4_lut_LC_11_9_2  (
            .in0(_gnd_net_),
            .in1(N__23252),
            .in2(N__9595),
            .in3(N__9568),
            .lcout(\receive_module.O_Y_2 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3712 ),
            .carryout(\receive_module.rx_counter.n3713 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.sub_23_add_2_5_lut_LC_11_9_3 .C_ON=1'b1;
    defparam \receive_module.rx_counter.sub_23_add_2_5_lut_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.sub_23_add_2_5_lut_LC_11_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.sub_23_add_2_5_lut_LC_11_9_3  (
            .in0(_gnd_net_),
            .in1(N__9562),
            .in2(_gnd_net_),
            .in3(N__9541),
            .lcout(\receive_module.O_Y_3 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3713 ),
            .carryout(\receive_module.rx_counter.n3714 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.sub_23_add_2_6_lut_LC_11_9_4 .C_ON=1'b1;
    defparam \receive_module.rx_counter.sub_23_add_2_6_lut_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.sub_23_add_2_6_lut_LC_11_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.sub_23_add_2_6_lut_LC_11_9_4  (
            .in0(_gnd_net_),
            .in1(N__9535),
            .in2(_gnd_net_),
            .in3(N__9517),
            .lcout(\receive_module.O_Y_4 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3714 ),
            .carryout(\receive_module.rx_counter.n3715 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.sub_23_add_2_7_lut_LC_11_9_5 .C_ON=1'b1;
    defparam \receive_module.rx_counter.sub_23_add_2_7_lut_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.sub_23_add_2_7_lut_LC_11_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.sub_23_add_2_7_lut_LC_11_9_5  (
            .in0(_gnd_net_),
            .in1(N__9512),
            .in2(N__23308),
            .in3(N__9496),
            .lcout(\receive_module.O_Y_5 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3715 ),
            .carryout(\receive_module.rx_counter.n3716 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.sub_23_add_2_8_lut_LC_11_9_6 .C_ON=1'b1;
    defparam \receive_module.rx_counter.sub_23_add_2_8_lut_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.sub_23_add_2_8_lut_LC_11_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.sub_23_add_2_8_lut_LC_11_9_6  (
            .in0(_gnd_net_),
            .in1(N__23256),
            .in2(N__9493),
            .in3(N__9472),
            .lcout(\receive_module.O_Y_6 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3716 ),
            .carryout(\receive_module.rx_counter.n3717 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.sub_23_add_2_9_lut_LC_11_9_7 .C_ON=1'b1;
    defparam \receive_module.rx_counter.sub_23_add_2_9_lut_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.sub_23_add_2_9_lut_LC_11_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.sub_23_add_2_9_lut_LC_11_9_7  (
            .in0(_gnd_net_),
            .in1(N__9466),
            .in2(N__23309),
            .in3(N__9448),
            .lcout(\receive_module.O_Y_7 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3717 ),
            .carryout(\receive_module.rx_counter.n3718 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.sub_23_add_2_10_LC_11_10_0 .C_ON=1'b1;
    defparam \receive_module.rx_counter.sub_23_add_2_10_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.sub_23_add_2_10_LC_11_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \receive_module.rx_counter.sub_23_add_2_10_LC_11_10_0  (
            .in0(_gnd_net_),
            .in1(N__9443),
            .in2(N__23306),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_10_0_),
            .carryout(\receive_module.rx_counter.O_VISIBLE_N_89 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i3_4_lut_LC_11_10_1 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i3_4_lut_LC_11_10_1 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i3_4_lut_LC_11_10_1 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \receive_module.rx_counter.i3_4_lut_LC_11_10_1  (
            .in0(N__10126),
            .in1(N__17386),
            .in2(N__9691),
            .in3(N__9679),
            .lcout(DEBUG_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.SYNC_BUFF1_57_LC_11_15_4 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.SYNC_BUFF1_57_LC_11_15_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.SYNC_BUFF1_57_LC_11_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.video_signal_controller.SYNC_BUFF1_57_LC_11_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9672),
            .lcout(\transmit_module.video_signal_controller.SYNC_BUFF1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22580),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.SYNC_BUFF2_58_LC_11_15_5 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.SYNC_BUFF2_58_LC_11_15_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.SYNC_BUFF2_58_LC_11_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.video_signal_controller.SYNC_BUFF2_58_LC_11_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9643),
            .lcout(\transmit_module.video_signal_controller.SYNC_BUFF2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22580),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i3_4_lut_LC_11_16_5 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i3_4_lut_LC_11_16_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i3_4_lut_LC_11_16_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \transmit_module.video_signal_controller.i3_4_lut_LC_11_16_5  (
            .in0(N__10560),
            .in1(N__10402),
            .in2(N__10527),
            .in3(N__10495),
            .lcout(),
            .ltout(\transmit_module.video_signal_controller.n3987_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.VGA_VS_61_LC_11_16_6 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.VGA_VS_61_LC_11_16_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_VS_61_LC_11_16_6 .LUT_INIT=16'b0000111100001100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_VS_61_LC_11_16_6  (
            .in0(_gnd_net_),
            .in1(N__10444),
            .in2(N__9637),
            .in3(N__10428),
            .lcout(ADV_VSYNC_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22438),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_3_lut_4_lut_adj_17_LC_11_17_0 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_3_lut_4_lut_adj_17_LC_11_17_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_3_lut_4_lut_adj_17_LC_11_17_0 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \transmit_module.video_signal_controller.i1_3_lut_4_lut_adj_17_LC_11_17_0  (
            .in0(N__10400),
            .in1(N__10516),
            .in2(N__10429),
            .in3(N__10555),
            .lcout(),
            .ltout(\transmit_module.video_signal_controller.n4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_4_lut_LC_11_17_1 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_4_lut_LC_11_17_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_4_lut_LC_11_17_1 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \transmit_module.video_signal_controller.i1_4_lut_LC_11_17_1  (
            .in0(N__10350),
            .in1(N__9631),
            .in2(N__9634),
            .in3(N__10371),
            .lcout(\transmit_module.video_signal_controller.n3936 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_2_lut_3_lut_LC_11_17_2 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_2_lut_3_lut_LC_11_17_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_2_lut_3_lut_LC_11_17_2 .LUT_INIT=16'b1111111011111110;
    LogicCell40 \transmit_module.video_signal_controller.i1_2_lut_3_lut_LC_11_17_2  (
            .in0(N__10901),
            .in1(N__10349),
            .in2(N__10924),
            .in3(_gnd_net_),
            .lcout(\transmit_module.video_signal_controller.n6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_24_LC_11_17_3 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_24_LC_11_17_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_24_LC_11_17_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \transmit_module.video_signal_controller.i1_2_lut_rep_24_LC_11_17_3  (
            .in0(_gnd_net_),
            .in1(N__10423),
            .in2(_gnd_net_),
            .in3(N__10399),
            .lcout(\transmit_module.video_signal_controller.n4215 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_2_lut_adj_12_LC_11_17_5 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_2_lut_adj_12_LC_11_17_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_2_lut_adj_12_LC_11_17_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \transmit_module.video_signal_controller.i1_2_lut_adj_12_LC_11_17_5  (
            .in0(_gnd_net_),
            .in1(N__10623),
            .in2(_gnd_net_),
            .in3(N__10608),
            .lcout(\transmit_module.video_signal_controller.n3935 ),
            .ltout(\transmit_module.video_signal_controller.n3935_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i4_4_lut_LC_11_17_6 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i4_4_lut_LC_11_17_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i4_4_lut_LC_11_17_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \transmit_module.video_signal_controller.i4_4_lut_LC_11_17_6  (
            .in0(N__10481),
            .in1(N__10370),
            .in2(N__9748),
            .in3(N__9745),
            .lcout(\transmit_module.video_signal_controller.n3892 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.Y_DELTA_PATTERN_i98_LC_11_18_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i98_LC_11_18_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i98_LC_11_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i98_LC_11_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19603),
            .lcout(\transmit_module.Y_DELTA_PATTERN_98 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22437),
            .ce(N__16038),
            .sr(N__21252));
    defparam \transmit_module.Y_DELTA_PATTERN_i76_LC_11_18_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i76_LC_11_18_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i76_LC_11_18_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i76_LC_11_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9697),
            .lcout(\transmit_module.Y_DELTA_PATTERN_76 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22437),
            .ce(N__16038),
            .sr(N__21252));
    defparam \transmit_module.Y_DELTA_PATTERN_i72_LC_11_18_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i72_LC_11_18_7 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i72_LC_11_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i72_LC_11_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9727),
            .lcout(\transmit_module.Y_DELTA_PATTERN_72 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22437),
            .ce(N__16038),
            .sr(N__21252));
    defparam \transmit_module.Y_DELTA_PATTERN_i75_LC_11_19_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i75_LC_11_19_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i75_LC_11_19_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i75_LC_11_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9733),
            .lcout(\transmit_module.Y_DELTA_PATTERN_75 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22434),
            .ce(N__21463),
            .sr(N__21093));
    defparam \transmit_module.Y_DELTA_PATTERN_i73_LC_11_19_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i73_LC_11_19_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i73_LC_11_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i73_LC_11_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9703),
            .lcout(\transmit_module.Y_DELTA_PATTERN_73 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22434),
            .ce(N__21463),
            .sr(N__21093));
    defparam \transmit_module.Y_DELTA_PATTERN_i81_LC_11_19_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i81_LC_11_19_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i81_LC_11_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i81_LC_11_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9721),
            .lcout(\transmit_module.Y_DELTA_PATTERN_81 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22434),
            .ce(N__21463),
            .sr(N__21093));
    defparam \transmit_module.Y_DELTA_PATTERN_i74_LC_11_19_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i74_LC_11_19_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i74_LC_11_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i74_LC_11_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9709),
            .lcout(\transmit_module.Y_DELTA_PATTERN_74 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22434),
            .ce(N__21463),
            .sr(N__21093));
    defparam \transmit_module.Y_DELTA_PATTERN_i77_LC_11_19_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i77_LC_11_19_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i77_LC_11_19_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i77_LC_11_19_7  (
            .in0(N__10969),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.Y_DELTA_PATTERN_77 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22434),
            .ce(N__21463),
            .sr(N__21093));
    defparam ADV_R__i1_LC_11_20_2.C_ON=1'b0;
    defparam ADV_R__i1_LC_11_20_2.SEQ_MODE=4'b1000;
    defparam ADV_R__i1_LC_11_20_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 ADV_R__i1_LC_11_20_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22960),
            .lcout(n1996),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVADV_R__i1C_net),
            .ce(),
            .sr(N__14604));
    defparam \transmit_module.Y_DELTA_PATTERN_i63_LC_11_21_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i63_LC_11_21_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i63_LC_11_21_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i63_LC_11_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10636),
            .lcout(\transmit_module.Y_DELTA_PATTERN_63 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22439),
            .ce(N__21458),
            .sr(N__21092));
    defparam \transmit_module.Y_DELTA_PATTERN_i70_LC_11_21_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i70_LC_11_21_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i70_LC_11_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i70_LC_11_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9991),
            .lcout(\transmit_module.Y_DELTA_PATTERN_70 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22439),
            .ce(N__21458),
            .sr(N__21092));
    defparam \transmit_module.Y_DELTA_PATTERN_i69_LC_11_21_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i69_LC_11_21_2 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i69_LC_11_21_2 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i69_LC_11_21_2  (
            .in0(_gnd_net_),
            .in1(N__10006),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.Y_DELTA_PATTERN_69 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22439),
            .ce(N__21458),
            .sr(N__21092));
    defparam \transmit_module.Y_DELTA_PATTERN_i71_LC_11_21_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i71_LC_11_21_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i71_LC_11_21_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i71_LC_11_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10000),
            .lcout(\transmit_module.Y_DELTA_PATTERN_71 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22439),
            .ce(N__21458),
            .sr(N__21092));
    defparam \transmit_module.Y_DELTA_PATTERN_i62_LC_11_21_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i62_LC_11_21_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i62_LC_11_21_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i62_LC_11_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9985),
            .lcout(\transmit_module.Y_DELTA_PATTERN_62 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22439),
            .ce(N__21458),
            .sr(N__21092));
    defparam \transmit_module.i1773_4_lut_LC_11_31_7 .C_ON=1'b0;
    defparam \transmit_module.i1773_4_lut_LC_11_31_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1773_4_lut_LC_11_31_7 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \transmit_module.i1773_4_lut_LC_11_31_7  (
            .in0(N__11713),
            .in1(N__11725),
            .in2(N__21335),
            .in3(N__20245),
            .lcout(n18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i29_1_lut_LC_12_9_5 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i29_1_lut_LC_12_9_5 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i29_1_lut_LC_12_9_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \receive_module.rx_counter.i29_1_lut_LC_12_9_5  (
            .in0(N__17110),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\receive_module.rx_counter.PULSE_1HZ_N_97 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.i667_3_lut_4_lut_LC_12_10_0 .C_ON=1'b0;
    defparam \receive_module.i667_3_lut_4_lut_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \receive_module.i667_3_lut_4_lut_LC_12_10_0 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \receive_module.i667_3_lut_4_lut_LC_12_10_0  (
            .in0(N__12236),
            .in1(N__11987),
            .in2(N__12516),
            .in3(N__12545),
            .lcout(\receive_module.n5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.i1_2_lut_rep_21_3_lut_LC_12_10_1 .C_ON=1'b0;
    defparam \receive_module.i1_2_lut_rep_21_3_lut_LC_12_10_1 .SEQ_MODE=4'b0000;
    defparam \receive_module.i1_2_lut_rep_21_3_lut_LC_12_10_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \receive_module.i1_2_lut_rep_21_3_lut_LC_12_10_1  (
            .in0(N__12512),
            .in1(N__11986),
            .in2(_gnd_net_),
            .in3(N__12237),
            .lcout(),
            .ltout(\receive_module.n4212_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.i681_4_lut_LC_12_10_2 .C_ON=1'b0;
    defparam \receive_module.i681_4_lut_LC_12_10_2 .SEQ_MODE=4'b0000;
    defparam \receive_module.i681_4_lut_LC_12_10_2 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \receive_module.i681_4_lut_LC_12_10_2  (
            .in0(N__13221),
            .in1(N__12963),
            .in2(N__10132),
            .in3(N__12547),
            .lcout(\receive_module.n3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.i1_2_lut_rep_22_LC_12_10_3 .C_ON=1'b0;
    defparam \receive_module.i1_2_lut_rep_22_LC_12_10_3 .SEQ_MODE=4'b0000;
    defparam \receive_module.i1_2_lut_rep_22_LC_12_10_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \receive_module.i1_2_lut_rep_22_LC_12_10_3  (
            .in0(_gnd_net_),
            .in1(N__12506),
            .in2(_gnd_net_),
            .in3(N__12235),
            .lcout(),
            .ltout(\receive_module.n4213_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.i674_3_lut_4_lut_LC_12_10_4 .C_ON=1'b0;
    defparam \receive_module.i674_3_lut_4_lut_LC_12_10_4 .SEQ_MODE=4'b0000;
    defparam \receive_module.i674_3_lut_4_lut_LC_12_10_4 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \receive_module.i674_3_lut_4_lut_LC_12_10_4  (
            .in0(N__13220),
            .in1(N__11988),
            .in2(N__10129),
            .in3(N__12546),
            .lcout(\receive_module.n4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.i660_3_lut_LC_12_10_5 .C_ON=1'b0;
    defparam \receive_module.i660_3_lut_LC_12_10_5 .SEQ_MODE=4'b0000;
    defparam \receive_module.i660_3_lut_LC_12_10_5 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \receive_module.i660_3_lut_LC_12_10_5  (
            .in0(N__12544),
            .in1(N__12508),
            .in2(_gnd_net_),
            .in3(N__12234),
            .lcout(\receive_module.n6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.i652_2_lut_org_LC_12_10_6 .C_ON=1'b0;
    defparam \receive_module.i652_2_lut_org_LC_12_10_6 .SEQ_MODE=4'b0000;
    defparam \receive_module.i652_2_lut_org_LC_12_10_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \receive_module.i652_2_lut_org_LC_12_10_6  (
            .in0(N__12507),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12543),
            .lcout(\receive_module.n7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i1831_4_lut_LC_12_10_7 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i1831_4_lut_LC_12_10_7 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i1831_4_lut_LC_12_10_7 .LUT_INIT=16'b1010100010001000;
    LogicCell40 \receive_module.rx_counter.i1831_4_lut_LC_12_10_7  (
            .in0(N__17476),
            .in1(N__17503),
            .in2(N__12529),
            .in3(N__17416),
            .lcout(\receive_module.rx_counter.n3204 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i1_2_lut_4_lut_adj_18_LC_12_11_0 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i1_2_lut_4_lut_adj_18_LC_12_11_0 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i1_2_lut_4_lut_adj_18_LC_12_11_0 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \receive_module.rx_counter.i1_2_lut_4_lut_adj_18_LC_12_11_0  (
            .in0(N__15760),
            .in1(N__15928),
            .in2(N__15807),
            .in3(N__15886),
            .lcout(n659),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \db5.i2_2_lut_rep_30_LC_12_11_1 .C_ON=1'b0;
    defparam \db5.i2_2_lut_rep_30_LC_12_11_1 .SEQ_MODE=4'b0000;
    defparam \db5.i2_2_lut_rep_30_LC_12_11_1 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \db5.i2_2_lut_rep_30_LC_12_11_1  (
            .in0(N__13426),
            .in1(_gnd_net_),
            .in2(N__13393),
            .in3(_gnd_net_),
            .lcout(\db5.n4221 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \db5.CLK_EN_13_LC_12_11_2 .C_ON=1'b0;
    defparam \db5.CLK_EN_13_LC_12_11_2 .SEQ_MODE=4'b1000;
    defparam \db5.CLK_EN_13_LC_12_11_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \db5.CLK_EN_13_LC_12_11_2  (
            .in0(N__13326),
            .in1(N__13388),
            .in2(N__13363),
            .in3(N__13425),
            .lcout(DEBUG_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19335),
            .ce(),
            .sr(_gnd_net_));
    defparam \db5.COUNTER_i2_LC_12_11_3 .C_ON=1'b0;
    defparam \db5.COUNTER_i2_LC_12_11_3 .SEQ_MODE=4'b1000;
    defparam \db5.COUNTER_i2_LC_12_11_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \db5.COUNTER_i2_LC_12_11_3  (
            .in0(N__13389),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\db5.COUNTER_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19335),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i1_2_lut_4_lut_LC_12_11_4 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i1_2_lut_4_lut_LC_12_11_4 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i1_2_lut_4_lut_LC_12_11_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \receive_module.rx_counter.i1_2_lut_4_lut_LC_12_11_4  (
            .in0(N__15759),
            .in1(N__15927),
            .in2(N__15806),
            .in3(N__15885),
            .lcout(n691),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \db5.COUNTER_i0_LC_12_11_5 .C_ON=1'b0;
    defparam \db5.COUNTER_i0_LC_12_11_5 .SEQ_MODE=4'b1000;
    defparam \db5.COUNTER_i0_LC_12_11_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \db5.COUNTER_i0_LC_12_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13327),
            .lcout(\db5.COUNTER_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19335),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_11_LC_12_11_7 .C_ON=1'b0;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_11_LC_12_11_7 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_adj_11_LC_12_11_7 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \line_buffer.i1_2_lut_3_lut_4_lut_adj_11_LC_12_11_7  (
            .in0(N__15887),
            .in1(N__15795),
            .in2(N__15931),
            .in3(N__15758),
            .lcout(\line_buffer.n626 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \db5.COUNTER_i1_LC_12_12_5 .C_ON=1'b0;
    defparam \db5.COUNTER_i1_LC_12_12_5 .SEQ_MODE=4'b1000;
    defparam \db5.COUNTER_i1_LC_12_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \db5.COUNTER_i1_LC_12_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13356),
            .lcout(\db5.COUNTER_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19339),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1_3_lut_4_lut_adj_10_LC_12_12_6 .C_ON=1'b0;
    defparam \line_buffer.i1_3_lut_4_lut_adj_10_LC_12_12_6 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1_3_lut_4_lut_adj_10_LC_12_12_6 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \line_buffer.i1_3_lut_4_lut_adj_10_LC_12_12_6  (
            .in0(N__15929),
            .in1(N__15892),
            .in2(N__15848),
            .in3(N__15762),
            .lcout(\line_buffer.n561 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_2_lut_LC_12_14_0 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_2_lut_LC_12_14_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_2_lut_LC_12_14_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \transmit_module.video_signal_controller.i1_2_lut_LC_12_14_0  (
            .in0(_gnd_net_),
            .in1(N__13630),
            .in2(_gnd_net_),
            .in3(N__13603),
            .lcout(\transmit_module.video_signal_controller.n3917 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i3_4_lut_adj_14_LC_12_14_2 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i3_4_lut_adj_14_LC_12_14_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i3_4_lut_adj_14_LC_12_14_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \transmit_module.video_signal_controller.i3_4_lut_adj_14_LC_12_14_2  (
            .in0(N__13583),
            .in1(N__13559),
            .in2(N__13303),
            .in3(N__13604),
            .lcout(),
            .ltout(\transmit_module.video_signal_controller.n3978_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i2578_3_lut_LC_12_14_3 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i2578_3_lut_LC_12_14_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i2578_3_lut_LC_12_14_3 .LUT_INIT=16'b1111110011001100;
    LogicCell40 \transmit_module.video_signal_controller.i2578_3_lut_LC_12_14_3  (
            .in0(_gnd_net_),
            .in1(N__10450),
            .in2(N__10135),
            .in3(N__13536),
            .lcout(\transmit_module.video_signal_controller.n4052 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_25_LC_12_14_5 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_25_LC_12_14_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_25_LC_12_14_5 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \transmit_module.video_signal_controller.i1_2_lut_rep_25_LC_12_14_5  (
            .in0(N__13560),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13537),
            .lcout(),
            .ltout(\transmit_module.video_signal_controller.n4216_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.VGA_HS_60_LC_12_14_6 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.VGA_HS_60_LC_12_14_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_HS_60_LC_12_14_6 .LUT_INIT=16'b1110111011101111;
    LogicCell40 \transmit_module.video_signal_controller.VGA_HS_60_LC_12_14_6  (
            .in0(N__13513),
            .in1(N__10333),
            .in2(N__10327),
            .in3(N__10324),
            .lcout(ADV_HSYNC_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22620),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i570_3_lut_LC_12_14_7 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i570_3_lut_LC_12_14_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i570_3_lut_LC_12_14_7 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \transmit_module.video_signal_controller.i570_3_lut_LC_12_14_7  (
            .in0(N__13605),
            .in1(N__13633),
            .in2(_gnd_net_),
            .in3(N__13584),
            .lcout(\transmit_module.video_signal_controller.n12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1859_4_lut_LC_12_15_0 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1859_4_lut_LC_12_15_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1859_4_lut_LC_12_15_0 .LUT_INIT=16'b1111111111001000;
    LogicCell40 \transmit_module.video_signal_controller.i1859_4_lut_LC_12_15_0  (
            .in0(N__13837),
            .in1(N__13811),
            .in2(N__10309),
            .in3(N__13784),
            .lcout(\transmit_module.video_signal_controller.n2274 ),
            .ltout(\transmit_module.video_signal_controller.n2274_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1227_2_lut_LC_12_15_1 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1227_2_lut_LC_12_15_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1227_2_lut_LC_12_15_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \transmit_module.video_signal_controller.i1227_2_lut_LC_12_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10318),
            .in3(N__10315),
            .lcout(\transmit_module.video_signal_controller.n2594 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1853_4_lut_LC_12_15_2 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1853_4_lut_LC_12_15_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1853_4_lut_LC_12_15_2 .LUT_INIT=16'b1111100000000000;
    LogicCell40 \transmit_module.video_signal_controller.i1853_4_lut_LC_12_15_2  (
            .in0(N__10291),
            .in1(N__13294),
            .in2(N__10300),
            .in3(N__13508),
            .lcout(\transmit_module.video_signal_controller.n3226 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i560_2_lut_rep_26_LC_12_15_3 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i560_2_lut_rep_26_LC_12_15_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i560_2_lut_rep_26_LC_12_15_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \transmit_module.video_signal_controller.i560_2_lut_rep_26_LC_12_15_3  (
            .in0(_gnd_net_),
            .in1(N__13654),
            .in2(_gnd_net_),
            .in3(N__13681),
            .lcout(\transmit_module.video_signal_controller.n4217 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_2_lut_3_lut_adj_15_LC_12_15_4 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_2_lut_3_lut_adj_15_LC_12_15_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_2_lut_3_lut_adj_15_LC_12_15_4 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \transmit_module.video_signal_controller.i1_2_lut_3_lut_adj_15_LC_12_15_4  (
            .in0(N__13582),
            .in1(N__13558),
            .in2(_gnd_net_),
            .in3(N__13534),
            .lcout(\transmit_module.video_signal_controller.n2260 ),
            .ltout(\transmit_module.video_signal_controller.n2260_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i557_4_lut_LC_12_15_5 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i557_4_lut_LC_12_15_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i557_4_lut_LC_12_15_5 .LUT_INIT=16'b1010100010100000;
    LogicCell40 \transmit_module.video_signal_controller.i557_4_lut_LC_12_15_5  (
            .in0(N__13507),
            .in1(N__10290),
            .in2(N__10282),
            .in3(N__10279),
            .lcout(),
            .ltout(\transmit_module.video_signal_controller.n18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i2_4_lut_4_lut_LC_12_15_6 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i2_4_lut_4_lut_LC_12_15_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i2_4_lut_4_lut_LC_12_15_6 .LUT_INIT=16'b0000000000110110;
    LogicCell40 \transmit_module.video_signal_controller.i2_4_lut_4_lut_LC_12_15_6  (
            .in0(N__13835),
            .in1(N__13807),
            .in2(N__10453),
            .in3(N__13783),
            .lcout(\transmit_module.n3910 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i2_3_lut_LC_12_15_7 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i2_3_lut_LC_12_15_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i2_3_lut_LC_12_15_7 .LUT_INIT=16'b1111111111111010;
    LogicCell40 \transmit_module.video_signal_controller.i2_3_lut_LC_12_15_7  (
            .in0(N__13785),
            .in1(_gnd_net_),
            .in2(N__13813),
            .in3(N__13836),
            .lcout(\transmit_module.video_signal_controller.n2219 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.VGA_Y_i0_LC_12_16_0 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i0_LC_12_16_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i0_LC_12_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i0_LC_12_16_0  (
            .in0(_gnd_net_),
            .in1(N__10443),
            .in2(_gnd_net_),
            .in3(N__10432),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_0 ),
            .ltout(),
            .carryin(bfn_12_16_0_),
            .carryout(\transmit_module.video_signal_controller.n3677 ),
            .clk(N__22561),
            .ce(N__13761),
            .sr(N__10584));
    defparam \transmit_module.video_signal_controller.VGA_Y_i1_LC_12_16_1 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i1_LC_12_16_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i1_LC_12_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i1_LC_12_16_1  (
            .in0(_gnd_net_),
            .in1(N__10427),
            .in2(_gnd_net_),
            .in3(N__10405),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_1 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3677 ),
            .carryout(\transmit_module.video_signal_controller.n3678 ),
            .clk(N__22561),
            .ce(N__13761),
            .sr(N__10584));
    defparam \transmit_module.video_signal_controller.VGA_Y_i2_LC_12_16_2 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i2_LC_12_16_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i2_LC_12_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i2_LC_12_16_2  (
            .in0(_gnd_net_),
            .in1(N__10401),
            .in2(_gnd_net_),
            .in3(N__10381),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_2 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3678 ),
            .carryout(\transmit_module.video_signal_controller.n3679 ),
            .clk(N__22561),
            .ce(N__13761),
            .sr(N__10584));
    defparam \transmit_module.video_signal_controller.VGA_Y_i3_LC_12_16_3 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i3_LC_12_16_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i3_LC_12_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i3_LC_12_16_3  (
            .in0(_gnd_net_),
            .in1(N__10559),
            .in2(_gnd_net_),
            .in3(N__10378),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_3 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3679 ),
            .carryout(\transmit_module.video_signal_controller.n3680 ),
            .clk(N__22561),
            .ce(N__13761),
            .sr(N__10584));
    defparam \transmit_module.video_signal_controller.VGA_Y_i4_LC_12_16_4 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i4_LC_12_16_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i4_LC_12_16_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i4_LC_12_16_4  (
            .in0(_gnd_net_),
            .in1(N__10520),
            .in2(_gnd_net_),
            .in3(N__10375),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_4 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3680 ),
            .carryout(\transmit_module.video_signal_controller.n3681 ),
            .clk(N__22561),
            .ce(N__13761),
            .sr(N__10584));
    defparam \transmit_module.video_signal_controller.VGA_Y_i5_LC_12_16_5 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i5_LC_12_16_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i5_LC_12_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i5_LC_12_16_5  (
            .in0(_gnd_net_),
            .in1(N__10372),
            .in2(_gnd_net_),
            .in3(N__10354),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_5 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3681 ),
            .carryout(\transmit_module.video_signal_controller.n3682 ),
            .clk(N__22561),
            .ce(N__13761),
            .sr(N__10584));
    defparam \transmit_module.video_signal_controller.VGA_Y_i6_LC_12_16_6 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i6_LC_12_16_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i6_LC_12_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i6_LC_12_16_6  (
            .in0(_gnd_net_),
            .in1(N__10351),
            .in2(_gnd_net_),
            .in3(N__10336),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_6 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3682 ),
            .carryout(\transmit_module.video_signal_controller.n3683 ),
            .clk(N__22561),
            .ce(N__13761),
            .sr(N__10584));
    defparam \transmit_module.video_signal_controller.VGA_Y_i7_LC_12_16_7 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i7_LC_12_16_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i7_LC_12_16_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i7_LC_12_16_7  (
            .in0(_gnd_net_),
            .in1(N__10624),
            .in2(_gnd_net_),
            .in3(N__10612),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_7 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3683 ),
            .carryout(\transmit_module.video_signal_controller.n3684 ),
            .clk(N__22561),
            .ce(N__13761),
            .sr(N__10584));
    defparam \transmit_module.video_signal_controller.VGA_Y_i8_LC_12_17_0 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i8_LC_12_17_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i8_LC_12_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i8_LC_12_17_0  (
            .in0(_gnd_net_),
            .in1(N__10609),
            .in2(_gnd_net_),
            .in3(N__10597),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_8 ),
            .ltout(),
            .carryin(bfn_12_17_0_),
            .carryout(\transmit_module.video_signal_controller.n3685 ),
            .clk(N__22499),
            .ce(N__13768),
            .sr(N__10585));
    defparam \transmit_module.video_signal_controller.VGA_Y_i9_LC_12_17_1 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i9_LC_12_17_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i9_LC_12_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i9_LC_12_17_1  (
            .in0(_gnd_net_),
            .in1(N__10483),
            .in2(_gnd_net_),
            .in3(N__10594),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_9 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3685 ),
            .carryout(\transmit_module.video_signal_controller.n3686 ),
            .clk(N__22499),
            .ce(N__13768),
            .sr(N__10585));
    defparam \transmit_module.video_signal_controller.VGA_Y_i10_LC_12_17_2 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_Y_i10_LC_12_17_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i10_LC_12_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i10_LC_12_17_2  (
            .in0(_gnd_net_),
            .in1(N__10903),
            .in2(_gnd_net_),
            .in3(N__10591),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_10 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3686 ),
            .carryout(\transmit_module.video_signal_controller.n3687 ),
            .clk(N__22499),
            .ce(N__13768),
            .sr(N__10585));
    defparam \transmit_module.video_signal_controller.VGA_Y_i11_LC_12_17_3 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.VGA_Y_i11_LC_12_17_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_Y_i11_LC_12_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_Y_i11_LC_12_17_3  (
            .in0(_gnd_net_),
            .in1(N__10923),
            .in2(_gnd_net_),
            .in3(N__10588),
            .lcout(\transmit_module.video_signal_controller.VGA_Y_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22499),
            .ce(N__13768),
            .sr(N__10585));
    defparam \transmit_module.video_signal_controller.i1_4_lut_adj_13_LC_12_18_1 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_4_lut_adj_13_LC_12_18_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_4_lut_adj_13_LC_12_18_1 .LUT_INIT=16'b1111111111100000;
    LogicCell40 \transmit_module.video_signal_controller.i1_4_lut_adj_13_LC_12_18_1  (
            .in0(N__10561),
            .in1(N__10534),
            .in2(N__10528),
            .in3(N__10494),
            .lcout(),
            .ltout(\transmit_module.video_signal_controller.VGA_VISIBLE_Y_N_553_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i2_4_lut_adj_16_LC_12_18_2 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i2_4_lut_adj_16_LC_12_18_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i2_4_lut_adj_16_LC_12_18_2 .LUT_INIT=16'b0001000001010000;
    LogicCell40 \transmit_module.video_signal_controller.i2_4_lut_adj_16_LC_12_18_2  (
            .in0(N__10885),
            .in1(N__10482),
            .in2(N__10465),
            .in3(N__10462),
            .lcout(\transmit_module.n3926 ),
            .ltout(\transmit_module.n3926_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.mux_14_i3_3_lut_4_lut_LC_12_18_3 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.mux_14_i3_3_lut_4_lut_LC_12_18_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.mux_14_i3_3_lut_4_lut_LC_12_18_3 .LUT_INIT=16'b1010110011001100;
    LogicCell40 \transmit_module.video_signal_controller.mux_14_i3_3_lut_4_lut_LC_12_18_3  (
            .in0(N__17797),
            .in1(N__17822),
            .in2(N__10456),
            .in3(N__19100),
            .lcout(\transmit_module.n217 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_27_LC_12_18_6 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_27_LC_12_18_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_27_LC_12_18_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \transmit_module.video_signal_controller.i1_2_lut_rep_27_LC_12_18_6  (
            .in0(_gnd_net_),
            .in1(N__10922),
            .in2(_gnd_net_),
            .in3(N__10902),
            .lcout(\transmit_module.video_signal_controller.n4218 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1211_1_lut_2_lut_LC_12_19_0 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1211_1_lut_2_lut_LC_12_19_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1211_1_lut_2_lut_LC_12_19_0 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \transmit_module.video_signal_controller.i1211_1_lut_2_lut_LC_12_19_0  (
            .in0(_gnd_net_),
            .in1(N__19095),
            .in2(_gnd_net_),
            .in3(N__19467),
            .lcout(n2587),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.mux_14_i1_3_lut_4_lut_LC_12_19_2 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.mux_14_i1_3_lut_4_lut_LC_12_19_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.mux_14_i1_3_lut_4_lut_LC_12_19_2 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \transmit_module.video_signal_controller.mux_14_i1_3_lut_4_lut_LC_12_19_2  (
            .in0(N__18420),
            .in1(N__19099),
            .in2(N__17521),
            .in3(N__19468),
            .lcout(\transmit_module.n219 ),
            .ltout(\transmit_module.n219_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1757_4_lut_LC_12_19_3 .C_ON=1'b0;
    defparam \transmit_module.i1757_4_lut_LC_12_19_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1757_4_lut_LC_12_19_3 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \transmit_module.i1757_4_lut_LC_12_19_3  (
            .in0(N__20167),
            .in1(N__21036),
            .in2(N__10879),
            .in3(N__17839),
            .lcout(n28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_19_LC_12_19_5 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_19_LC_12_19_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_19_LC_12_19_5 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \transmit_module.video_signal_controller.i1_2_lut_rep_19_LC_12_19_5  (
            .in0(N__19469),
            .in1(_gnd_net_),
            .in2(N__19121),
            .in3(_gnd_net_),
            .lcout(n4210),
            .ltout(n4210_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1762_4_lut_LC_12_19_6 .C_ON=1'b0;
    defparam \transmit_module.i1762_4_lut_LC_12_19_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1762_4_lut_LC_12_19_6 .LUT_INIT=16'b1101110111111100;
    LogicCell40 \transmit_module.i1762_4_lut_LC_12_19_6  (
            .in0(N__19716),
            .in1(N__21037),
            .in2(N__10639),
            .in3(N__20166),
            .lcout(\transmit_module.n2277 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i13_LC_12_20_0 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i13_LC_12_20_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i13_LC_12_20_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \transmit_module.BRAM_ADDR__i13_LC_12_20_0  (
            .in0(N__22793),
            .in1(N__19150),
            .in2(_gnd_net_),
            .in3(N__19397),
            .lcout(DEBUG_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22534),
            .ce(),
            .sr(N__21167));
    defparam \transmit_module.Y_DELTA_PATTERN_i64_LC_12_21_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i64_LC_12_21_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i64_LC_12_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i64_LC_12_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10948),
            .lcout(\transmit_module.Y_DELTA_PATTERN_64 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22348),
            .ce(N__21456),
            .sr(N__21306));
    defparam \transmit_module.Y_DELTA_PATTERN_i66_LC_12_21_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i66_LC_12_21_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i66_LC_12_21_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i66_LC_12_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10630),
            .lcout(\transmit_module.Y_DELTA_PATTERN_66 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22348),
            .ce(N__21456),
            .sr(N__21306));
    defparam \transmit_module.Y_DELTA_PATTERN_i67_LC_12_21_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i67_LC_12_21_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i67_LC_12_21_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i67_LC_12_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10975),
            .lcout(\transmit_module.Y_DELTA_PATTERN_67 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22348),
            .ce(N__21456),
            .sr(N__21306));
    defparam \transmit_module.Y_DELTA_PATTERN_i80_LC_12_21_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i80_LC_12_21_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i80_LC_12_21_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i80_LC_12_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10993),
            .lcout(\transmit_module.Y_DELTA_PATTERN_80 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22348),
            .ce(N__21456),
            .sr(N__21306));
    defparam \transmit_module.Y_DELTA_PATTERN_i68_LC_12_21_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i68_LC_12_21_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i68_LC_12_21_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i68_LC_12_21_7  (
            .in0(N__10981),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.Y_DELTA_PATTERN_68 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22348),
            .ce(N__21456),
            .sr(N__21306));
    defparam \transmit_module.Y_DELTA_PATTERN_i78_LC_12_22_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i78_LC_12_22_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i78_LC_12_22_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i78_LC_12_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10936),
            .lcout(\transmit_module.Y_DELTA_PATTERN_78 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22315),
            .ce(N__21489),
            .sr(N__21278));
    defparam \transmit_module.Y_DELTA_PATTERN_i61_LC_12_22_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i61_LC_12_22_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i61_LC_12_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i61_LC_12_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10960),
            .lcout(\transmit_module.Y_DELTA_PATTERN_61 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22315),
            .ce(N__21489),
            .sr(N__21278));
    defparam \transmit_module.Y_DELTA_PATTERN_i51_LC_12_22_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i51_LC_12_22_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i51_LC_12_22_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i51_LC_12_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14545),
            .lcout(\transmit_module.Y_DELTA_PATTERN_51 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22315),
            .ce(N__21489),
            .sr(N__21278));
    defparam \transmit_module.Y_DELTA_PATTERN_i65_LC_12_22_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i65_LC_12_22_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i65_LC_12_22_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i65_LC_12_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10954),
            .lcout(\transmit_module.Y_DELTA_PATTERN_65 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22315),
            .ce(N__21489),
            .sr(N__21278));
    defparam \transmit_module.Y_DELTA_PATTERN_i79_LC_12_22_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i79_LC_12_22_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i79_LC_12_22_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i79_LC_12_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10942),
            .lcout(\transmit_module.Y_DELTA_PATTERN_79 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22315),
            .ce(N__21489),
            .sr(N__21278));
    defparam \transmit_module.Y_DELTA_PATTERN_i56_LC_12_23_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i56_LC_12_23_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i56_LC_12_23_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i56_LC_12_23_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10930),
            .lcout(\transmit_module.Y_DELTA_PATTERN_56 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21958),
            .ce(N__21493),
            .sr(N__21288));
    defparam \transmit_module.Y_DELTA_PATTERN_i57_LC_12_23_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i57_LC_12_23_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i57_LC_12_23_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i57_LC_12_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14656),
            .lcout(\transmit_module.Y_DELTA_PATTERN_57 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__21958),
            .ce(N__21493),
            .sr(N__21288));
    defparam \transmit_module.ADDR_Y_COMPONENT__i10_LC_12_24_6 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i10_LC_12_24_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i10_LC_12_24_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i10_LC_12_24_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17951),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22230),
            .ce(N__19881),
            .sr(N__21325));
    defparam \transmit_module.mux_12_i11_3_lut_LC_12_25_2 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i11_3_lut_LC_12_25_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i11_3_lut_LC_12_25_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_12_i11_3_lut_LC_12_25_2  (
            .in0(N__19717),
            .in1(N__11731),
            .in2(_gnd_net_),
            .in3(N__17944),
            .lcout(\transmit_module.n178 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.mux_14_i11_3_lut_4_lut_LC_12_26_1 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.mux_14_i11_3_lut_4_lut_LC_12_26_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.mux_14_i11_3_lut_4_lut_LC_12_26_1 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \transmit_module.video_signal_controller.mux_14_i11_3_lut_4_lut_LC_12_26_1  (
            .in0(N__17920),
            .in1(N__19129),
            .in2(N__17955),
            .in3(N__19520),
            .lcout(\transmit_module.n209 ),
            .ltout(\transmit_module.n209_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i10_LC_12_26_2 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i10_LC_12_26_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i10_LC_12_26_2 .LUT_INIT=16'b0010001000110000;
    LogicCell40 \transmit_module.BRAM_ADDR__i10_LC_12_26_2  (
            .in0(N__11709),
            .in1(N__21268),
            .in2(N__11695),
            .in3(N__20239),
            .lcout(\transmit_module.TX_ADDR_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22229),
            .ce(),
            .sr(_gnd_net_));
    defparam i284_3_lut_3_lut_LC_13_9_3.C_ON=1'b0;
    defparam i284_3_lut_3_lut_LC_13_9_3.SEQ_MODE=4'b0000;
    defparam i284_3_lut_3_lut_LC_13_9_3.LUT_INIT=16'b0111011101010101;
    LogicCell40 i284_3_lut_3_lut_LC_13_9_3 (
            .in0(N__17106),
            .in1(N__15441),
            .in2(_gnd_net_),
            .in3(N__11668),
            .lcout(n2283),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.old_HS_50_LC_13_9_6 .C_ON=1'b0;
    defparam \receive_module.rx_counter.old_HS_50_LC_13_9_6 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.old_HS_50_LC_13_9_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \receive_module.rx_counter.old_HS_50_LC_13_9_6  (
            .in0(N__15442),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(old_HS),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19329),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.sub_29_add_2_2_lut_LC_13_10_0 .C_ON=1'b1;
    defparam \receive_module.rx_counter.sub_29_add_2_2_lut_LC_13_10_0 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.sub_29_add_2_2_lut_LC_13_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.sub_29_add_2_2_lut_LC_13_10_0  (
            .in0(_gnd_net_),
            .in1(N__17026),
            .in2(_gnd_net_),
            .in3(N__11434),
            .lcout(RX_ADDR_3),
            .ltout(),
            .carryin(bfn_13_10_0_),
            .carryout(\receive_module.rx_counter.n3650 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.sub_29_add_2_3_lut_LC_13_10_1 .C_ON=1'b1;
    defparam \receive_module.rx_counter.sub_29_add_2_3_lut_LC_13_10_1 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.sub_29_add_2_3_lut_LC_13_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.sub_29_add_2_3_lut_LC_13_10_1  (
            .in0(_gnd_net_),
            .in1(N__17047),
            .in2(N__23303),
            .in3(N__11212),
            .lcout(RX_ADDR_4),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3650 ),
            .carryout(\receive_module.rx_counter.n3651 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.sub_29_add_2_4_lut_LC_13_10_2 .C_ON=1'b1;
    defparam \receive_module.rx_counter.sub_29_add_2_4_lut_LC_13_10_2 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.sub_29_add_2_4_lut_LC_13_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.sub_29_add_2_4_lut_LC_13_10_2  (
            .in0(_gnd_net_),
            .in1(N__23238),
            .in2(N__17074),
            .in3(N__10996),
            .lcout(RX_ADDR_5),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3651 ),
            .carryout(\receive_module.rx_counter.n3652 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.sub_29_add_2_5_lut_LC_13_10_3 .C_ON=1'b1;
    defparam \receive_module.rx_counter.sub_29_add_2_5_lut_LC_13_10_3 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.sub_29_add_2_5_lut_LC_13_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.sub_29_add_2_5_lut_LC_13_10_3  (
            .in0(_gnd_net_),
            .in1(N__17407),
            .in2(N__23304),
            .in3(N__12559),
            .lcout(\receive_module.O_X_6 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3652 ),
            .carryout(\receive_module.rx_counter.n3653 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.sub_29_add_2_6_lut_LC_13_10_4 .C_ON=1'b1;
    defparam \receive_module.rx_counter.sub_29_add_2_6_lut_LC_13_10_4 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.sub_29_add_2_6_lut_LC_13_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.sub_29_add_2_6_lut_LC_13_10_4  (
            .in0(_gnd_net_),
            .in1(N__17437),
            .in2(_gnd_net_),
            .in3(N__12556),
            .lcout(\receive_module.O_X_7 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3653 ),
            .carryout(\receive_module.rx_counter.n3654 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.sub_29_add_2_7_lut_LC_13_10_5 .C_ON=1'b1;
    defparam \receive_module.rx_counter.sub_29_add_2_7_lut_LC_13_10_5 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.sub_29_add_2_7_lut_LC_13_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.sub_29_add_2_7_lut_LC_13_10_5  (
            .in0(_gnd_net_),
            .in1(N__17497),
            .in2(N__23305),
            .in3(N__12553),
            .lcout(\receive_module.O_X_8 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3654 ),
            .carryout(\receive_module.rx_counter.n3655 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.sub_29_add_2_8_lut_LC_13_10_6 .C_ON=1'b0;
    defparam \receive_module.rx_counter.sub_29_add_2_8_lut_LC_13_10_6 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.sub_29_add_2_8_lut_LC_13_10_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \receive_module.rx_counter.sub_29_add_2_8_lut_LC_13_10_6  (
            .in0(N__17470),
            .in1(N__23245),
            .in2(_gnd_net_),
            .in3(N__12550),
            .lcout(\receive_module.O_X_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i1_2_lut_4_lut_adj_19_LC_13_10_7 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i1_2_lut_4_lut_adj_19_LC_13_10_7 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i1_2_lut_4_lut_adj_19_LC_13_10_7 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \receive_module.rx_counter.i1_2_lut_4_lut_adj_19_LC_13_10_7  (
            .in0(N__17027),
            .in1(N__17071),
            .in2(N__17443),
            .in3(N__17048),
            .lcout(\receive_module.rx_counter.n4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_629_2_lut_LC_13_11_0 .C_ON=1'b1;
    defparam \receive_module.add_629_2_lut_LC_13_11_0 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_629_2_lut_LC_13_11_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_629_2_lut_LC_13_11_0  (
            .in0(_gnd_net_),
            .in1(N__12520),
            .in2(N__12484),
            .in3(_gnd_net_),
            .lcout(RX_ADDR_6),
            .ltout(),
            .carryin(bfn_13_11_0_),
            .carryout(\receive_module.n3699 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_629_3_lut_LC_13_11_1 .C_ON=1'b1;
    defparam \receive_module.add_629_3_lut_LC_13_11_1 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_629_3_lut_LC_13_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_629_3_lut_LC_13_11_1  (
            .in0(_gnd_net_),
            .in1(N__12250),
            .in2(N__12244),
            .in3(N__11998),
            .lcout(RX_ADDR_7),
            .ltout(),
            .carryin(\receive_module.n3699 ),
            .carryout(\receive_module.n3700 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_629_4_lut_LC_13_11_2 .C_ON=1'b1;
    defparam \receive_module.add_629_4_lut_LC_13_11_2 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_629_4_lut_LC_13_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_629_4_lut_LC_13_11_2  (
            .in0(_gnd_net_),
            .in1(N__11995),
            .in2(N__11968),
            .in3(N__11734),
            .lcout(RX_ADDR_8),
            .ltout(),
            .carryin(\receive_module.n3700 ),
            .carryout(\receive_module.n3701 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_629_5_lut_LC_13_11_3 .C_ON=1'b1;
    defparam \receive_module.add_629_5_lut_LC_13_11_3 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_629_5_lut_LC_13_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_629_5_lut_LC_13_11_3  (
            .in0(_gnd_net_),
            .in1(N__13237),
            .in2(N__13231),
            .in3(N__12982),
            .lcout(RX_ADDR_9),
            .ltout(),
            .carryin(\receive_module.n3701 ),
            .carryout(\receive_module.n3702 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_629_6_lut_LC_13_11_4 .C_ON=1'b1;
    defparam \receive_module.add_629_6_lut_LC_13_11_4 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_629_6_lut_LC_13_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_629_6_lut_LC_13_11_4  (
            .in0(_gnd_net_),
            .in1(N__12979),
            .in2(N__12973),
            .in3(N__12730),
            .lcout(RX_ADDR_10),
            .ltout(),
            .carryin(\receive_module.n3702 ),
            .carryout(\receive_module.n3703 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_629_7_lut_LC_13_11_5 .C_ON=1'b1;
    defparam \receive_module.add_629_7_lut_LC_13_11_5 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_629_7_lut_LC_13_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_629_7_lut_LC_13_11_5  (
            .in0(_gnd_net_),
            .in1(N__12727),
            .in2(N__12721),
            .in3(N__12706),
            .lcout(RX_ADDR_11),
            .ltout(),
            .carryin(\receive_module.n3703 ),
            .carryout(\receive_module.n3704 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_629_8_lut_LC_13_11_6 .C_ON=1'b1;
    defparam \receive_module.add_629_8_lut_LC_13_11_6 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_629_8_lut_LC_13_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.add_629_8_lut_LC_13_11_6  (
            .in0(_gnd_net_),
            .in1(N__12703),
            .in2(N__12697),
            .in3(N__12682),
            .lcout(RX_ADDR_12),
            .ltout(),
            .carryin(\receive_module.n3704 ),
            .carryout(\receive_module.n3705 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.add_629_9_lut_LC_13_11_7 .C_ON=1'b0;
    defparam \receive_module.add_629_9_lut_LC_13_11_7 .SEQ_MODE=4'b0000;
    defparam \receive_module.add_629_9_lut_LC_13_11_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \receive_module.add_629_9_lut_LC_13_11_7  (
            .in0(N__12679),
            .in1(N__12673),
            .in2(_gnd_net_),
            .in3(N__12661),
            .lcout(DEBUG_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_LC_13_12_0 .C_ON=1'b0;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_LC_13_12_0 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1_2_lut_3_lut_4_lut_LC_13_12_0 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \line_buffer.i1_2_lut_3_lut_4_lut_LC_13_12_0  (
            .in0(N__15923),
            .in1(N__15889),
            .in2(N__15843),
            .in3(N__15755),
            .lcout(\line_buffer.n627 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i1_3_lut_4_lut_LC_13_12_2 .C_ON=1'b0;
    defparam \line_buffer.i1_3_lut_4_lut_LC_13_12_2 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i1_3_lut_4_lut_LC_13_12_2 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \line_buffer.i1_3_lut_4_lut_LC_13_12_2  (
            .in0(N__15922),
            .in1(N__15890),
            .in2(N__15844),
            .in3(N__15756),
            .lcout(\line_buffer.n562 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \db5.COUNTER_i3_LC_13_12_5 .C_ON=1'b0;
    defparam \db5.COUNTER_i3_LC_13_12_5 .SEQ_MODE=4'b1000;
    defparam \db5.COUNTER_i3_LC_13_12_5 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \db5.COUNTER_i3_LC_13_12_5  (
            .in0(_gnd_net_),
            .in1(N__13424),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\db5.COUNTER_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19336),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i1_2_lut_4_lut_adj_22_LC_13_12_6 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i1_2_lut_4_lut_adj_22_LC_13_12_6 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i1_2_lut_4_lut_adj_22_LC_13_12_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \receive_module.rx_counter.i1_2_lut_4_lut_adj_22_LC_13_12_6  (
            .in0(N__15921),
            .in1(N__15888),
            .in2(N__15842),
            .in3(N__15757),
            .lcout(n690),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \db5.NEXT_COUNTER__i3_LC_13_13_0 .C_ON=1'b0;
    defparam \db5.NEXT_COUNTER__i3_LC_13_13_0 .SEQ_MODE=4'b1000;
    defparam \db5.NEXT_COUNTER__i3_LC_13_13_0 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \db5.NEXT_COUNTER__i3_LC_13_13_0  (
            .in0(N__13345),
            .in1(N__13408),
            .in2(N__13435),
            .in3(N__13375),
            .lcout(\db5.NEXT_COUNTER_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVdb5.NEXT_COUNTER__i3C_net ),
            .ce(),
            .sr(N__13315));
    defparam \db5.NEXT_COUNTER__i2_LC_13_13_1 .C_ON=1'b0;
    defparam \db5.NEXT_COUNTER__i2_LC_13_13_1 .SEQ_MODE=4'b1000;
    defparam \db5.NEXT_COUNTER__i2_LC_13_13_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \db5.NEXT_COUNTER__i2_LC_13_13_1  (
            .in0(N__13374),
            .in1(N__13407),
            .in2(_gnd_net_),
            .in3(N__13344),
            .lcout(\db5.NEXT_COUNTER_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVdb5.NEXT_COUNTER__i3C_net ),
            .ce(),
            .sr(N__13315));
    defparam \db5.NEXT_COUNTER__i1_LC_13_13_2 .C_ON=1'b0;
    defparam \db5.NEXT_COUNTER__i1_LC_13_13_2 .SEQ_MODE=4'b1000;
    defparam \db5.NEXT_COUNTER__i1_LC_13_13_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \db5.NEXT_COUNTER__i1_LC_13_13_2  (
            .in0(N__13343),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13373),
            .lcout(\db5.NEXT_COUNTER_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVdb5.NEXT_COUNTER__i3C_net ),
            .ce(),
            .sr(N__13315));
    defparam \db5.NEXT_COUNTER__i0_LC_13_13_3 .C_ON=1'b0;
    defparam \db5.NEXT_COUNTER__i0_LC_13_13_3 .SEQ_MODE=4'b1000;
    defparam \db5.NEXT_COUNTER__i0_LC_13_13_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \db5.NEXT_COUNTER__i0_LC_13_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13342),
            .lcout(\db5.NEXT_COUNTER_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVdb5.NEXT_COUNTER__i3C_net ),
            .ce(),
            .sr(N__13315));
    defparam \transmit_module.video_signal_controller.i2_4_lut_LC_13_14_0 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i2_4_lut_LC_13_14_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i2_4_lut_LC_13_14_0 .LUT_INIT=16'b1100000010000000;
    LogicCell40 \transmit_module.video_signal_controller.i2_4_lut_LC_13_14_0  (
            .in0(N__13683),
            .in1(N__13631),
            .in2(N__13660),
            .in3(N__13254),
            .lcout(\transmit_module.video_signal_controller.n3997 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1823_2_lut_3_lut_LC_13_14_1 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1823_2_lut_3_lut_LC_13_14_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1823_2_lut_3_lut_LC_13_14_1 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \transmit_module.video_signal_controller.i1823_2_lut_3_lut_LC_13_14_1  (
            .in0(N__13253),
            .in1(N__13655),
            .in2(_gnd_net_),
            .in3(N__13682),
            .lcout(\transmit_module.video_signal_controller.n3196 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2628_3_lut_LC_13_14_5 .C_ON=1'b0;
    defparam \line_buffer.i2628_3_lut_LC_13_14_5 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2628_3_lut_LC_13_14_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \line_buffer.i2628_3_lut_LC_13_14_5  (
            .in0(N__13288),
            .in1(N__13270),
            .in2(_gnd_net_),
            .in3(N__23591),
            .lcout(\line_buffer.n4102 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.VGA_X_i0_LC_13_15_0 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i0_LC_13_15_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i0_LC_13_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i0_LC_13_15_0  (
            .in0(_gnd_net_),
            .in1(N__13255),
            .in2(_gnd_net_),
            .in3(N__13240),
            .lcout(\transmit_module.video_signal_controller.VGA_X_0 ),
            .ltout(),
            .carryin(bfn_13_15_0_),
            .carryout(\transmit_module.video_signal_controller.n3688 ),
            .clk(N__22422),
            .ce(),
            .sr(N__13753));
    defparam \transmit_module.video_signal_controller.VGA_X_i1_LC_13_15_1 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i1_LC_13_15_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i1_LC_13_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i1_LC_13_15_1  (
            .in0(_gnd_net_),
            .in1(N__13684),
            .in2(_gnd_net_),
            .in3(N__13663),
            .lcout(\transmit_module.video_signal_controller.VGA_X_1 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3688 ),
            .carryout(\transmit_module.video_signal_controller.n3689 ),
            .clk(N__22422),
            .ce(),
            .sr(N__13753));
    defparam \transmit_module.video_signal_controller.VGA_X_i2_LC_13_15_2 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i2_LC_13_15_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i2_LC_13_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i2_LC_13_15_2  (
            .in0(_gnd_net_),
            .in1(N__13659),
            .in2(_gnd_net_),
            .in3(N__13636),
            .lcout(\transmit_module.video_signal_controller.VGA_X_2 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3689 ),
            .carryout(\transmit_module.video_signal_controller.n3690 ),
            .clk(N__22422),
            .ce(),
            .sr(N__13753));
    defparam \transmit_module.video_signal_controller.VGA_X_i3_LC_13_15_3 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i3_LC_13_15_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i3_LC_13_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i3_LC_13_15_3  (
            .in0(_gnd_net_),
            .in1(N__13632),
            .in2(_gnd_net_),
            .in3(N__13609),
            .lcout(\transmit_module.video_signal_controller.VGA_X_3 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3690 ),
            .carryout(\transmit_module.video_signal_controller.n3691 ),
            .clk(N__22422),
            .ce(),
            .sr(N__13753));
    defparam \transmit_module.video_signal_controller.VGA_X_i4_LC_13_15_4 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i4_LC_13_15_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i4_LC_13_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i4_LC_13_15_4  (
            .in0(_gnd_net_),
            .in1(N__13606),
            .in2(_gnd_net_),
            .in3(N__13588),
            .lcout(\transmit_module.video_signal_controller.VGA_X_4 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3691 ),
            .carryout(\transmit_module.video_signal_controller.n3692 ),
            .clk(N__22422),
            .ce(),
            .sr(N__13753));
    defparam \transmit_module.video_signal_controller.VGA_X_i5_LC_13_15_5 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i5_LC_13_15_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i5_LC_13_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i5_LC_13_15_5  (
            .in0(_gnd_net_),
            .in1(N__13585),
            .in2(_gnd_net_),
            .in3(N__13564),
            .lcout(\transmit_module.video_signal_controller.VGA_X_5 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3692 ),
            .carryout(\transmit_module.video_signal_controller.n3693 ),
            .clk(N__22422),
            .ce(),
            .sr(N__13753));
    defparam \transmit_module.video_signal_controller.VGA_X_i6_LC_13_15_6 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i6_LC_13_15_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i6_LC_13_15_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i6_LC_13_15_6  (
            .in0(_gnd_net_),
            .in1(N__13561),
            .in2(_gnd_net_),
            .in3(N__13540),
            .lcout(\transmit_module.video_signal_controller.VGA_X_6 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3693 ),
            .carryout(\transmit_module.video_signal_controller.n3694 ),
            .clk(N__22422),
            .ce(),
            .sr(N__13753));
    defparam \transmit_module.video_signal_controller.VGA_X_i7_LC_13_15_7 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i7_LC_13_15_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i7_LC_13_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i7_LC_13_15_7  (
            .in0(_gnd_net_),
            .in1(N__13535),
            .in2(_gnd_net_),
            .in3(N__13516),
            .lcout(\transmit_module.video_signal_controller.VGA_X_7 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3694 ),
            .carryout(\transmit_module.video_signal_controller.n3695 ),
            .clk(N__22422),
            .ce(),
            .sr(N__13753));
    defparam \transmit_module.video_signal_controller.VGA_X_i8_LC_13_16_0 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i8_LC_13_16_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i8_LC_13_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i8_LC_13_16_0  (
            .in0(_gnd_net_),
            .in1(N__13509),
            .in2(_gnd_net_),
            .in3(N__13489),
            .lcout(\transmit_module.video_signal_controller.VGA_X_8 ),
            .ltout(),
            .carryin(bfn_13_16_0_),
            .carryout(\transmit_module.video_signal_controller.n3696 ),
            .clk(N__22609),
            .ce(),
            .sr(N__13754));
    defparam \transmit_module.video_signal_controller.VGA_X_i9_LC_13_16_1 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i9_LC_13_16_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i9_LC_13_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i9_LC_13_16_1  (
            .in0(_gnd_net_),
            .in1(N__13834),
            .in2(_gnd_net_),
            .in3(N__13816),
            .lcout(\transmit_module.video_signal_controller.VGA_X_9 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3696 ),
            .carryout(\transmit_module.video_signal_controller.n3697 ),
            .clk(N__22609),
            .ce(),
            .sr(N__13754));
    defparam \transmit_module.video_signal_controller.VGA_X_i10_LC_13_16_2 .C_ON=1'b1;
    defparam \transmit_module.video_signal_controller.VGA_X_i10_LC_13_16_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i10_LC_13_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i10_LC_13_16_2  (
            .in0(_gnd_net_),
            .in1(N__13812),
            .in2(_gnd_net_),
            .in3(N__13792),
            .lcout(\transmit_module.video_signal_controller.VGA_X_10 ),
            .ltout(),
            .carryin(\transmit_module.video_signal_controller.n3697 ),
            .carryout(\transmit_module.video_signal_controller.n3698 ),
            .clk(N__22609),
            .ce(),
            .sr(N__13754));
    defparam \transmit_module.video_signal_controller.VGA_X_i11_LC_13_16_3 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.VGA_X_i11_LC_13_16_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.video_signal_controller.VGA_X_i11_LC_13_16_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.video_signal_controller.VGA_X_i11_LC_13_16_3  (
            .in0(_gnd_net_),
            .in1(N__13786),
            .in2(_gnd_net_),
            .in3(N__13789),
            .lcout(\transmit_module.video_signal_controller.VGA_X_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22609),
            .ce(),
            .sr(N__13754));
    defparam \transmit_module.video_signal_controller.mux_14_i7_3_lut_4_lut_LC_13_17_1 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.mux_14_i7_3_lut_4_lut_LC_13_17_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.mux_14_i7_3_lut_4_lut_LC_13_17_1 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \transmit_module.video_signal_controller.mux_14_i7_3_lut_4_lut_LC_13_17_1  (
            .in0(N__17725),
            .in1(N__19101),
            .in2(N__17756),
            .in3(N__19500),
            .lcout(\transmit_module.n213 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i2_LC_13_17_3 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i2_LC_13_17_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i2_LC_13_17_3 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \transmit_module.BRAM_ADDR__i2_LC_13_17_3  (
            .in0(N__14122),
            .in1(N__14107),
            .in2(N__21259),
            .in3(N__20215),
            .lcout(\transmit_module.TX_ADDR_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22533),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i6_LC_13_17_5 .C_ON=1'b0;
    defparam \line_buffer.dout_i6_LC_13_17_5 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i6_LC_13_17_5 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \line_buffer.dout_i6_LC_13_17_5  (
            .in0(N__13726),
            .in1(N__22829),
            .in2(N__15670),
            .in3(N__16051),
            .lcout(TX_DATA_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22533),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i143_2_lut_3_lut_4_lut_LC_13_17_6 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i143_2_lut_3_lut_4_lut_LC_13_17_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i143_2_lut_3_lut_4_lut_LC_13_17_6 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \transmit_module.video_signal_controller.i143_2_lut_3_lut_4_lut_LC_13_17_6  (
            .in0(N__19501),
            .in1(N__16762),
            .in2(N__21219),
            .in3(N__16705),
            .lcout(\transmit_module.n2361 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2703_LC_13_17_7 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2703_LC_13_17_7 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2703_LC_13_17_7 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_2703_LC_13_17_7  (
            .in0(N__13717),
            .in1(N__23807),
            .in2(N__13702),
            .in3(N__23576),
            .lcout(\line_buffer.n4182 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.mux_14_i9_3_lut_4_lut_LC_13_18_1 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.mux_14_i9_3_lut_4_lut_LC_13_18_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.mux_14_i9_3_lut_4_lut_LC_13_18_1 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \transmit_module.video_signal_controller.mux_14_i9_3_lut_4_lut_LC_13_18_1  (
            .in0(N__17668),
            .in1(N__19103),
            .in2(N__17893),
            .in3(N__19494),
            .lcout(\transmit_module.n211 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.mux_14_i8_3_lut_4_lut_LC_13_18_2 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.mux_14_i8_3_lut_4_lut_LC_13_18_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.mux_14_i8_3_lut_4_lut_LC_13_18_2 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \transmit_module.video_signal_controller.mux_14_i8_3_lut_4_lut_LC_13_18_2  (
            .in0(N__19493),
            .in1(N__17683),
            .in2(N__17712),
            .in3(N__19104),
            .lcout(\transmit_module.n212 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i3_3_lut_LC_13_18_3 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i3_3_lut_LC_13_18_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i3_3_lut_LC_13_18_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_12_i3_3_lut_LC_13_18_3  (
            .in0(N__19714),
            .in1(N__16366),
            .in2(_gnd_net_),
            .in3(N__17821),
            .lcout(\transmit_module.n186 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_3_lut_4_lut_LC_13_18_4 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_3_lut_4_lut_LC_13_18_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_3_lut_4_lut_LC_13_18_4 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \transmit_module.video_signal_controller.i1_3_lut_4_lut_LC_13_18_4  (
            .in0(N__19496),
            .in1(N__19715),
            .in2(N__21196),
            .in3(N__19572),
            .lcout(\transmit_module.n2305 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.mux_14_i10_3_lut_4_lut_LC_13_18_5 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.mux_14_i10_3_lut_4_lut_LC_13_18_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.mux_14_i10_3_lut_4_lut_LC_13_18_5 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \transmit_module.video_signal_controller.mux_14_i10_3_lut_4_lut_LC_13_18_5  (
            .in0(N__17653),
            .in1(N__19102),
            .in2(N__18465),
            .in3(N__19492),
            .lcout(\transmit_module.n210 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i143_2_lut_3_lut_4_lut_rep_34_LC_13_18_6 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i143_2_lut_3_lut_4_lut_rep_34_LC_13_18_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i143_2_lut_3_lut_4_lut_rep_34_LC_13_18_6 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \transmit_module.video_signal_controller.i143_2_lut_3_lut_4_lut_rep_34_LC_13_18_6  (
            .in0(N__19495),
            .in1(N__16761),
            .in2(N__21195),
            .in3(N__16717),
            .lcout(\transmit_module.n4225 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i9_3_lut_LC_13_19_1 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i9_3_lut_LC_13_19_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i9_3_lut_LC_13_19_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \transmit_module.mux_12_i9_3_lut_LC_13_19_1  (
            .in0(N__17886),
            .in1(N__19692),
            .in2(_gnd_net_),
            .in3(N__17866),
            .lcout(\transmit_module.n180 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_20_3_lut_LC_13_19_2 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_20_3_lut_LC_13_19_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_20_3_lut_LC_13_19_2 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \transmit_module.video_signal_controller.i1_2_lut_rep_20_3_lut_LC_13_19_2  (
            .in0(N__16712),
            .in1(N__16756),
            .in2(_gnd_net_),
            .in3(N__19470),
            .lcout(\transmit_module.n4211 ),
            .ltout(\transmit_module.n4211_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1765_4_lut_LC_13_19_3 .C_ON=1'b0;
    defparam \transmit_module.i1765_4_lut_LC_13_19_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1765_4_lut_LC_13_19_3 .LUT_INIT=16'b0100010101000000;
    LogicCell40 \transmit_module.i1765_4_lut_LC_13_19_3  (
            .in0(N__21035),
            .in1(N__14121),
            .in2(N__14110),
            .in3(N__14106),
            .lcout(n26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.mux_14_i4_3_lut_4_lut_LC_13_19_4 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.mux_14_i4_3_lut_4_lut_LC_13_19_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.mux_14_i4_3_lut_4_lut_LC_13_19_4 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \transmit_module.video_signal_controller.mux_14_i4_3_lut_4_lut_LC_13_19_4  (
            .in0(N__18375),
            .in1(N__19122),
            .in2(N__17782),
            .in3(N__19471),
            .lcout(\transmit_module.n216 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n4182_bdd_4_lut_LC_13_19_5 .C_ON=1'b0;
    defparam \line_buffer.n4182_bdd_4_lut_LC_13_19_5 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n4182_bdd_4_lut_LC_13_19_5 .LUT_INIT=16'b1100110010111000;
    LogicCell40 \line_buffer.n4182_bdd_4_lut_LC_13_19_5  (
            .in0(N__13876),
            .in1(N__13861),
            .in2(N__13852),
            .in3(N__23855),
            .lcout(),
            .ltout(\line_buffer.n4185_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i7_LC_13_19_6 .C_ON=1'b0;
    defparam \line_buffer.dout_i7_LC_13_19_6 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i7_LC_13_19_6 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \line_buffer.dout_i7_LC_13_19_6  (
            .in0(_gnd_net_),
            .in1(N__22764),
            .in2(N__14539),
            .in3(N__14536),
            .lcout(TX_DATA_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22266),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.old_VGA_HS_34_LC_13_19_7 .C_ON=1'b0;
    defparam \transmit_module.old_VGA_HS_34_LC_13_19_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.old_VGA_HS_34_LC_13_19_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.old_VGA_HS_34_LC_13_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16713),
            .lcout(\transmit_module.old_VGA_HS ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22266),
            .ce(),
            .sr(_gnd_net_));
    defparam ADV_R__i2_LC_13_20_1.C_ON=1'b0;
    defparam ADV_R__i2_LC_13_20_1.SEQ_MODE=4'b1000;
    defparam ADV_R__i2_LC_13_20_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 ADV_R__i2_LC_13_20_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20404),
            .lcout(n1995),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVADV_R__i2C_net),
            .ce(),
            .sr(N__14605));
    defparam ADV_R__i3_LC_13_20_2.C_ON=1'b0;
    defparam ADV_R__i3_LC_13_20_2.SEQ_MODE=4'b1000;
    defparam ADV_R__i3_LC_13_20_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 ADV_R__i3_LC_13_20_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14479),
            .lcout(n1994),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVADV_R__i2C_net),
            .ce(),
            .sr(N__14605));
    defparam ADV_R__i4_LC_13_20_3.C_ON=1'b0;
    defparam ADV_R__i4_LC_13_20_3.SEQ_MODE=4'b1000;
    defparam ADV_R__i4_LC_13_20_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 ADV_R__i4_LC_13_20_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21580),
            .lcout(n1993),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVADV_R__i2C_net),
            .ce(),
            .sr(N__14605));
    defparam ADV_R__i5_LC_13_20_4.C_ON=1'b0;
    defparam ADV_R__i5_LC_13_20_4.SEQ_MODE=4'b1000;
    defparam ADV_R__i5_LC_13_20_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 ADV_R__i5_LC_13_20_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22708),
            .lcout(n1992),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVADV_R__i2C_net),
            .ce(),
            .sr(N__14605));
    defparam ADV_R__i6_LC_13_20_5.C_ON=1'b0;
    defparam ADV_R__i6_LC_13_20_5.SEQ_MODE=4'b1000;
    defparam ADV_R__i6_LC_13_20_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 ADV_R__i6_LC_13_20_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17971),
            .lcout(n1991),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVADV_R__i2C_net),
            .ce(),
            .sr(N__14605));
    defparam ADV_R__i7_LC_13_20_6.C_ON=1'b0;
    defparam ADV_R__i7_LC_13_20_6.SEQ_MODE=4'b1000;
    defparam ADV_R__i7_LC_13_20_6.LUT_INIT=16'b1010101010101010;
    LogicCell40 ADV_R__i7_LC_13_20_6 (
            .in0(N__14254),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n1990),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVADV_R__i2C_net),
            .ce(),
            .sr(N__14605));
    defparam ADV_R__i8_LC_13_20_7.C_ON=1'b0;
    defparam ADV_R__i8_LC_13_20_7.SEQ_MODE=4'b1000;
    defparam ADV_R__i8_LC_13_20_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 ADV_R__i8_LC_13_20_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14188),
            .lcout(ADV_B_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVADV_R__i2C_net),
            .ce(),
            .sr(N__14605));
    defparam \transmit_module.Y_DELTA_PATTERN_i42_LC_13_21_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i42_LC_13_21_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i42_LC_13_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i42_LC_13_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14587),
            .lcout(\transmit_module.Y_DELTA_PATTERN_42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22486),
            .ce(N__21436),
            .sr(N__21344));
    defparam \transmit_module.Y_DELTA_PATTERN_i43_LC_13_21_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i43_LC_13_21_2 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i43_LC_13_21_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i43_LC_13_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14581),
            .lcout(\transmit_module.Y_DELTA_PATTERN_43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22486),
            .ce(N__21436),
            .sr(N__21344));
    defparam \transmit_module.Y_DELTA_PATTERN_i46_LC_13_21_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i46_LC_13_21_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i46_LC_13_21_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i46_LC_13_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14563),
            .lcout(\transmit_module.Y_DELTA_PATTERN_46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22486),
            .ce(N__21436),
            .sr(N__21344));
    defparam \transmit_module.Y_DELTA_PATTERN_i44_LC_13_21_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i44_LC_13_21_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i44_LC_13_21_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i44_LC_13_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14569),
            .lcout(\transmit_module.Y_DELTA_PATTERN_44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22486),
            .ce(N__21436),
            .sr(N__21344));
    defparam \transmit_module.Y_DELTA_PATTERN_i45_LC_13_21_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i45_LC_13_21_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i45_LC_13_21_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i45_LC_13_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14575),
            .lcout(\transmit_module.Y_DELTA_PATTERN_45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22486),
            .ce(N__21436),
            .sr(N__21344));
    defparam \transmit_module.Y_DELTA_PATTERN_i47_LC_13_21_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i47_LC_13_21_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i47_LC_13_21_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i47_LC_13_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14557),
            .lcout(\transmit_module.Y_DELTA_PATTERN_47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22486),
            .ce(N__21436),
            .sr(N__21344));
    defparam \transmit_module.Y_DELTA_PATTERN_i53_LC_13_22_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i53_LC_13_22_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i53_LC_13_22_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i53_LC_13_22_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14692),
            .lcout(\transmit_module.Y_DELTA_PATTERN_53 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22322),
            .ce(N__21464),
            .sr(N__21166));
    defparam \transmit_module.Y_DELTA_PATTERN_i48_LC_13_22_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i48_LC_13_22_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i48_LC_13_22_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i48_LC_13_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14698),
            .lcout(\transmit_module.Y_DELTA_PATTERN_48 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22322),
            .ce(N__21464),
            .sr(N__21166));
    defparam \transmit_module.Y_DELTA_PATTERN_i52_LC_13_22_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i52_LC_13_22_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i52_LC_13_22_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i52_LC_13_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14551),
            .lcout(\transmit_module.Y_DELTA_PATTERN_52 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22322),
            .ce(N__21464),
            .sr(N__21166));
    defparam \transmit_module.Y_DELTA_PATTERN_i49_LC_13_22_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i49_LC_13_22_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i49_LC_13_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i49_LC_13_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14680),
            .lcout(\transmit_module.Y_DELTA_PATTERN_49 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22322),
            .ce(N__21464),
            .sr(N__21166));
    defparam \transmit_module.Y_DELTA_PATTERN_i54_LC_13_22_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i54_LC_13_22_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i54_LC_13_22_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i54_LC_13_22_5  (
            .in0(N__14668),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.Y_DELTA_PATTERN_54 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22322),
            .ce(N__21464),
            .sr(N__21166));
    defparam \transmit_module.Y_DELTA_PATTERN_i50_LC_13_22_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i50_LC_13_22_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i50_LC_13_22_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i50_LC_13_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14686),
            .lcout(\transmit_module.Y_DELTA_PATTERN_50 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22322),
            .ce(N__21464),
            .sr(N__21166));
    defparam \transmit_module.Y_DELTA_PATTERN_i59_LC_13_23_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i59_LC_13_23_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i59_LC_13_23_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i59_LC_13_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14644),
            .lcout(\transmit_module.Y_DELTA_PATTERN_59 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22409),
            .ce(N__21437),
            .sr(N__21345));
    defparam \transmit_module.Y_DELTA_PATTERN_i55_LC_13_23_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i55_LC_13_23_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i55_LC_13_23_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i55_LC_13_23_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14674),
            .lcout(\transmit_module.Y_DELTA_PATTERN_55 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22409),
            .ce(N__21437),
            .sr(N__21345));
    defparam \transmit_module.Y_DELTA_PATTERN_i58_LC_13_23_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i58_LC_13_23_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i58_LC_13_23_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i58_LC_13_23_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14662),
            .lcout(\transmit_module.Y_DELTA_PATTERN_58 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22409),
            .ce(N__21437),
            .sr(N__21345));
    defparam \transmit_module.Y_DELTA_PATTERN_i60_LC_13_23_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i60_LC_13_23_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i60_LC_13_23_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i60_LC_13_23_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14650),
            .lcout(\transmit_module.Y_DELTA_PATTERN_60 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22409),
            .ce(N__21437),
            .sr(N__21345));
    defparam \transmit_module.ADDR_Y_COMPONENT__i6_LC_13_24_0 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i6_LC_13_24_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i6_LC_13_24_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i6_LC_13_24_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17758),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22282),
            .ce(N__19882),
            .sr(N__21269));
    defparam \line_buffer.i2627_3_lut_LC_13_25_7 .C_ON=1'b0;
    defparam \line_buffer.i2627_3_lut_LC_13_25_7 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2627_3_lut_LC_13_25_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \line_buffer.i2627_3_lut_LC_13_25_7  (
            .in0(N__14638),
            .in1(N__14620),
            .in2(_gnd_net_),
            .in3(N__23553),
            .lcout(\line_buffer.n4101 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1769_4_lut_LC_13_31_7 .C_ON=1'b0;
    defparam \transmit_module.i1769_4_lut_LC_13_31_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1769_4_lut_LC_13_31_7 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \transmit_module.i1769_4_lut_LC_13_31_7  (
            .in0(N__16414),
            .in1(N__16345),
            .in2(N__21346),
            .in3(N__20241),
            .lcout(n22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i1_2_lut_adj_25_LC_14_8_0 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i1_2_lut_adj_25_LC_14_8_0 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i1_2_lut_adj_25_LC_14_8_0 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \receive_module.rx_counter.i1_2_lut_adj_25_LC_14_8_0  (
            .in0(_gnd_net_),
            .in1(N__17157),
            .in2(_gnd_net_),
            .in3(N__17187),
            .lcout(),
            .ltout(\receive_module.rx_counter.n5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i3_4_lut_adj_26_LC_14_8_1 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i3_4_lut_adj_26_LC_14_8_1 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i3_4_lut_adj_26_LC_14_8_1 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \receive_module.rx_counter.i3_4_lut_adj_26_LC_14_8_1  (
            .in0(N__16392),
            .in1(N__17139),
            .in2(N__15445),
            .in3(N__15403),
            .lcout(\receive_module.rx_counter.n11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i28_1_lut_rep_23_LC_14_8_6.C_ON=1'b0;
    defparam i28_1_lut_rep_23_LC_14_8_6.SEQ_MODE=4'b0000;
    defparam i28_1_lut_rep_23_LC_14_8_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 i28_1_lut_rep_23_LC_14_8_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15440),
            .lcout(n4214),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i1_2_lut_adj_24_LC_14_8_7 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i1_2_lut_adj_24_LC_14_8_7 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i1_2_lut_adj_24_LC_14_8_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \receive_module.rx_counter.i1_2_lut_adj_24_LC_14_8_7  (
            .in0(_gnd_net_),
            .in1(N__16377),
            .in2(_gnd_net_),
            .in3(N__17172),
            .lcout(\receive_module.rx_counter.n4_adj_576 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.X_277__i1_LC_14_9_0 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_277__i1_LC_14_9_0 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_277__i1_LC_14_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_277__i1_LC_14_9_0  (
            .in0(_gnd_net_),
            .in1(N__15185),
            .in2(_gnd_net_),
            .in3(N__15166),
            .lcout(RX_ADDR_0),
            .ltout(),
            .carryin(bfn_14_9_0_),
            .carryout(\receive_module.rx_counter.n3720 ),
            .clk(N__19326),
            .ce(),
            .sr(N__15952));
    defparam \receive_module.rx_counter.X_277__i2_LC_14_9_1 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_277__i2_LC_14_9_1 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_277__i2_LC_14_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_277__i2_LC_14_9_1  (
            .in0(_gnd_net_),
            .in1(N__14954),
            .in2(_gnd_net_),
            .in3(N__14932),
            .lcout(RX_ADDR_1),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3720 ),
            .carryout(\receive_module.rx_counter.n3721 ),
            .clk(N__19326),
            .ce(),
            .sr(N__15952));
    defparam \receive_module.rx_counter.X_277__i3_LC_14_9_2 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_277__i3_LC_14_9_2 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_277__i3_LC_14_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_277__i3_LC_14_9_2  (
            .in0(_gnd_net_),
            .in1(N__14723),
            .in2(_gnd_net_),
            .in3(N__14701),
            .lcout(RX_ADDR_2),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3721 ),
            .carryout(\receive_module.rx_counter.n3722 ),
            .clk(N__19326),
            .ce(),
            .sr(N__15952));
    defparam \receive_module.rx_counter.X_277__i4_LC_14_9_3 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_277__i4_LC_14_9_3 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_277__i4_LC_14_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_277__i4_LC_14_9_3  (
            .in0(_gnd_net_),
            .in1(N__17029),
            .in2(_gnd_net_),
            .in3(N__15973),
            .lcout(\receive_module.rx_counter.X_3 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3722 ),
            .carryout(\receive_module.rx_counter.n3723 ),
            .clk(N__19326),
            .ce(),
            .sr(N__15952));
    defparam \receive_module.rx_counter.X_277__i5_LC_14_9_4 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_277__i5_LC_14_9_4 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_277__i5_LC_14_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_277__i5_LC_14_9_4  (
            .in0(_gnd_net_),
            .in1(N__17050),
            .in2(_gnd_net_),
            .in3(N__15970),
            .lcout(\receive_module.rx_counter.X_4 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3723 ),
            .carryout(\receive_module.rx_counter.n3724 ),
            .clk(N__19326),
            .ce(),
            .sr(N__15952));
    defparam \receive_module.rx_counter.X_277__i6_LC_14_9_5 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_277__i6_LC_14_9_5 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_277__i6_LC_14_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_277__i6_LC_14_9_5  (
            .in0(_gnd_net_),
            .in1(N__17073),
            .in2(_gnd_net_),
            .in3(N__15967),
            .lcout(\receive_module.rx_counter.X_5 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3724 ),
            .carryout(\receive_module.rx_counter.n3725 ),
            .clk(N__19326),
            .ce(),
            .sr(N__15952));
    defparam \receive_module.rx_counter.X_277__i7_LC_14_9_6 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_277__i7_LC_14_9_6 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_277__i7_LC_14_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_277__i7_LC_14_9_6  (
            .in0(_gnd_net_),
            .in1(N__17412),
            .in2(_gnd_net_),
            .in3(N__15964),
            .lcout(\receive_module.rx_counter.X_6 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3725 ),
            .carryout(\receive_module.rx_counter.n3726 ),
            .clk(N__19326),
            .ce(),
            .sr(N__15952));
    defparam \receive_module.rx_counter.X_277__i8_LC_14_9_7 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_277__i8_LC_14_9_7 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_277__i8_LC_14_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_277__i8_LC_14_9_7  (
            .in0(_gnd_net_),
            .in1(N__17442),
            .in2(_gnd_net_),
            .in3(N__15961),
            .lcout(\receive_module.rx_counter.X_7 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3726 ),
            .carryout(\receive_module.rx_counter.n3727 ),
            .clk(N__19326),
            .ce(),
            .sr(N__15952));
    defparam \receive_module.rx_counter.X_277__i9_LC_14_10_0 .C_ON=1'b1;
    defparam \receive_module.rx_counter.X_277__i9_LC_14_10_0 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_277__i9_LC_14_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_277__i9_LC_14_10_0  (
            .in0(_gnd_net_),
            .in1(N__17502),
            .in2(_gnd_net_),
            .in3(N__15958),
            .lcout(\receive_module.rx_counter.X_8 ),
            .ltout(),
            .carryin(bfn_14_10_0_),
            .carryout(\receive_module.rx_counter.n3728 ),
            .clk(N__19330),
            .ce(),
            .sr(N__15948));
    defparam \receive_module.rx_counter.X_277__i10_LC_14_10_1 .C_ON=1'b0;
    defparam \receive_module.rx_counter.X_277__i10_LC_14_10_1 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.X_277__i10_LC_14_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.X_277__i10_LC_14_10_1  (
            .in0(_gnd_net_),
            .in1(N__17475),
            .in2(_gnd_net_),
            .in3(N__15955),
            .lcout(\receive_module.rx_counter.X_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19330),
            .ce(),
            .sr(N__15948));
    defparam \receive_module.rx_counter.i1_2_lut_4_lut_adj_27_LC_14_11_2 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i1_2_lut_4_lut_adj_27_LC_14_11_2 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i1_2_lut_4_lut_adj_27_LC_14_11_2 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \receive_module.rx_counter.i1_2_lut_4_lut_adj_27_LC_14_11_2  (
            .in0(N__15930),
            .in1(N__15891),
            .in2(N__15852),
            .in3(N__15761),
            .lcout(n658),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.X_DELTA_PATTERN_i9_LC_14_14_0 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i9_LC_14_14_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i9_LC_14_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i9_LC_14_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16066),
            .lcout(\transmit_module.X_DELTA_PATTERN_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22619),
            .ce(N__17578),
            .sr(N__20565));
    defparam \transmit_module.X_DELTA_PATTERN_i12_LC_14_14_3 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i12_LC_14_14_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.X_DELTA_PATTERN_i12_LC_14_14_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i12_LC_14_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16090),
            .lcout(\transmit_module.X_DELTA_PATTERN_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22619),
            .ce(N__17578),
            .sr(N__20565));
    defparam \transmit_module.X_DELTA_PATTERN_i13_LC_14_14_4 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i13_LC_14_14_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i13_LC_14_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i13_LC_14_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17629),
            .lcout(\transmit_module.X_DELTA_PATTERN_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22619),
            .ce(N__17578),
            .sr(N__20565));
    defparam \transmit_module.X_DELTA_PATTERN_i8_LC_14_14_5 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i8_LC_14_14_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.X_DELTA_PATTERN_i8_LC_14_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i8_LC_14_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16084),
            .lcout(\transmit_module.X_DELTA_PATTERN_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22619),
            .ce(N__17578),
            .sr(N__20565));
    defparam \transmit_module.X_DELTA_PATTERN_i11_LC_14_14_6 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i11_LC_14_14_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i11_LC_14_14_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i11_LC_14_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16078),
            .lcout(\transmit_module.X_DELTA_PATTERN_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22619),
            .ce(N__17578),
            .sr(N__20565));
    defparam \transmit_module.X_DELTA_PATTERN_i10_LC_14_14_7 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i10_LC_14_14_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.X_DELTA_PATTERN_i10_LC_14_14_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i10_LC_14_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16072),
            .lcout(\transmit_module.X_DELTA_PATTERN_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22619),
            .ce(N__17578),
            .sr(N__20565));
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_2663_LC_14_15_2 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_2663_LC_14_15_2 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_2663_LC_14_15_2 .LUT_INIT=16'b1100111110100000;
    LogicCell40 \line_buffer.TX_ADDR_12__bdd_4_lut_2663_LC_14_15_2  (
            .in0(N__17281),
            .in1(N__16060),
            .in2(N__22858),
            .in3(N__23836),
            .lcout(\line_buffer.n4134 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i2_4_lut_LC_14_15_5 .C_ON=1'b0;
    defparam \transmit_module.i2_4_lut_LC_14_15_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i2_4_lut_LC_14_15_5 .LUT_INIT=16'b1111111011110000;
    LogicCell40 \transmit_module.i2_4_lut_LC_14_15_5  (
            .in0(N__19583),
            .in1(N__19120),
            .in2(N__21194),
            .in3(N__19525),
            .lcout(\transmit_module.n2315 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.X_DELTA_PATTERN_i0_LC_14_16_0 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i0_LC_14_16_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i0_LC_14_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i0_LC_14_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17614),
            .lcout(\transmit_module.X_DELTA_PATTERN_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22560),
            .ce(N__17583),
            .sr(N__16025));
    defparam \transmit_module.ADDR_Y_COMPONENT__i4_LC_14_17_3 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i4_LC_14_17_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i4_LC_14_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i4_LC_14_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18991),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22498),
            .ce(N__19876),
            .sr(N__21317));
    defparam \transmit_module.ADDR_Y_COMPONENT__i2_LC_14_17_6 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i2_LC_14_17_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i2_LC_14_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i2_LC_14_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17824),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22498),
            .ce(N__19876),
            .sr(N__21317));
    defparam \transmit_module.BRAM_ADDR__i8_LC_14_18_0 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i8_LC_14_18_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i8_LC_14_18_0 .LUT_INIT=16'b0000000011100100;
    LogicCell40 \transmit_module.BRAM_ADDR__i8_LC_14_18_0  (
            .in0(N__20195),
            .in1(N__16987),
            .in2(N__17008),
            .in3(N__21209),
            .lcout(\transmit_module.TX_ADDR_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22470),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i0_LC_14_18_1 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i0_LC_14_18_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i0_LC_14_18_1 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \transmit_module.BRAM_ADDR__i0_LC_14_18_1  (
            .in0(N__17838),
            .in1(N__16360),
            .in2(N__21292),
            .in3(N__20191),
            .lcout(\transmit_module.TX_ADDR_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22470),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i10_3_lut_LC_14_18_2 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i10_3_lut_LC_14_18_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i10_3_lut_LC_14_18_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_12_i10_3_lut_LC_14_18_2  (
            .in0(N__19697),
            .in1(N__18433),
            .in2(_gnd_net_),
            .in3(N__18457),
            .lcout(\transmit_module.n179 ),
            .ltout(\transmit_module.n179_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i9_LC_14_18_3 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i9_LC_14_18_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i9_LC_14_18_3 .LUT_INIT=16'b0101000001000100;
    LogicCell40 \transmit_module.BRAM_ADDR__i9_LC_14_18_3  (
            .in0(N__21198),
            .in1(N__16321),
            .in2(N__16348),
            .in3(N__20196),
            .lcout(\transmit_module.TX_ADDR_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22470),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i7_LC_14_18_4 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i7_LC_14_18_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i7_LC_14_18_4 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \transmit_module.BRAM_ADDR__i7_LC_14_18_4  (
            .in0(N__20194),
            .in1(N__21199),
            .in2(N__16663),
            .in3(N__16654),
            .lcout(\transmit_module.TX_ADDR_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22470),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i6_LC_14_18_5 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i6_LC_14_18_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i6_LC_14_18_5 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \transmit_module.BRAM_ADDR__i6_LC_14_18_5  (
            .in0(N__16413),
            .in1(N__16341),
            .in2(N__21294),
            .in3(N__20193),
            .lcout(\transmit_module.TX_ADDR_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22470),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i143_2_lut_3_lut_4_lut_rep_33_LC_14_18_6 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i143_2_lut_3_lut_4_lut_rep_33_LC_14_18_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i143_2_lut_3_lut_4_lut_rep_33_LC_14_18_6 .LUT_INIT=16'b1100110011101100;
    LogicCell40 \transmit_module.video_signal_controller.i143_2_lut_3_lut_4_lut_rep_33_LC_14_18_6  (
            .in0(N__16760),
            .in1(N__21197),
            .in2(N__19533),
            .in3(N__16719),
            .lcout(\transmit_module.n4224 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i3_LC_14_18_7 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i3_LC_14_18_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i3_LC_14_18_7 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \transmit_module.BRAM_ADDR__i3_LC_14_18_7  (
            .in0(N__20274),
            .in1(N__20259),
            .in2(N__21293),
            .in3(N__20192),
            .lcout(\transmit_module.TX_ADDR_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22470),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1772_4_lut_LC_14_19_0 .C_ON=1'b0;
    defparam \transmit_module.i1772_4_lut_LC_14_19_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1772_4_lut_LC_14_19_0 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \transmit_module.i1772_4_lut_LC_14_19_0  (
            .in0(N__16327),
            .in1(N__16320),
            .in2(N__21180),
            .in3(N__20170),
            .lcout(n19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1771_4_lut_LC_14_19_1 .C_ON=1'b0;
    defparam \transmit_module.i1771_4_lut_LC_14_19_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1771_4_lut_LC_14_19_1 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \transmit_module.i1771_4_lut_LC_14_19_1  (
            .in0(N__20169),
            .in1(N__21034),
            .in2(N__17004),
            .in3(N__16986),
            .lcout(n20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_29_LC_14_19_2 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_29_LC_14_19_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.i1_2_lut_rep_29_LC_14_19_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \transmit_module.video_signal_controller.i1_2_lut_rep_29_LC_14_19_2  (
            .in0(_gnd_net_),
            .in1(N__16755),
            .in2(_gnd_net_),
            .in3(N__16718),
            .lcout(\transmit_module.n4220 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i8_3_lut_LC_14_19_3 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i8_3_lut_LC_14_19_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i8_3_lut_LC_14_19_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_12_i8_3_lut_LC_14_19_3  (
            .in0(N__19701),
            .in1(N__16429),
            .in2(_gnd_net_),
            .in3(N__17708),
            .lcout(\transmit_module.n181 ),
            .ltout(\transmit_module.n181_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1770_4_lut_LC_14_19_4 .C_ON=1'b0;
    defparam \transmit_module.i1770_4_lut_LC_14_19_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1770_4_lut_LC_14_19_4 .LUT_INIT=16'b0101000001000100;
    LogicCell40 \transmit_module.i1770_4_lut_LC_14_19_4  (
            .in0(N__21033),
            .in1(N__16653),
            .in2(N__16642),
            .in3(N__20168),
            .lcout(n21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.ADDR_Y_COMPONENT__i7_LC_14_21_3 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i7_LC_14_21_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i7_LC_14_21_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i7_LC_14_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17713),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22347),
            .ce(N__19869),
            .sr(N__21307));
    defparam \transmit_module.ADDR_Y_COMPONENT__i1_LC_14_22_7 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i1_LC_14_22_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i1_LC_14_22_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i1_LC_14_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18322),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22314),
            .ce(N__19875),
            .sr(N__21340));
    defparam \transmit_module.mux_12_i7_3_lut_LC_14_24_3 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i7_3_lut_LC_14_24_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i7_3_lut_LC_14_24_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_12_i7_3_lut_LC_14_24_3  (
            .in0(N__19713),
            .in1(N__16420),
            .in2(_gnd_net_),
            .in3(N__17757),
            .lcout(\transmit_module.n182 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.FRAME_COUNTER_278__i0_LC_15_8_0 .C_ON=1'b1;
    defparam \receive_module.rx_counter.FRAME_COUNTER_278__i0_LC_15_8_0 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.FRAME_COUNTER_278__i0_LC_15_8_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.FRAME_COUNTER_278__i0_LC_15_8_0  (
            .in0(_gnd_net_),
            .in1(N__16393),
            .in2(_gnd_net_),
            .in3(N__16381),
            .lcout(\receive_module.rx_counter.FRAME_COUNTER_0 ),
            .ltout(),
            .carryin(bfn_15_8_0_),
            .carryout(\receive_module.rx_counter.n3706 ),
            .clk(N__19322),
            .ce(N__17332),
            .sr(N__17128));
    defparam \receive_module.rx_counter.FRAME_COUNTER_278__i1_LC_15_8_1 .C_ON=1'b1;
    defparam \receive_module.rx_counter.FRAME_COUNTER_278__i1_LC_15_8_1 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.FRAME_COUNTER_278__i1_LC_15_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.FRAME_COUNTER_278__i1_LC_15_8_1  (
            .in0(_gnd_net_),
            .in1(N__16378),
            .in2(_gnd_net_),
            .in3(N__17191),
            .lcout(\receive_module.rx_counter.FRAME_COUNTER_1 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3706 ),
            .carryout(\receive_module.rx_counter.n3707 ),
            .clk(N__19322),
            .ce(N__17332),
            .sr(N__17128));
    defparam \receive_module.rx_counter.FRAME_COUNTER_278__i2_LC_15_8_2 .C_ON=1'b1;
    defparam \receive_module.rx_counter.FRAME_COUNTER_278__i2_LC_15_8_2 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.FRAME_COUNTER_278__i2_LC_15_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.FRAME_COUNTER_278__i2_LC_15_8_2  (
            .in0(_gnd_net_),
            .in1(N__17188),
            .in2(_gnd_net_),
            .in3(N__17176),
            .lcout(\receive_module.rx_counter.FRAME_COUNTER_2 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3707 ),
            .carryout(\receive_module.rx_counter.n3708 ),
            .clk(N__19322),
            .ce(N__17332),
            .sr(N__17128));
    defparam \receive_module.rx_counter.FRAME_COUNTER_278__i3_LC_15_8_3 .C_ON=1'b1;
    defparam \receive_module.rx_counter.FRAME_COUNTER_278__i3_LC_15_8_3 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.FRAME_COUNTER_278__i3_LC_15_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.FRAME_COUNTER_278__i3_LC_15_8_3  (
            .in0(_gnd_net_),
            .in1(N__17173),
            .in2(_gnd_net_),
            .in3(N__17161),
            .lcout(\receive_module.rx_counter.FRAME_COUNTER_3 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3708 ),
            .carryout(\receive_module.rx_counter.n3709 ),
            .clk(N__19322),
            .ce(N__17332),
            .sr(N__17128));
    defparam \receive_module.rx_counter.FRAME_COUNTER_278__i4_LC_15_8_4 .C_ON=1'b1;
    defparam \receive_module.rx_counter.FRAME_COUNTER_278__i4_LC_15_8_4 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.FRAME_COUNTER_278__i4_LC_15_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.FRAME_COUNTER_278__i4_LC_15_8_4  (
            .in0(_gnd_net_),
            .in1(N__17158),
            .in2(_gnd_net_),
            .in3(N__17146),
            .lcout(\receive_module.rx_counter.FRAME_COUNTER_4 ),
            .ltout(),
            .carryin(\receive_module.rx_counter.n3709 ),
            .carryout(\receive_module.rx_counter.n3710 ),
            .clk(N__19322),
            .ce(N__17332),
            .sr(N__17128));
    defparam \receive_module.rx_counter.FRAME_COUNTER_278__i5_LC_15_8_5 .C_ON=1'b0;
    defparam \receive_module.rx_counter.FRAME_COUNTER_278__i5_LC_15_8_5 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.FRAME_COUNTER_278__i5_LC_15_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \receive_module.rx_counter.FRAME_COUNTER_278__i5_LC_15_8_5  (
            .in0(_gnd_net_),
            .in1(N__17140),
            .in2(_gnd_net_),
            .in3(N__17143),
            .lcout(\receive_module.rx_counter.FRAME_COUNTER_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19322),
            .ce(N__17332),
            .sr(N__17128));
    defparam \receive_module.rx_counter.old_VS_51_LC_15_9_0 .C_ON=1'b0;
    defparam \receive_module.rx_counter.old_VS_51_LC_15_9_0 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.old_VS_51_LC_15_9_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \receive_module.rx_counter.old_VS_51_LC_15_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17099),
            .lcout(\receive_module.rx_counter.old_VS ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19324),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i1360_2_lut_3_lut_LC_15_9_1 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i1360_2_lut_3_lut_LC_15_9_1 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i1360_2_lut_3_lut_LC_15_9_1 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \receive_module.rx_counter.i1360_2_lut_3_lut_LC_15_9_1  (
            .in0(N__17097),
            .in1(N__17118),
            .in2(_gnd_net_),
            .in3(N__17370),
            .lcout(\receive_module.rx_counter.n2605 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i150_2_lut_rep_31_LC_15_9_2 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i150_2_lut_rep_31_LC_15_9_2 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i150_2_lut_rep_31_LC_15_9_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \receive_module.rx_counter.i150_2_lut_rep_31_LC_15_9_2  (
            .in0(N__17119),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17098),
            .lcout(\receive_module.rx_counter.n4222 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i2_3_lut_rep_28_LC_15_9_3 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i2_3_lut_rep_28_LC_15_9_3 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i2_3_lut_rep_28_LC_15_9_3 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \receive_module.rx_counter.i2_3_lut_rep_28_LC_15_9_3  (
            .in0(N__17072),
            .in1(N__17049),
            .in2(_gnd_net_),
            .in3(N__17028),
            .lcout(\receive_module.rx_counter.n4219 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i1_2_lut_adj_20_LC_15_10_1 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i1_2_lut_adj_20_LC_15_10_1 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i1_2_lut_adj_20_LC_15_10_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \receive_module.rx_counter.i1_2_lut_adj_20_LC_15_10_1  (
            .in0(_gnd_net_),
            .in1(N__17498),
            .in2(_gnd_net_),
            .in3(N__17471),
            .lcout(),
            .ltout(\receive_module.rx_counter.n4_adj_575_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.i2_4_lut_adj_21_LC_15_10_2 .C_ON=1'b0;
    defparam \receive_module.rx_counter.i2_4_lut_adj_21_LC_15_10_2 .SEQ_MODE=4'b0000;
    defparam \receive_module.rx_counter.i2_4_lut_adj_21_LC_15_10_2 .LUT_INIT=16'b1111110011111000;
    LogicCell40 \receive_module.rx_counter.i2_4_lut_adj_21_LC_15_10_2  (
            .in0(N__17449),
            .in1(N__17441),
            .in2(N__17419),
            .in3(N__17408),
            .lcout(\receive_module.rx_counter.O_VISIBLE_N_86 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \receive_module.rx_counter.PULSE_1HZ_48_LC_15_10_3 .C_ON=1'b0;
    defparam \receive_module.rx_counter.PULSE_1HZ_48_LC_15_10_3 .SEQ_MODE=4'b1000;
    defparam \receive_module.rx_counter.PULSE_1HZ_48_LC_15_10_3 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \receive_module.rx_counter.PULSE_1HZ_48_LC_15_10_3  (
            .in0(N__17374),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17343),
            .lcout(LED_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__19327),
            .ce(N__17331),
            .sr(_gnd_net_));
    defparam \line_buffer.i2597_3_lut_LC_15_13_1 .C_ON=1'b0;
    defparam \line_buffer.i2597_3_lut_LC_15_13_1 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2597_3_lut_LC_15_13_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \line_buffer.i2597_3_lut_LC_15_13_1  (
            .in0(N__23492),
            .in1(N__17320),
            .in2(_gnd_net_),
            .in3(N__17302),
            .lcout(\line_buffer.n4071 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2698_LC_15_13_6 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2698_LC_15_13_6 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2698_LC_15_13_6 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_2698_LC_15_13_6  (
            .in0(N__17272),
            .in1(N__23846),
            .in2(N__17260),
            .in3(N__23493),
            .lcout(),
            .ltout(\line_buffer.n4176_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n4176_bdd_4_lut_LC_15_13_7 .C_ON=1'b0;
    defparam \line_buffer.n4176_bdd_4_lut_LC_15_13_7 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n4176_bdd_4_lut_LC_15_13_7 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \line_buffer.n4176_bdd_4_lut_LC_15_13_7  (
            .in0(N__23847),
            .in1(N__17239),
            .in2(N__17218),
            .in3(N__17215),
            .lcout(\line_buffer.n4179 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.X_DELTA_PATTERN_i7_LC_15_14_1 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i7_LC_15_14_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i7_LC_15_14_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i7_LC_15_14_1  (
            .in0(N__17197),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.X_DELTA_PATTERN_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22514),
            .ce(N__17582),
            .sr(N__20587));
    defparam \transmit_module.X_DELTA_PATTERN_i5_LC_15_15_5 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i5_LC_15_15_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.X_DELTA_PATTERN_i5_LC_15_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i5_LC_15_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17635),
            .lcout(\transmit_module.X_DELTA_PATTERN_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22513),
            .ce(N__17571),
            .sr(N__20583));
    defparam \transmit_module.X_DELTA_PATTERN_i6_LC_15_15_6 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i6_LC_15_15_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i6_LC_15_15_6 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i6_LC_15_15_6  (
            .in0(_gnd_net_),
            .in1(N__17641),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.X_DELTA_PATTERN_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22513),
            .ce(N__17571),
            .sr(N__20583));
    defparam \transmit_module.X_DELTA_PATTERN_i14_LC_15_16_0 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i14_LC_15_16_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.X_DELTA_PATTERN_i14_LC_15_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i14_LC_15_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17602),
            .lcout(\transmit_module.X_DELTA_PATTERN_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22248),
            .ce(N__17584),
            .sr(N__20550));
    defparam \transmit_module.X_DELTA_PATTERN_i2_LC_15_16_1 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i2_LC_15_16_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i2_LC_15_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i2_LC_15_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17608),
            .lcout(\transmit_module.X_DELTA_PATTERN_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22248),
            .ce(N__17584),
            .sr(N__20550));
    defparam \transmit_module.X_DELTA_PATTERN_i1_LC_15_16_4 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i1_LC_15_16_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.X_DELTA_PATTERN_i1_LC_15_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i1_LC_15_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17620),
            .lcout(\transmit_module.X_DELTA_PATTERN_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22248),
            .ce(N__17584),
            .sr(N__20550));
    defparam \transmit_module.X_DELTA_PATTERN_i3_LC_15_16_5 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i3_LC_15_16_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.X_DELTA_PATTERN_i3_LC_15_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i3_LC_15_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17590),
            .lcout(\transmit_module.X_DELTA_PATTERN_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22248),
            .ce(N__17584),
            .sr(N__20550));
    defparam \transmit_module.X_DELTA_PATTERN_i15_LC_15_16_6 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i15_LC_15_16_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i15_LC_15_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i15_LC_15_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17535),
            .lcout(\transmit_module.X_DELTA_PATTERN_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22248),
            .ce(N__17584),
            .sr(N__20550));
    defparam \transmit_module.X_DELTA_PATTERN_i4_LC_15_16_7 .C_ON=1'b0;
    defparam \transmit_module.X_DELTA_PATTERN_i4_LC_15_16_7 .SEQ_MODE=4'b1001;
    defparam \transmit_module.X_DELTA_PATTERN_i4_LC_15_16_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \transmit_module.X_DELTA_PATTERN_i4_LC_15_16_7  (
            .in0(N__17596),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.X_DELTA_PATTERN_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22248),
            .ce(N__17584),
            .sr(N__20550));
    defparam \transmit_module.add_13_2_lut_LC_15_17_0 .C_ON=1'b1;
    defparam \transmit_module.add_13_2_lut_LC_15_17_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_2_lut_LC_15_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_2_lut_LC_15_17_0  (
            .in0(_gnd_net_),
            .in1(N__18406),
            .in2(N__17536),
            .in3(_gnd_net_),
            .lcout(\transmit_module.n204 ),
            .ltout(),
            .carryin(bfn_15_17_0_),
            .carryout(\transmit_module.n3656 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_3_lut_LC_15_17_1 .C_ON=1'b1;
    defparam \transmit_module.add_13_3_lut_LC_15_17_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_3_lut_LC_15_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_3_lut_LC_15_17_1  (
            .in0(_gnd_net_),
            .in1(N__18320),
            .in2(_gnd_net_),
            .in3(N__17506),
            .lcout(\transmit_module.n203 ),
            .ltout(),
            .carryin(\transmit_module.n3656 ),
            .carryout(\transmit_module.n3657 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_4_lut_LC_15_17_2 .C_ON=1'b1;
    defparam \transmit_module.add_13_4_lut_LC_15_17_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_4_lut_LC_15_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_4_lut_LC_15_17_2  (
            .in0(_gnd_net_),
            .in1(N__17823),
            .in2(_gnd_net_),
            .in3(N__17785),
            .lcout(\transmit_module.n202 ),
            .ltout(),
            .carryin(\transmit_module.n3657 ),
            .carryout(\transmit_module.n3658 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_5_lut_LC_15_17_3 .C_ON=1'b1;
    defparam \transmit_module.add_13_5_lut_LC_15_17_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_5_lut_LC_15_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_5_lut_LC_15_17_3  (
            .in0(_gnd_net_),
            .in1(N__18373),
            .in2(_gnd_net_),
            .in3(N__17767),
            .lcout(\transmit_module.n201 ),
            .ltout(),
            .carryin(\transmit_module.n3658 ),
            .carryout(\transmit_module.n3659 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_6_lut_LC_15_17_4 .C_ON=1'b1;
    defparam \transmit_module.add_13_6_lut_LC_15_17_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_6_lut_LC_15_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_6_lut_LC_15_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18987),
            .in3(N__17764),
            .lcout(\transmit_module.n200 ),
            .ltout(),
            .carryin(\transmit_module.n3659 ),
            .carryout(\transmit_module.n3660 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_7_lut_LC_15_17_5 .C_ON=1'b1;
    defparam \transmit_module.add_13_7_lut_LC_15_17_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_7_lut_LC_15_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_7_lut_LC_15_17_5  (
            .in0(_gnd_net_),
            .in1(N__19021),
            .in2(_gnd_net_),
            .in3(N__17761),
            .lcout(\transmit_module.n199 ),
            .ltout(),
            .carryin(\transmit_module.n3660 ),
            .carryout(\transmit_module.n3661 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_8_lut_LC_15_17_6 .C_ON=1'b1;
    defparam \transmit_module.add_13_8_lut_LC_15_17_6 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_8_lut_LC_15_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_8_lut_LC_15_17_6  (
            .in0(_gnd_net_),
            .in1(N__17741),
            .in2(_gnd_net_),
            .in3(N__17716),
            .lcout(\transmit_module.n198 ),
            .ltout(),
            .carryin(\transmit_module.n3661 ),
            .carryout(\transmit_module.n3662 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_9_lut_LC_15_17_7 .C_ON=1'b1;
    defparam \transmit_module.add_13_9_lut_LC_15_17_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_9_lut_LC_15_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_9_lut_LC_15_17_7  (
            .in0(_gnd_net_),
            .in1(N__17704),
            .in2(_gnd_net_),
            .in3(N__17671),
            .lcout(\transmit_module.n197 ),
            .ltout(),
            .carryin(\transmit_module.n3662 ),
            .carryout(\transmit_module.n3663 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_10_lut_LC_15_18_0 .C_ON=1'b1;
    defparam \transmit_module.add_13_10_lut_LC_15_18_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_10_lut_LC_15_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_10_lut_LC_15_18_0  (
            .in0(_gnd_net_),
            .in1(N__17884),
            .in2(_gnd_net_),
            .in3(N__17656),
            .lcout(\transmit_module.n196 ),
            .ltout(),
            .carryin(bfn_15_18_0_),
            .carryout(\transmit_module.n3664 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_11_lut_LC_15_18_1 .C_ON=1'b1;
    defparam \transmit_module.add_13_11_lut_LC_15_18_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_11_lut_LC_15_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_11_lut_LC_15_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18464),
            .in3(N__17644),
            .lcout(\transmit_module.n195 ),
            .ltout(),
            .carryin(\transmit_module.n3664 ),
            .carryout(\transmit_module.n3665 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_12_lut_LC_15_18_2 .C_ON=1'b1;
    defparam \transmit_module.add_13_12_lut_LC_15_18_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_12_lut_LC_15_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_12_lut_LC_15_18_2  (
            .in0(_gnd_net_),
            .in1(N__17956),
            .in2(_gnd_net_),
            .in3(N__17905),
            .lcout(\transmit_module.n194 ),
            .ltout(),
            .carryin(\transmit_module.n3665 ),
            .carryout(\transmit_module.n3666 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_13_lut_LC_15_18_3 .C_ON=1'b1;
    defparam \transmit_module.add_13_13_lut_LC_15_18_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_13_lut_LC_15_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_13_lut_LC_15_18_3  (
            .in0(_gnd_net_),
            .in1(N__23518),
            .in2(_gnd_net_),
            .in3(N__17902),
            .lcout(\transmit_module.n193 ),
            .ltout(),
            .carryin(\transmit_module.n3666 ),
            .carryout(\transmit_module.n3667 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_14_lut_LC_15_18_4 .C_ON=1'b1;
    defparam \transmit_module.add_13_14_lut_LC_15_18_4 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_14_lut_LC_15_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \transmit_module.add_13_14_lut_LC_15_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23806),
            .in3(N__17899),
            .lcout(\transmit_module.n192 ),
            .ltout(),
            .carryin(\transmit_module.n3667 ),
            .carryout(\transmit_module.n3668 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.add_13_15_lut_LC_15_18_5 .C_ON=1'b0;
    defparam \transmit_module.add_13_15_lut_LC_15_18_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.add_13_15_lut_LC_15_18_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \transmit_module.add_13_15_lut_LC_15_18_5  (
            .in0(N__22802),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17896),
            .lcout(\transmit_module.n191 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.ADDR_Y_COMPONENT__i8_LC_15_18_7 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i8_LC_15_18_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i8_LC_15_18_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i8_LC_15_18_7  (
            .in0(N__17885),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22445),
            .ce(N__19853),
            .sr(N__21210));
    defparam \transmit_module.mux_12_i4_3_lut_LC_15_19_1 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i4_3_lut_LC_15_19_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i4_3_lut_LC_15_19_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \transmit_module.mux_12_i4_3_lut_LC_15_19_1  (
            .in0(N__18352),
            .in1(N__19670),
            .in2(_gnd_net_),
            .in3(N__18374),
            .lcout(\transmit_module.n185 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.mux_14_i2_3_lut_4_lut_LC_15_19_3 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.mux_14_i2_3_lut_4_lut_LC_15_19_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.mux_14_i2_3_lut_4_lut_LC_15_19_3 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \transmit_module.video_signal_controller.mux_14_i2_3_lut_4_lut_LC_15_19_3  (
            .in0(N__18319),
            .in1(N__19128),
            .in2(N__17854),
            .in3(N__19521),
            .lcout(\transmit_module.n218 ),
            .ltout(\transmit_module.n218_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i1_LC_15_19_4 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i1_LC_15_19_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i1_LC_15_19_4 .LUT_INIT=16'b0100010001010000;
    LogicCell40 \transmit_module.BRAM_ADDR__i1_LC_15_19_4  (
            .in0(N__21179),
            .in1(N__18292),
            .in2(N__17842),
            .in3(N__20209),
            .lcout(\transmit_module.TX_ADDR_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22352),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i1_3_lut_LC_15_19_7 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i1_3_lut_LC_15_19_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i1_3_lut_LC_15_19_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_12_i1_3_lut_LC_15_19_7  (
            .in0(N__19691),
            .in1(N__18385),
            .in2(_gnd_net_),
            .in3(N__18407),
            .lcout(\transmit_module.n188 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.ADDR_Y_COMPONENT__i0_LC_15_20_0 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i0_LC_15_20_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i0_LC_15_20_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i0_LC_15_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18421),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22070),
            .ce(N__19874),
            .sr(N__21181));
    defparam \transmit_module.ADDR_Y_COMPONENT__i11_LC_15_20_1 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i11_LC_15_20_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i11_LC_15_20_1 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i11_LC_15_20_1  (
            .in0(_gnd_net_),
            .in1(N__23485),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22070),
            .ce(N__19874),
            .sr(N__21181));
    defparam \transmit_module.ADDR_Y_COMPONENT__i3_LC_15_20_6 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i3_LC_15_20_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i3_LC_15_20_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i3_LC_15_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18379),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22070),
            .ce(N__19874),
            .sr(N__21181));
    defparam \transmit_module.BRAM_ADDR__rep_1_i0_LC_15_21_0 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__rep_1_i0_LC_15_21_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__rep_1_i0_LC_15_21_0 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \transmit_module.BRAM_ADDR__rep_1_i0_LC_15_21_0  (
            .in0(N__19582),
            .in1(N__18346),
            .in2(N__18337),
            .in3(N__19532),
            .lcout(TX_ADDR_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22062),
            .ce(N__19410),
            .sr(N__21338));
    defparam \transmit_module.mux_12_i2_3_lut_LC_15_22_2 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i2_3_lut_LC_15_22_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i2_3_lut_LC_15_22_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_12_i2_3_lut_LC_15_22_2  (
            .in0(N__19693),
            .in1(N__18328),
            .in2(_gnd_net_),
            .in3(N__18321),
            .lcout(\transmit_module.n187 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1764_4_lut_LC_15_27_1 .C_ON=1'b0;
    defparam \transmit_module.i1764_4_lut_LC_15_27_1 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1764_4_lut_LC_15_27_1 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \transmit_module.i1764_4_lut_LC_15_27_1  (
            .in0(N__18291),
            .in1(N__18274),
            .in2(N__21336),
            .in3(N__20240),
            .lcout(n27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_LC_16_13_3 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_LC_16_13_3 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_LC_16_13_3 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_LC_16_13_3  (
            .in0(N__18049),
            .in1(N__23848),
            .in2(N__18031),
            .in3(N__23611),
            .lcout(),
            .ltout(\line_buffer.n4188_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n4188_bdd_4_lut_LC_16_13_4 .C_ON=1'b0;
    defparam \line_buffer.n4188_bdd_4_lut_LC_16_13_4 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n4188_bdd_4_lut_LC_16_13_4 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \line_buffer.n4188_bdd_4_lut_LC_16_13_4  (
            .in0(N__23849),
            .in1(N__18019),
            .in2(N__18001),
            .in3(N__17998),
            .lcout(),
            .ltout(\line_buffer.n4191_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i5_LC_16_13_5 .C_ON=1'b0;
    defparam \line_buffer.dout_i5_LC_16_13_5 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i5_LC_16_13_5 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \line_buffer.dout_i5_LC_16_13_5  (
            .in0(_gnd_net_),
            .in1(N__22856),
            .in2(N__17980),
            .in3(N__17977),
            .lcout(TX_DATA_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22421),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.Y_DELTA_PATTERN_i18_LC_16_16_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i18_LC_16_16_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i18_LC_16_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i18_LC_16_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18481),
            .lcout(\transmit_module.Y_DELTA_PATTERN_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22247),
            .ce(N__20597),
            .sr(N__21147));
    defparam \transmit_module.Y_DELTA_PATTERN_i20_LC_16_16_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i20_LC_16_16_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i20_LC_16_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i20_LC_16_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18493),
            .lcout(\transmit_module.Y_DELTA_PATTERN_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22247),
            .ce(N__20597),
            .sr(N__21147));
    defparam \transmit_module.Y_DELTA_PATTERN_i0_LC_16_16_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i0_LC_16_16_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i0_LC_16_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i0_LC_16_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18475),
            .lcout(\transmit_module.Y_DELTA_PATTERN_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22247),
            .ce(N__20597),
            .sr(N__21147));
    defparam \transmit_module.Y_DELTA_PATTERN_i17_LC_16_16_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i17_LC_16_16_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i17_LC_16_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i17_LC_16_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18499),
            .lcout(\transmit_module.Y_DELTA_PATTERN_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22247),
            .ce(N__20597),
            .sr(N__21147));
    defparam \transmit_module.Y_DELTA_PATTERN_i21_LC_16_16_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i21_LC_16_16_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i21_LC_16_16_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i21_LC_16_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20647),
            .lcout(\transmit_module.Y_DELTA_PATTERN_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22247),
            .ce(N__20597),
            .sr(N__21147));
    defparam \transmit_module.Y_DELTA_PATTERN_i19_LC_16_16_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i19_LC_16_16_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i19_LC_16_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i19_LC_16_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18487),
            .lcout(\transmit_module.Y_DELTA_PATTERN_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22247),
            .ce(N__20597),
            .sr(N__21147));
    defparam \transmit_module.Y_DELTA_PATTERN_i1_LC_16_16_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i1_LC_16_16_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i1_LC_16_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i1_LC_16_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20656),
            .lcout(\transmit_module.Y_DELTA_PATTERN_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22247),
            .ce(N__20597),
            .sr(N__21147));
    defparam \transmit_module.ADDR_Y_COMPONENT__i5_LC_16_17_5 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i5_LC_16_17_5 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i5_LC_16_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i5_LC_16_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19026),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22243),
            .ce(N__19877),
            .sr(N__21341));
    defparam \transmit_module.ADDR_Y_COMPONENT__i9_LC_16_17_6 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i9_LC_16_17_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i9_LC_16_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i9_LC_16_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18469),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22243),
            .ce(N__19877),
            .sr(N__21341));
    defparam \transmit_module.video_signal_controller.mux_14_i5_3_lut_4_lut_LC_16_18_0 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.mux_14_i5_3_lut_4_lut_LC_16_18_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.mux_14_i5_3_lut_4_lut_LC_16_18_0 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \transmit_module.video_signal_controller.mux_14_i5_3_lut_4_lut_LC_16_18_0  (
            .in0(N__18983),
            .in1(N__19126),
            .in2(N__19174),
            .in3(N__19512),
            .lcout(\transmit_module.n215 ),
            .ltout(\transmit_module.n215_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i4_LC_16_18_1 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i4_LC_16_18_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i4_LC_16_18_1 .LUT_INIT=16'b0100010001010000;
    LogicCell40 \transmit_module.BRAM_ADDR__i4_LC_16_18_1  (
            .in0(N__21217),
            .in1(N__18961),
            .in2(N__19165),
            .in3(N__20228),
            .lcout(\transmit_module.TX_ADDR_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22444),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i6_3_lut_LC_16_18_2 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i6_3_lut_LC_16_18_2 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i6_3_lut_LC_16_18_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_12_i6_3_lut_LC_16_18_2  (
            .in0(N__19663),
            .in1(N__19162),
            .in2(_gnd_net_),
            .in3(N__19022),
            .lcout(\transmit_module.n183 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.mux_18_i14_3_lut_4_lut_LC_16_18_3 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.mux_18_i14_3_lut_4_lut_LC_16_18_3 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.mux_18_i14_3_lut_4_lut_LC_16_18_3 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \transmit_module.video_signal_controller.mux_18_i14_3_lut_4_lut_LC_16_18_3  (
            .in0(N__19513),
            .in1(N__19587),
            .in2(N__19897),
            .in3(N__19156),
            .lcout(\transmit_module.BRAM_ADDR_13_N_258_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.video_signal_controller.mux_14_i6_3_lut_4_lut_LC_16_18_5 .C_ON=1'b0;
    defparam \transmit_module.video_signal_controller.mux_14_i6_3_lut_4_lut_LC_16_18_5 .SEQ_MODE=4'b0000;
    defparam \transmit_module.video_signal_controller.mux_14_i6_3_lut_4_lut_LC_16_18_5 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \transmit_module.video_signal_controller.mux_14_i6_3_lut_4_lut_LC_16_18_5  (
            .in0(N__19511),
            .in1(N__19138),
            .in2(N__19027),
            .in3(N__19127),
            .lcout(\transmit_module.n214 ),
            .ltout(\transmit_module.n214_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i5_LC_16_18_6 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i5_LC_16_18_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i5_LC_16_18_6 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \transmit_module.BRAM_ADDR__i5_LC_16_18_6  (
            .in0(N__20229),
            .in1(N__21218),
            .in2(N__19030),
            .in3(N__18732),
            .lcout(\transmit_module.TX_ADDR_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22444),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.mux_12_i5_3_lut_LC_16_18_7 .C_ON=1'b0;
    defparam \transmit_module.mux_12_i5_3_lut_LC_16_18_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.mux_12_i5_3_lut_LC_16_18_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \transmit_module.mux_12_i5_3_lut_LC_16_18_7  (
            .in0(N__19662),
            .in1(N__19003),
            .in2(_gnd_net_),
            .in3(N__18982),
            .lcout(\transmit_module.n184 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1767_4_lut_LC_16_19_0 .C_ON=1'b0;
    defparam \transmit_module.i1767_4_lut_LC_16_19_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1767_4_lut_LC_16_19_0 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \transmit_module.i1767_4_lut_LC_16_19_0  (
            .in0(N__18960),
            .in1(N__18949),
            .in2(N__21280),
            .in3(N__20197),
            .lcout(n24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.i1768_4_lut_LC_16_19_7 .C_ON=1'b0;
    defparam \transmit_module.i1768_4_lut_LC_16_19_7 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1768_4_lut_LC_16_19_7 .LUT_INIT=16'b0011000100100000;
    LogicCell40 \transmit_module.i1768_4_lut_LC_16_19_7  (
            .in0(N__20198),
            .in1(N__21172),
            .in2(N__18733),
            .in3(N__18718),
            .lcout(n23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.BRAM_ADDR__i12_LC_16_20_7 .C_ON=1'b0;
    defparam \transmit_module.BRAM_ADDR__i12_LC_16_20_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.BRAM_ADDR__i12_LC_16_20_7 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \transmit_module.BRAM_ADDR__i12_LC_16_20_7  (
            .in0(N__19588),
            .in1(N__19543),
            .in2(N__19906),
            .in3(N__19534),
            .lcout(TX_ADDR_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22069),
            .ce(N__19411),
            .sr(N__21260));
    defparam \transmit_module.Y_DELTA_PATTERN_i41_LC_16_21_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i41_LC_16_21_6 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i41_LC_16_21_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i41_LC_16_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19381),
            .lcout(\transmit_module.Y_DELTA_PATTERN_41 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22061),
            .ce(N__21459),
            .sr(N__21339));
    defparam GB_BUFFER_DEBUG_c_1_c_THRU_LUT4_0_LC_16_30_5.C_ON=1'b0;
    defparam GB_BUFFER_DEBUG_c_1_c_THRU_LUT4_0_LC_16_30_5.SEQ_MODE=4'b0000;
    defparam GB_BUFFER_DEBUG_c_1_c_THRU_LUT4_0_LC_16_30_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 GB_BUFFER_DEBUG_c_1_c_THRU_LUT4_0_LC_16_30_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19372),
            .lcout(GB_BUFFER_DEBUG_c_1_c_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.Y_DELTA_PATTERN_i5_LC_17_14_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i5_LC_17_14_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i5_LC_17_14_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i5_LC_17_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20350),
            .lcout(\transmit_module.Y_DELTA_PATTERN_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22565),
            .ce(N__20622),
            .sr(N__21295));
    defparam \transmit_module.Y_DELTA_PATTERN_i28_LC_17_15_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i28_LC_17_15_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i28_LC_17_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i28_LC_17_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19192),
            .lcout(\transmit_module.Y_DELTA_PATTERN_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22420),
            .ce(N__20599),
            .sr(N__21266));
    defparam \transmit_module.Y_DELTA_PATTERN_i31_LC_17_15_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i31_LC_17_15_1 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i31_LC_17_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i31_LC_17_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19762),
            .lcout(\transmit_module.Y_DELTA_PATTERN_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22420),
            .ce(N__20599),
            .sr(N__21266));
    defparam \transmit_module.Y_DELTA_PATTERN_i29_LC_17_15_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i29_LC_17_15_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i29_LC_17_15_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i29_LC_17_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19180),
            .lcout(\transmit_module.Y_DELTA_PATTERN_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22420),
            .ce(N__20599),
            .sr(N__21266));
    defparam \transmit_module.Y_DELTA_PATTERN_i30_LC_17_15_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i30_LC_17_15_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i30_LC_17_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i30_LC_17_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19186),
            .lcout(\transmit_module.Y_DELTA_PATTERN_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22420),
            .ce(N__20599),
            .sr(N__21266));
    defparam \transmit_module.Y_DELTA_PATTERN_i12_LC_17_16_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i12_LC_17_16_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i12_LC_17_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i12_LC_17_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19756),
            .lcout(\transmit_module.Y_DELTA_PATTERN_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22548),
            .ce(N__20614),
            .sr(N__21324));
    defparam \transmit_module.Y_DELTA_PATTERN_i11_LC_17_16_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i11_LC_17_16_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i11_LC_17_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i11_LC_17_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19768),
            .lcout(\transmit_module.Y_DELTA_PATTERN_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22548),
            .ce(N__20614),
            .sr(N__21324));
    defparam \transmit_module.Y_DELTA_PATTERN_i32_LC_17_16_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i32_LC_17_16_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i32_LC_17_16_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i32_LC_17_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21523),
            .lcout(\transmit_module.Y_DELTA_PATTERN_32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22548),
            .ce(N__20614),
            .sr(N__21324));
    defparam \transmit_module.Y_DELTA_PATTERN_i13_LC_17_16_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i13_LC_17_16_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i13_LC_17_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i13_LC_17_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19750),
            .lcout(\transmit_module.Y_DELTA_PATTERN_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22548),
            .ce(N__20614),
            .sr(N__21324));
    defparam \transmit_module.Y_DELTA_PATTERN_i14_LC_17_16_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i14_LC_17_16_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i14_LC_17_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i14_LC_17_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20308),
            .lcout(\transmit_module.Y_DELTA_PATTERN_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22548),
            .ce(N__20614),
            .sr(N__21324));
    defparam \transmit_module.Y_DELTA_PATTERN_i26_LC_17_17_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i26_LC_17_17_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i26_LC_17_17_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i26_LC_17_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19723),
            .lcout(\transmit_module.Y_DELTA_PATTERN_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22573),
            .ce(N__20598),
            .sr(N__21343));
    defparam \transmit_module.Y_DELTA_PATTERN_i24_LC_17_17_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i24_LC_17_17_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i24_LC_17_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i24_LC_17_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19738),
            .lcout(\transmit_module.Y_DELTA_PATTERN_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22573),
            .ce(N__20598),
            .sr(N__21343));
    defparam \transmit_module.Y_DELTA_PATTERN_i25_LC_17_17_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i25_LC_17_17_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i25_LC_17_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i25_LC_17_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19744),
            .lcout(\transmit_module.Y_DELTA_PATTERN_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22573),
            .ce(N__20598),
            .sr(N__21343));
    defparam \transmit_module.Y_DELTA_PATTERN_i27_LC_17_17_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i27_LC_17_17_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i27_LC_17_17_5 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i27_LC_17_17_5  (
            .in0(_gnd_net_),
            .in1(N__19732),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.Y_DELTA_PATTERN_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22573),
            .ce(N__20598),
            .sr(N__21343));
    defparam \transmit_module.Y_DELTA_PATTERN_i99_LC_17_17_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i99_LC_17_17_7 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i99_LC_17_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i99_LC_17_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19661),
            .lcout(\transmit_module.Y_DELTA_PATTERN_99 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22573),
            .ce(N__20598),
            .sr(N__21343));
    defparam \transmit_module.Y_DELTA_PATTERN_i37_LC_17_18_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i37_LC_17_18_0 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i37_LC_17_18_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i37_LC_17_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20281),
            .lcout(\transmit_module.Y_DELTA_PATTERN_37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22466),
            .ce(N__21473),
            .sr(N__21262));
    defparam \transmit_module.Y_DELTA_PATTERN_i35_LC_17_18_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i35_LC_17_18_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i35_LC_17_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i35_LC_17_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20287),
            .lcout(\transmit_module.Y_DELTA_PATTERN_35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22466),
            .ce(N__21473),
            .sr(N__21262));
    defparam \transmit_module.Y_DELTA_PATTERN_i36_LC_17_18_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i36_LC_17_18_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i36_LC_17_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i36_LC_17_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20293),
            .lcout(\transmit_module.Y_DELTA_PATTERN_36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22466),
            .ce(N__21473),
            .sr(N__21262));
    defparam \transmit_module.Y_DELTA_PATTERN_i38_LC_17_18_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i38_LC_17_18_7 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i38_LC_17_18_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i38_LC_17_18_7  (
            .in0(N__19789),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.Y_DELTA_PATTERN_38 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22466),
            .ce(N__21473),
            .sr(N__21262));
    defparam \transmit_module.i1766_4_lut_LC_17_19_0 .C_ON=1'b0;
    defparam \transmit_module.i1766_4_lut_LC_17_19_0 .SEQ_MODE=4'b0000;
    defparam \transmit_module.i1766_4_lut_LC_17_19_0 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \transmit_module.i1766_4_lut_LC_17_19_0  (
            .in0(N__20275),
            .in1(N__20260),
            .in2(N__21281),
            .in3(N__20216),
            .lcout(n25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.ADDR_Y_COMPONENT__i12_LC_17_20_2 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i12_LC_17_20_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i12_LC_17_20_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i12_LC_17_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23741),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22440),
            .ce(N__19870),
            .sr(N__21261));
    defparam \transmit_module.ADDR_Y_COMPONENT__i13_LC_17_20_3 .C_ON=1'b0;
    defparam \transmit_module.ADDR_Y_COMPONENT__i13_LC_17_20_3 .SEQ_MODE=4'b1000;
    defparam \transmit_module.ADDR_Y_COMPONENT__i13_LC_17_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.ADDR_Y_COMPONENT__i13_LC_17_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22818),
            .lcout(\transmit_module.ADDR_Y_COMPONENT_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22440),
            .ce(N__19870),
            .sr(N__21261));
    defparam \transmit_module.Y_DELTA_PATTERN_i39_LC_17_21_2 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i39_LC_17_21_2 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i39_LC_17_21_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i39_LC_17_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19774),
            .lcout(\transmit_module.Y_DELTA_PATTERN_39 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22340),
            .ce(N__21487),
            .sr(N__21337));
    defparam \transmit_module.Y_DELTA_PATTERN_i40_LC_17_21_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i40_LC_17_21_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i40_LC_17_21_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i40_LC_17_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19780),
            .lcout(\transmit_module.Y_DELTA_PATTERN_40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22340),
            .ce(N__21487),
            .sr(N__21337));
    defparam \line_buffer.i2591_3_lut_LC_18_9_4 .C_ON=1'b0;
    defparam \line_buffer.i2591_3_lut_LC_18_9_4 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2591_3_lut_LC_18_9_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \line_buffer.i2591_3_lut_LC_18_9_4  (
            .in0(N__20377),
            .in1(N__20359),
            .in2(_gnd_net_),
            .in3(N__23535),
            .lcout(\line_buffer.n4065 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.Y_DELTA_PATTERN_i6_LC_18_14_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i6_LC_18_14_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i6_LC_18_14_0 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i6_LC_18_14_0  (
            .in0(_gnd_net_),
            .in1(N__20338),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.Y_DELTA_PATTERN_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22572),
            .ce(N__20623),
            .sr(N__21296));
    defparam \transmit_module.Y_DELTA_PATTERN_i4_LC_18_14_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i4_LC_18_14_7 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i4_LC_18_14_7 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i4_LC_18_14_7  (
            .in0(_gnd_net_),
            .in1(N__20344),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.Y_DELTA_PATTERN_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22572),
            .ce(N__20623),
            .sr(N__21296));
    defparam \transmit_module.Y_DELTA_PATTERN_i9_LC_18_15_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i9_LC_18_15_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i9_LC_18_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i9_LC_18_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20326),
            .lcout(\transmit_module.Y_DELTA_PATTERN_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22419),
            .ce(N__20618),
            .sr(N__21323));
    defparam \transmit_module.Y_DELTA_PATTERN_i7_LC_18_15_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i7_LC_18_15_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i7_LC_18_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i7_LC_18_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20314),
            .lcout(\transmit_module.Y_DELTA_PATTERN_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22419),
            .ce(N__20618),
            .sr(N__21323));
    defparam \transmit_module.Y_DELTA_PATTERN_i10_LC_18_15_3 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i10_LC_18_15_3 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i10_LC_18_15_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i10_LC_18_15_3  (
            .in0(N__20332),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\transmit_module.Y_DELTA_PATTERN_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22419),
            .ce(N__20618),
            .sr(N__21323));
    defparam \transmit_module.Y_DELTA_PATTERN_i8_LC_18_15_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i8_LC_18_15_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i8_LC_18_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i8_LC_18_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20320),
            .lcout(\transmit_module.Y_DELTA_PATTERN_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22419),
            .ce(N__20618),
            .sr(N__21323));
    defparam \transmit_module.Y_DELTA_PATTERN_i15_LC_18_16_1 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i15_LC_18_16_1 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i15_LC_18_16_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i15_LC_18_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20668),
            .lcout(\transmit_module.Y_DELTA_PATTERN_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22562),
            .ce(N__20607),
            .sr(N__21267));
    defparam \transmit_module.Y_DELTA_PATTERN_i3_LC_18_16_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i3_LC_18_16_4 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i3_LC_18_16_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i3_LC_18_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20302),
            .lcout(\transmit_module.Y_DELTA_PATTERN_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22562),
            .ce(N__20607),
            .sr(N__21267));
    defparam \transmit_module.Y_DELTA_PATTERN_i16_LC_18_16_6 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i16_LC_18_16_6 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i16_LC_18_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i16_LC_18_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20677),
            .lcout(\transmit_module.Y_DELTA_PATTERN_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22562),
            .ce(N__20607),
            .sr(N__21267));
    defparam \transmit_module.Y_DELTA_PATTERN_i2_LC_18_16_7 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i2_LC_18_16_7 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i2_LC_18_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i2_LC_18_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20662),
            .lcout(\transmit_module.Y_DELTA_PATTERN_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22562),
            .ce(N__20607),
            .sr(N__21267));
    defparam \transmit_module.Y_DELTA_PATTERN_i22_LC_18_17_4 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i22_LC_18_17_4 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i22_LC_18_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i22_LC_18_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20629),
            .lcout(\transmit_module.Y_DELTA_PATTERN_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22512),
            .ce(N__20606),
            .sr(N__21342));
    defparam \transmit_module.Y_DELTA_PATTERN_i23_LC_18_17_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i23_LC_18_17_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i23_LC_18_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i23_LC_18_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20635),
            .lcout(\transmit_module.Y_DELTA_PATTERN_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22512),
            .ce(N__20606),
            .sr(N__21342));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2688_LC_18_18_5 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2688_LC_18_18_5 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2688_LC_18_18_5 .LUT_INIT=16'b1110010010101010;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_2688_LC_18_18_5  (
            .in0(N__23602),
            .in1(N__20485),
            .in2(N__20470),
            .in3(N__23842),
            .lcout(),
            .ltout(\line_buffer.n4164_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n4164_bdd_4_lut_LC_18_18_6 .C_ON=1'b0;
    defparam \line_buffer.n4164_bdd_4_lut_LC_18_18_6 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n4164_bdd_4_lut_LC_18_18_6 .LUT_INIT=16'b1111010010100100;
    LogicCell40 \line_buffer.n4164_bdd_4_lut_LC_18_18_6  (
            .in0(N__23843),
            .in1(N__20449),
            .in2(N__20428),
            .in3(N__20425),
            .lcout(),
            .ltout(\line_buffer.n4167_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i1_LC_18_18_7 .C_ON=1'b0;
    defparam \line_buffer.dout_i1_LC_18_18_7 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i1_LC_18_18_7 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \line_buffer.dout_i1_LC_18_18_7  (
            .in0(_gnd_net_),
            .in1(N__22835),
            .in2(N__20407),
            .in3(N__20683),
            .lcout(TX_DATA_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22474),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_2658_LC_18_19_0 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_2658_LC_18_19_0 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_2658_LC_18_19_0 .LUT_INIT=16'b1100111110100000;
    LogicCell40 \line_buffer.TX_ADDR_12__bdd_4_lut_2658_LC_18_19_0  (
            .in0(N__20389),
            .in1(N__21628),
            .in2(N__22857),
            .in3(N__23829),
            .lcout(\line_buffer.n4128 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2592_3_lut_LC_18_20_0 .C_ON=1'b0;
    defparam \line_buffer.i2592_3_lut_LC_18_20_0 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2592_3_lut_LC_18_20_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \line_buffer.i2592_3_lut_LC_18_20_0  (
            .in0(N__21664),
            .in1(N__21646),
            .in2(_gnd_net_),
            .in3(N__23598),
            .lcout(\line_buffer.n4066 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2600_3_lut_LC_18_20_1 .C_ON=1'b0;
    defparam \line_buffer.i2600_3_lut_LC_18_20_1 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2600_3_lut_LC_18_20_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \line_buffer.i2600_3_lut_LC_18_20_1  (
            .in0(N__23600),
            .in1(N__21622),
            .in2(_gnd_net_),
            .in3(N__21607),
            .lcout(),
            .ltout(\line_buffer.n4074_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i3_LC_18_20_2 .C_ON=1'b0;
    defparam \line_buffer.dout_i3_LC_18_20_2 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i3_LC_18_20_2 .LUT_INIT=16'b1110111001010000;
    LogicCell40 \line_buffer.dout_i3_LC_18_20_2  (
            .in0(N__22819),
            .in1(N__21529),
            .in2(N__21589),
            .in3(N__21586),
            .lcout(TX_DATA_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22465),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2601_3_lut_LC_18_20_3 .C_ON=1'b0;
    defparam \line_buffer.i2601_3_lut_LC_18_20_3 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2601_3_lut_LC_18_20_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \line_buffer.i2601_3_lut_LC_18_20_3  (
            .in0(N__23599),
            .in1(N__21571),
            .in2(_gnd_net_),
            .in3(N__21547),
            .lcout(\line_buffer.n4075 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \transmit_module.Y_DELTA_PATTERN_i33_LC_19_17_0 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i33_LC_19_17_0 .SEQ_MODE=4'b1000;
    defparam \transmit_module.Y_DELTA_PATTERN_i33_LC_19_17_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i33_LC_19_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21499),
            .lcout(\transmit_module.Y_DELTA_PATTERN_33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22574),
            .ce(N__21488),
            .sr(N__21322));
    defparam \transmit_module.Y_DELTA_PATTERN_i34_LC_19_17_5 .C_ON=1'b0;
    defparam \transmit_module.Y_DELTA_PATTERN_i34_LC_19_17_5 .SEQ_MODE=4'b1001;
    defparam \transmit_module.Y_DELTA_PATTERN_i34_LC_19_17_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \transmit_module.Y_DELTA_PATTERN_i34_LC_19_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21511),
            .lcout(\transmit_module.Y_DELTA_PATTERN_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22574),
            .ce(N__21488),
            .sr(N__21322));
    defparam \line_buffer.n4146_bdd_4_lut_LC_19_18_6 .C_ON=1'b0;
    defparam \line_buffer.n4146_bdd_4_lut_LC_19_18_6 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n4146_bdd_4_lut_LC_19_18_6 .LUT_INIT=16'b1100110010111000;
    LogicCell40 \line_buffer.n4146_bdd_4_lut_LC_19_18_6  (
            .in0(N__20761),
            .in1(N__22972),
            .in2(N__20746),
            .in3(N__23841),
            .lcout(\line_buffer.n4149 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n4158_bdd_4_lut_LC_19_18_7 .C_ON=1'b0;
    defparam \line_buffer.n4158_bdd_4_lut_LC_19_18_7 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n4158_bdd_4_lut_LC_19_18_7 .LUT_INIT=16'b1111101001000100;
    LogicCell40 \line_buffer.n4158_bdd_4_lut_LC_19_18_7  (
            .in0(N__23840),
            .in1(N__20725),
            .in2(N__20707),
            .in3(N__23659),
            .lcout(\line_buffer.n4161 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2673_LC_19_19_0 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2673_LC_19_19_0 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2673_LC_19_19_0 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_2673_LC_19_19_0  (
            .in0(N__23011),
            .in1(N__23828),
            .in2(N__22990),
            .in3(N__23601),
            .lcout(\line_buffer.n4146 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i0_LC_19_19_6 .C_ON=1'b0;
    defparam \line_buffer.dout_i0_LC_19_19_6 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i0_LC_19_19_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \line_buffer.dout_i0_LC_19_19_6  (
            .in0(N__22842),
            .in1(N__21670),
            .in2(_gnd_net_),
            .in3(N__22966),
            .lcout(TX_DATA_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22487),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2588_3_lut_LC_20_9_0 .C_ON=1'b0;
    defparam \line_buffer.i2588_3_lut_LC_20_9_0 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2588_3_lut_LC_20_9_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \line_buffer.i2588_3_lut_LC_20_9_0  (
            .in0(N__22945),
            .in1(N__22933),
            .in2(_gnd_net_),
            .in3(N__23536),
            .lcout(\line_buffer.n4062 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2604_3_lut_LC_20_11_2 .C_ON=1'b0;
    defparam \line_buffer.i2604_3_lut_LC_20_11_2 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2604_3_lut_LC_20_11_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \line_buffer.i2604_3_lut_LC_20_11_2  (
            .in0(N__22918),
            .in1(N__22906),
            .in2(_gnd_net_),
            .in3(N__23614),
            .lcout(\line_buffer.n4078 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_LC_20_13_1 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_LC_20_13_1 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_12__bdd_4_lut_LC_20_13_1 .LUT_INIT=16'b1010111111000000;
    LogicCell40 \line_buffer.TX_ADDR_12__bdd_4_lut_LC_20_13_1  (
            .in0(N__23401),
            .in1(N__22891),
            .in2(N__22869),
            .in3(N__23859),
            .lcout(\line_buffer.n4140 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.dout_i4_LC_20_14_1 .C_ON=1'b0;
    defparam \line_buffer.dout_i4_LC_20_14_1 .SEQ_MODE=4'b1000;
    defparam \line_buffer.dout_i4_LC_20_14_1 .LUT_INIT=16'b1110111000110000;
    LogicCell40 \line_buffer.dout_i4_LC_20_14_1  (
            .in0(N__22882),
            .in1(N__22865),
            .in2(N__23893),
            .in3(N__22714),
            .lcout(TX_DATA_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__22621),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2649_LC_20_17_5 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2649_LC_20_17_5 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2649_LC_20_17_5 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_2649_LC_20_17_5  (
            .in0(N__21739),
            .in1(N__23850),
            .in2(N__21724),
            .in3(N__23577),
            .lcout(\line_buffer.n4116 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.n4116_bdd_4_lut_LC_20_18_1 .C_ON=1'b0;
    defparam \line_buffer.n4116_bdd_4_lut_LC_20_18_1 .SEQ_MODE=4'b0000;
    defparam \line_buffer.n4116_bdd_4_lut_LC_20_18_1 .LUT_INIT=16'b1100110010111000;
    LogicCell40 \line_buffer.n4116_bdd_4_lut_LC_20_18_1  (
            .in0(N__21709),
            .in1(N__21694),
            .in2(N__21688),
            .in3(N__23851),
            .lcout(\line_buffer.n4119 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2603_3_lut_LC_20_18_7 .C_ON=1'b0;
    defparam \line_buffer.i2603_3_lut_LC_20_18_7 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2603_3_lut_LC_20_18_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \line_buffer.i2603_3_lut_LC_20_18_7  (
            .in0(N__23590),
            .in1(N__23923),
            .in2(_gnd_net_),
            .in3(N__23908),
            .lcout(\line_buffer.n4077 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2683_LC_20_19_6 .C_ON=1'b0;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2683_LC_20_19_6 .SEQ_MODE=4'b0000;
    defparam \line_buffer.TX_ADDR_11__bdd_4_lut_2683_LC_20_19_6 .LUT_INIT=16'b1111001110001000;
    LogicCell40 \line_buffer.TX_ADDR_11__bdd_4_lut_2683_LC_20_19_6  (
            .in0(N__23881),
            .in1(N__23818),
            .in2(N__23674),
            .in3(N__23586),
            .lcout(\line_buffer.n4158 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \line_buffer.i2589_3_lut_LC_21_13_3 .C_ON=1'b0;
    defparam \line_buffer.i2589_3_lut_LC_21_13_3 .SEQ_MODE=4'b0000;
    defparam \line_buffer.i2589_3_lut_LC_21_13_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \line_buffer.i2589_3_lut_LC_21_13_3  (
            .in0(N__23653),
            .in1(N__23635),
            .in2(_gnd_net_),
            .in3(N__23612),
            .lcout(\line_buffer.n4063 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_24_24_1.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_24_24_1.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_24_24_1.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_24_24_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // main
